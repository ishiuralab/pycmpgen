module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    compressor_CLA486_32 compressor_CLA486_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA486_32(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [0:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [0:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], 1'h0, comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], 1'h0}),
        .dst({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [0:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [0:0] dst39,
      output wire [0:0] dst40);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [126:0] stage1_0;
   wire [137:0] stage1_1;
   wire [227:0] stage1_2;
   wire [187:0] stage1_3;
   wire [225:0] stage1_4;
   wire [217:0] stage1_5;
   wire [246:0] stage1_6;
   wire [223:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [187:0] stage1_10;
   wire [219:0] stage1_11;
   wire [281:0] stage1_12;
   wire [204:0] stage1_13;
   wire [296:0] stage1_14;
   wire [171:0] stage1_15;
   wire [264:0] stage1_16;
   wire [270:0] stage1_17;
   wire [200:0] stage1_18;
   wire [299:0] stage1_19;
   wire [188:0] stage1_20;
   wire [198:0] stage1_21;
   wire [250:0] stage1_22;
   wire [177:0] stage1_23;
   wire [211:0] stage1_24;
   wire [234:0] stage1_25;
   wire [214:0] stage1_26;
   wire [158:0] stage1_27;
   wire [251:0] stage1_28;
   wire [235:0] stage1_29;
   wire [171:0] stage1_30;
   wire [160:0] stage1_31;
   wire [150:0] stage1_32;
   wire [80:0] stage1_33;
   wire [21:0] stage2_0;
   wire [106:0] stage2_1;
   wire [50:0] stage2_2;
   wire [87:0] stage2_3;
   wire [90:0] stage2_4;
   wire [83:0] stage2_5;
   wire [93:0] stage2_6;
   wire [109:0] stage2_7;
   wire [107:0] stage2_8;
   wire [74:0] stage2_9;
   wire [88:0] stage2_10;
   wire [91:0] stage2_11;
   wire [102:0] stage2_12;
   wire [101:0] stage2_13;
   wire [138:0] stage2_14;
   wire [135:0] stage2_15;
   wire [103:0] stage2_16;
   wire [121:0] stage2_17;
   wire [81:0] stage2_18;
   wire [109:0] stage2_19;
   wire [127:0] stage2_20;
   wire [78:0] stage2_21;
   wire [78:0] stage2_22;
   wire [109:0] stage2_23;
   wire [99:0] stage2_24;
   wire [87:0] stage2_25;
   wire [98:0] stage2_26;
   wire [96:0] stage2_27;
   wire [74:0] stage2_28;
   wire [120:0] stage2_29;
   wire [129:0] stage2_30;
   wire [83:0] stage2_31;
   wire [64:0] stage2_32;
   wire [45:0] stage2_33;
   wire [35:0] stage2_34;
   wire [13:0] stage2_35;
   wire [7:0] stage3_0;
   wire [17:0] stage3_1;
   wire [31:0] stage3_2;
   wire [26:0] stage3_3;
   wire [43:0] stage3_4;
   wire [48:0] stage3_5;
   wire [42:0] stage3_6;
   wire [68:0] stage3_7;
   wire [37:0] stage3_8;
   wire [69:0] stage3_9;
   wire [28:0] stage3_10;
   wire [43:0] stage3_11;
   wire [41:0] stage3_12;
   wire [40:0] stage3_13;
   wire [50:0] stage3_14;
   wire [89:0] stage3_15;
   wire [61:0] stage3_16;
   wire [49:0] stage3_17;
   wire [49:0] stage3_18;
   wire [49:0] stage3_19;
   wire [45:0] stage3_20;
   wire [58:0] stage3_21;
   wire [46:0] stage3_22;
   wire [47:0] stage3_23;
   wire [40:0] stage3_24;
   wire [39:0] stage3_25;
   wire [31:0] stage3_26;
   wire [66:0] stage3_27;
   wire [42:0] stage3_28;
   wire [38:0] stage3_29;
   wire [59:0] stage3_30;
   wire [39:0] stage3_31;
   wire [35:0] stage3_32;
   wire [39:0] stage3_33;
   wire [21:0] stage3_34;
   wire [12:0] stage3_35;
   wire [6:0] stage3_36;
   wire [1:0] stage3_37;
   wire [2:0] stage4_0;
   wire [8:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [22:0] stage4_5;
   wire [20:0] stage4_6;
   wire [26:0] stage4_7;
   wire [22:0] stage4_8;
   wire [26:0] stage4_9;
   wire [28:0] stage4_10;
   wire [20:0] stage4_11;
   wire [13:0] stage4_12;
   wire [27:0] stage4_13;
   wire [12:0] stage4_14;
   wire [47:0] stage4_15;
   wire [28:0] stage4_16;
   wire [34:0] stage4_17;
   wire [18:0] stage4_18;
   wire [28:0] stage4_19;
   wire [25:0] stage4_20;
   wire [21:0] stage4_21;
   wire [22:0] stage4_22;
   wire [21:0] stage4_23;
   wire [30:0] stage4_24;
   wire [16:0] stage4_25;
   wire [23:0] stage4_26;
   wire [27:0] stage4_27;
   wire [17:0] stage4_28;
   wire [20:0] stage4_29;
   wire [22:0] stage4_30;
   wire [20:0] stage4_31;
   wire [18:0] stage4_32;
   wire [13:0] stage4_33;
   wire [16:0] stage4_34;
   wire [13:0] stage4_35;
   wire [9:0] stage4_36;
   wire [1:0] stage4_37;
   wire [0:0] stage4_38;
   wire [2:0] stage5_0;
   wire [8:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [3:0] stage5_4;
   wire [8:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [12:0] stage5_8;
   wire [11:0] stage5_9;
   wire [22:0] stage5_10;
   wire [8:0] stage5_11;
   wire [10:0] stage5_12;
   wire [15:0] stage5_13;
   wire [7:0] stage5_14;
   wire [10:0] stage5_15;
   wire [21:0] stage5_16;
   wire [14:0] stage5_17;
   wire [12:0] stage5_18;
   wire [12:0] stage5_19;
   wire [9:0] stage5_20;
   wire [10:0] stage5_21;
   wire [11:0] stage5_22;
   wire [13:0] stage5_23;
   wire [7:0] stage5_24;
   wire [7:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [11:0] stage5_30;
   wire [10:0] stage5_31;
   wire [10:0] stage5_32;
   wire [8:0] stage5_33;
   wire [7:0] stage5_34;
   wire [14:0] stage5_35;
   wire [3:0] stage5_36;
   wire [5:0] stage5_37;
   wire [1:0] stage5_38;
   wire [2:0] stage6_0;
   wire [6:0] stage6_1;
   wire [0:0] stage6_2;
   wire [3:0] stage6_3;
   wire [1:0] stage6_4;
   wire [5:0] stage6_5;
   wire [4:0] stage6_6;
   wire [2:0] stage6_7;
   wire [5:0] stage6_8;
   wire [4:0] stage6_9;
   wire [6:0] stage6_10;
   wire [5:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [4:0] stage6_22;
   wire [8:0] stage6_23;
   wire [3:0] stage6_24;
   wire [4:0] stage6_25;
   wire [11:0] stage6_26;
   wire [8:0] stage6_27;
   wire [6:0] stage6_28;
   wire [3:0] stage6_29;
   wire [4:0] stage6_30;
   wire [7:0] stage6_31;
   wire [3:0] stage6_32;
   wire [5:0] stage6_33;
   wire [10:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [1:0] stage6_37;
   wire [2:0] stage6_38;
   wire [0:0] stage6_39;
   wire [2:0] stage7_0;
   wire [6:0] stage7_1;
   wire [0:0] stage7_2;
   wire [3:0] stage7_3;
   wire [1:0] stage7_4;
   wire [3:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [1:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [2:0] stage7_19;
   wire [6:0] stage7_20;
   wire [0:0] stage7_21;
   wire [5:0] stage7_22;
   wire [5:0] stage7_23;
   wire [3:0] stage7_24;
   wire [0:0] stage7_25;
   wire [2:0] stage7_26;
   wire [5:0] stage7_27;
   wire [5:0] stage7_28;
   wire [3:0] stage7_29;
   wire [2:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [3:0] stage7_38;
   wire [0:0] stage7_39;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [0:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [0:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [0:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc1343_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3]},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[4]},
      {stage0_2[3]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[5]},
      {stage0_2[4]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[6]},
      {stage0_2[5]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_1[7]},
      {stage0_2[6]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[8]},
      {stage0_2[7]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[9]},
      {stage0_2[8]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[10]},
      {stage0_2[9]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[11]},
      {stage0_2[10]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[12]},
      {stage0_2[11]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[13]},
      {stage0_2[12]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[14]},
      {stage0_2[13]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[15]},
      {stage0_2[14]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[16]},
      {stage0_2[15]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc117_4 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[17]},
      {stage0_2[16]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc117_4 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[18]},
      {stage0_2[17]},
      {stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc117_4 gpc16 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[19]},
      {stage0_2[18]},
      {stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[19]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[20]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[21]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[22]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[23]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[24]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[25]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[26]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[27]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[28]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[29]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[30]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[31]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[32]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[33]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[34]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[35]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[36]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[37]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[38]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[39]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[40]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[41]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[42]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[43]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[44]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[27],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[28],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[29],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[30],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[31],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[32],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[33],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[34],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[35],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[36],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[37],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[38],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[39],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[40],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[41],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[42],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[43],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[44],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[45],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[46],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[47],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[48],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[49],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[50],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[51],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[52],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[53],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[54],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[55],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[56],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[57],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[58],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[59],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[60],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[61],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[62],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[63],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[64],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[65],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[66],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437], stage0_0[438]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[67],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc1325_5 gpc84 (
      {stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_1[176], stage0_1[177]},
      {stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage0_3[27]},
      {stage1_4[68],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[0],stage1_4[69],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[1],stage1_4[70],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[2],stage1_4[71],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[3],stage1_4[72],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[4],stage1_4[73],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[5],stage1_4[74],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[6],stage1_4[75],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[7],stage1_4[76],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[8],stage1_4[77],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[9],stage1_4[78],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[10],stage1_4[79],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[11],stage1_4[80],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[12],stage1_4[81],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[13],stage1_4[82],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[14],stage1_4[83],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[15],stage1_4[84],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279]},
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage1_5[16],stage1_4[85],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285]},
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135]},
      {stage1_5[17],stage1_4[86],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291]},
      {stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141]},
      {stage1_5[18],stage1_4[87],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297]},
      {stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147]},
      {stage1_5[19],stage1_4[88],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303]},
      {stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153]},
      {stage1_5[20],stage1_4[89],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309]},
      {stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159]},
      {stage1_5[21],stage1_4[90],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315]},
      {stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165]},
      {stage1_5[22],stage1_4[91],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321]},
      {stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage1_5[23],stage1_4[92],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327]},
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177]},
      {stage1_5[24],stage1_4[93],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333]},
      {stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183]},
      {stage1_5[25],stage1_4[94],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339]},
      {stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189]},
      {stage1_5[26],stage1_4[95],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345]},
      {stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195]},
      {stage1_5[27],stage1_4[96],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351]},
      {stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage1_5[28],stage1_4[97],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357]},
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207]},
      {stage1_5[29],stage1_4[98],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363]},
      {stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213]},
      {stage1_5[30],stage1_4[99],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369]},
      {stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219]},
      {stage1_5[31],stage1_4[100],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375]},
      {stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage1_5[32],stage1_4[101],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381]},
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage1_5[33],stage1_4[102],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387]},
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage1_5[34],stage1_4[103],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393]},
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243]},
      {stage1_5[35],stage1_4[104],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399]},
      {stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249]},
      {stage1_5[36],stage1_4[105],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405]},
      {stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255]},
      {stage1_5[37],stage1_4[106],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411]},
      {stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage1_5[38],stage1_4[107],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417]},
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267]},
      {stage1_5[39],stage1_4[108],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423]},
      {stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273]},
      {stage1_5[40],stage1_4[109],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429]},
      {stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279]},
      {stage1_5[41],stage1_4[110],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435]},
      {stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage1_5[42],stage1_4[111],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441]},
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage1_5[43],stage1_4[112],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447]},
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296], stage0_3[297]},
      {stage1_5[44],stage1_4[113],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453]},
      {stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302], stage0_3[303]},
      {stage1_5[45],stage1_4[114],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459]},
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309]},
      {stage1_5[46],stage1_4[115],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465]},
      {stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage1_5[47],stage1_4[116],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471]},
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage1_5[48],stage1_4[117],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477]},
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327]},
      {stage1_5[49],stage1_4[118],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[478], stage0_1[479], stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483]},
      {stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage1_5[50],stage1_4[119],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[51],stage1_4[120],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[52],stage1_4[121],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[53],stage1_4[122],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[54],stage1_4[123],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[55],stage1_4[124],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[56],stage1_4[125],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[57],stage1_4[126],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[58],stage1_4[127],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[59],stage1_4[128],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[60],stage1_4[129],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[61],stage1_4[130],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[62],stage1_4[131],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[63],stage1_4[132],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[64],stage1_4[133],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[65],stage1_4[134],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[66],stage1_4[135],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394]},
      {stage0_3[334]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[67],stage1_4[136],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399]},
      {stage0_3[335]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[68],stage1_4[137],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage0_3[336]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[69],stage1_4[138],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409]},
      {stage0_3[337]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[70],stage1_4[139],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage0_3[338]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[71],stage1_4[140],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[126]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[21],stage1_5[72],stage1_4[141],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[127]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[22],stage1_5[73],stage1_4[142],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[128]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[23],stage1_5[74],stage1_4[143],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[129]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[24],stage1_5[75],stage1_4[144],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[130]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[25],stage1_5[76],stage1_4[145],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[131]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[26],stage1_5[77],stage1_4[146],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[132]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[27],stage1_5[78],stage1_4[147],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[133]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[28],stage1_5[79],stage1_4[148],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[134]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[29],stage1_5[80],stage1_4[149],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[135]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[30],stage1_5[81],stage1_4[150],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[136]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[31],stage1_5[82],stage1_4[151],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[137]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[32],stage1_5[83],stage1_4[152],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[138]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[33],stage1_5[84],stage1_4[153],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[139]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[34],stage1_5[85],stage1_4[154],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[140]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[35],stage1_5[86],stage1_4[155],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[414], stage0_3[415], stage0_3[416], stage0_3[417], stage0_3[418]},
      {stage0_4[141]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[36],stage1_5[87],stage1_4[156],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422], stage0_3[423]},
      {stage0_4[142]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[37],stage1_5[88],stage1_4[157],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage0_4[143]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[38],stage1_5[89],stage1_4[158],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433]},
      {stage0_4[144]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[39],stage1_5[90],stage1_4[159],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[434], stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438]},
      {stage0_4[145]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[40],stage1_5[91],stage1_4[160],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[439], stage0_3[440], stage0_3[441], stage0_3[442], stage0_3[443]},
      {stage0_4[146]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[41],stage1_5[92],stage1_4[161],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[444], stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448]},
      {stage0_4[147]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[42],stage1_5[93],stage1_4[162],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[449], stage0_3[450], stage0_3[451], stage0_3[452], stage0_3[453]},
      {stage0_4[148]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[43],stage1_5[94],stage1_4[163],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[454], stage0_3[455], stage0_3[456], stage0_3[457], stage0_3[458]},
      {stage0_4[149]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[44],stage1_5[95],stage1_4[164],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[459], stage0_3[460], stage0_3[461], stage0_3[462], stage0_3[463]},
      {stage0_4[150]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[45],stage1_5[96],stage1_4[165],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[464], stage0_3[465], stage0_3[466], stage0_3[467], stage0_3[468]},
      {stage0_4[151]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[46],stage1_5[97],stage1_4[166],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[469], stage0_3[470], stage0_3[471], stage0_3[472], stage0_3[473]},
      {stage0_4[152]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[47],stage1_5[98],stage1_4[167],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[474], stage0_3[475], stage0_3[476], stage0_3[477], stage0_3[478]},
      {stage0_4[153]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[48],stage1_5[99],stage1_4[168],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[479], stage0_3[480], stage0_3[481], stage0_3[482], stage0_3[483]},
      {stage0_4[154]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[49],stage1_5[100],stage1_4[169],stage1_3[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[29],stage1_6[50],stage1_5[101],stage1_4[170]}
   );
   gpc606_5 gpc187 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[30],stage1_6[51],stage1_5[102],stage1_4[171]}
   );
   gpc606_5 gpc188 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[31],stage1_6[52],stage1_5[103],stage1_4[172]}
   );
   gpc606_5 gpc189 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[32],stage1_6[53],stage1_5[104],stage1_4[173]}
   );
   gpc606_5 gpc190 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[33],stage1_6[54],stage1_5[105],stage1_4[174]}
   );
   gpc606_5 gpc191 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[34],stage1_6[55],stage1_5[106],stage1_4[175]}
   );
   gpc606_5 gpc192 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[35],stage1_6[56],stage1_5[107],stage1_4[176]}
   );
   gpc606_5 gpc193 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[36],stage1_6[57],stage1_5[108],stage1_4[177]}
   );
   gpc606_5 gpc194 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[37],stage1_6[58],stage1_5[109],stage1_4[178]}
   );
   gpc606_5 gpc195 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[38],stage1_6[59],stage1_5[110],stage1_4[179]}
   );
   gpc606_5 gpc196 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[39],stage1_6[60],stage1_5[111],stage1_4[180]}
   );
   gpc606_5 gpc197 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[40],stage1_6[61],stage1_5[112],stage1_4[181]}
   );
   gpc606_5 gpc198 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[41],stage1_6[62],stage1_5[113],stage1_4[182]}
   );
   gpc606_5 gpc199 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[42],stage1_6[63],stage1_5[114],stage1_4[183]}
   );
   gpc606_5 gpc200 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[43],stage1_6[64],stage1_5[115],stage1_4[184]}
   );
   gpc606_5 gpc201 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[44],stage1_6[65],stage1_5[116],stage1_4[185]}
   );
   gpc606_5 gpc202 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[45],stage1_6[66],stage1_5[117],stage1_4[186]}
   );
   gpc606_5 gpc203 (
      {stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[46],stage1_6[67],stage1_5[118],stage1_4[187]}
   );
   gpc606_5 gpc204 (
      {stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[47],stage1_6[68],stage1_5[119],stage1_4[188]}
   );
   gpc606_5 gpc205 (
      {stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[48],stage1_6[69],stage1_5[120],stage1_4[189]}
   );
   gpc606_5 gpc206 (
      {stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[49],stage1_6[70],stage1_5[121],stage1_4[190]}
   );
   gpc606_5 gpc207 (
      {stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[50],stage1_6[71],stage1_5[122],stage1_4[191]}
   );
   gpc606_5 gpc208 (
      {stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[51],stage1_6[72],stage1_5[123],stage1_4[192]}
   );
   gpc606_5 gpc209 (
      {stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[52],stage1_6[73],stage1_5[124],stage1_4[193]}
   );
   gpc606_5 gpc210 (
      {stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[53],stage1_6[74],stage1_5[125],stage1_4[194]}
   );
   gpc606_5 gpc211 (
      {stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[54],stage1_6[75],stage1_5[126],stage1_4[195]}
   );
   gpc606_5 gpc212 (
      {stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[55],stage1_6[76],stage1_5[127],stage1_4[196]}
   );
   gpc606_5 gpc213 (
      {stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[56],stage1_6[77],stage1_5[128],stage1_4[197]}
   );
   gpc606_5 gpc214 (
      {stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[57],stage1_6[78],stage1_5[129],stage1_4[198]}
   );
   gpc606_5 gpc215 (
      {stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[58],stage1_6[79],stage1_5[130],stage1_4[199]}
   );
   gpc606_5 gpc216 (
      {stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[59],stage1_6[80],stage1_5[131],stage1_4[200]}
   );
   gpc606_5 gpc217 (
      {stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[60],stage1_6[81],stage1_5[132],stage1_4[201]}
   );
   gpc606_5 gpc218 (
      {stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[61],stage1_6[82],stage1_5[133],stage1_4[202]}
   );
   gpc606_5 gpc219 (
      {stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[62],stage1_6[83],stage1_5[134],stage1_4[203]}
   );
   gpc606_5 gpc220 (
      {stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[63],stage1_6[84],stage1_5[135],stage1_4[204]}
   );
   gpc606_5 gpc221 (
      {stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[64],stage1_6[85],stage1_5[136],stage1_4[205]}
   );
   gpc606_5 gpc222 (
      {stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[65],stage1_6[86],stage1_5[137],stage1_4[206]}
   );
   gpc606_5 gpc223 (
      {stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[66],stage1_6[87],stage1_5[138],stage1_4[207]}
   );
   gpc606_5 gpc224 (
      {stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[67],stage1_6[88],stage1_5[139],stage1_4[208]}
   );
   gpc606_5 gpc225 (
      {stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[68],stage1_6[89],stage1_5[140],stage1_4[209]}
   );
   gpc606_5 gpc226 (
      {stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[69],stage1_6[90],stage1_5[141],stage1_4[210]}
   );
   gpc606_5 gpc227 (
      {stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[70],stage1_6[91],stage1_5[142],stage1_4[211]}
   );
   gpc606_5 gpc228 (
      {stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[71],stage1_6[92],stage1_5[143],stage1_4[212]}
   );
   gpc606_5 gpc229 (
      {stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[72],stage1_6[93],stage1_5[144],stage1_4[213]}
   );
   gpc606_5 gpc230 (
      {stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[73],stage1_6[94],stage1_5[145],stage1_4[214]}
   );
   gpc606_5 gpc231 (
      {stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[74],stage1_6[95],stage1_5[146],stage1_4[215]}
   );
   gpc606_5 gpc232 (
      {stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[75],stage1_6[96],stage1_5[147],stage1_4[216]}
   );
   gpc606_5 gpc233 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[76],stage1_6[97],stage1_5[148],stage1_4[217]}
   );
   gpc606_5 gpc234 (
      {stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[77],stage1_6[98],stage1_5[149],stage1_4[218]}
   );
   gpc606_5 gpc235 (
      {stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[78],stage1_6[99],stage1_5[150],stage1_4[219]}
   );
   gpc606_5 gpc236 (
      {stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[79],stage1_6[100],stage1_5[151],stage1_4[220]}
   );
   gpc606_5 gpc237 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[80],stage1_6[101],stage1_5[152],stage1_4[221]}
   );
   gpc606_5 gpc238 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[81],stage1_6[102],stage1_5[153],stage1_4[222]}
   );
   gpc606_5 gpc239 (
      {stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[82],stage1_6[103],stage1_5[154],stage1_4[223]}
   );
   gpc606_5 gpc240 (
      {stage0_4[479], stage0_4[480], stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[83],stage1_6[104],stage1_5[155],stage1_4[224]}
   );
   gpc606_5 gpc241 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[84],stage1_6[105],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[85],stage1_6[106],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[86],stage1_6[107],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[87],stage1_6[108],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[88],stage1_6[109],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[89],stage1_6[110],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[90],stage1_6[111],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[91],stage1_6[112],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[92],stage1_6[113],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[93],stage1_6[114],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[94],stage1_6[115],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[95],stage1_6[116],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[96],stage1_6[117],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[97],stage1_6[118],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[98],stage1_6[119],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[99],stage1_6[120],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[100],stage1_6[121],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[101],stage1_6[122],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[102],stage1_6[123],stage1_5[174]}
   );
   gpc606_5 gpc260 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[103],stage1_6[124],stage1_5[175]}
   );
   gpc606_5 gpc261 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[104],stage1_6[125],stage1_5[176]}
   );
   gpc606_5 gpc262 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[105],stage1_6[126],stage1_5[177]}
   );
   gpc606_5 gpc263 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[106],stage1_6[127],stage1_5[178]}
   );
   gpc606_5 gpc264 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[107],stage1_6[128],stage1_5[179]}
   );
   gpc606_5 gpc265 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[108],stage1_6[129],stage1_5[180]}
   );
   gpc606_5 gpc266 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[109],stage1_6[130],stage1_5[181]}
   );
   gpc606_5 gpc267 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[110],stage1_6[131],stage1_5[182]}
   );
   gpc606_5 gpc268 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[111],stage1_6[132],stage1_5[183]}
   );
   gpc606_5 gpc269 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[112],stage1_6[133],stage1_5[184]}
   );
   gpc606_5 gpc270 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[113],stage1_6[134],stage1_5[185]}
   );
   gpc606_5 gpc271 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[114],stage1_6[135],stage1_5[186]}
   );
   gpc606_5 gpc272 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[115],stage1_6[136],stage1_5[187]}
   );
   gpc606_5 gpc273 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[116],stage1_6[137],stage1_5[188]}
   );
   gpc606_5 gpc274 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[117],stage1_6[138],stage1_5[189]}
   );
   gpc606_5 gpc275 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[118],stage1_6[139],stage1_5[190]}
   );
   gpc606_5 gpc276 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[119],stage1_6[140],stage1_5[191]}
   );
   gpc606_5 gpc277 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[120],stage1_6[141],stage1_5[192]}
   );
   gpc606_5 gpc278 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[121],stage1_6[142],stage1_5[193]}
   );
   gpc606_5 gpc279 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[122],stage1_6[143],stage1_5[194]}
   );
   gpc606_5 gpc280 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[123],stage1_6[144],stage1_5[195]}
   );
   gpc606_5 gpc281 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[124],stage1_6[145],stage1_5[196]}
   );
   gpc606_5 gpc282 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[125],stage1_6[146],stage1_5[197]}
   );
   gpc606_5 gpc283 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[126],stage1_6[147],stage1_5[198]}
   );
   gpc606_5 gpc284 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[127],stage1_6[148],stage1_5[199]}
   );
   gpc606_5 gpc285 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[128],stage1_6[149],stage1_5[200]}
   );
   gpc606_5 gpc286 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[129],stage1_6[150],stage1_5[201]}
   );
   gpc606_5 gpc287 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[130],stage1_6[151],stage1_5[202]}
   );
   gpc606_5 gpc288 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[131],stage1_6[152],stage1_5[203]}
   );
   gpc606_5 gpc289 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[132],stage1_6[153],stage1_5[204]}
   );
   gpc606_5 gpc290 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[133],stage1_6[154],stage1_5[205]}
   );
   gpc615_5 gpc291 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[105],stage1_7[134],stage1_6[155]}
   );
   gpc615_5 gpc292 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[106],stage1_7[135],stage1_6[156]}
   );
   gpc615_5 gpc293 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[107],stage1_7[136],stage1_6[157]}
   );
   gpc615_5 gpc294 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[108],stage1_7[137],stage1_6[158]}
   );
   gpc615_5 gpc295 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[109],stage1_7[138],stage1_6[159]}
   );
   gpc615_5 gpc296 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[110],stage1_7[139],stage1_6[160]}
   );
   gpc615_5 gpc297 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[111],stage1_7[140],stage1_6[161]}
   );
   gpc615_5 gpc298 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[112],stage1_7[141],stage1_6[162]}
   );
   gpc615_5 gpc299 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[113],stage1_7[142],stage1_6[163]}
   );
   gpc615_5 gpc300 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[114],stage1_7[143],stage1_6[164]}
   );
   gpc615_5 gpc301 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[115],stage1_7[144],stage1_6[165]}
   );
   gpc615_5 gpc302 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[116],stage1_7[145],stage1_6[166]}
   );
   gpc615_5 gpc303 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[117],stage1_7[146],stage1_6[167]}
   );
   gpc615_5 gpc304 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[118],stage1_7[147],stage1_6[168]}
   );
   gpc615_5 gpc305 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[119],stage1_7[148],stage1_6[169]}
   );
   gpc615_5 gpc306 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[120],stage1_7[149],stage1_6[170]}
   );
   gpc615_5 gpc307 (
      {stage0_7[316], stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320]},
      {stage0_8[96]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[16],stage1_9[66],stage1_8[121],stage1_7[150]}
   );
   gpc615_5 gpc308 (
      {stage0_7[321], stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325]},
      {stage0_8[97]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[17],stage1_9[67],stage1_8[122],stage1_7[151]}
   );
   gpc615_5 gpc309 (
      {stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330]},
      {stage0_8[98]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[18],stage1_9[68],stage1_8[123],stage1_7[152]}
   );
   gpc615_5 gpc310 (
      {stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage0_8[99]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[19],stage1_9[69],stage1_8[124],stage1_7[153]}
   );
   gpc615_5 gpc311 (
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340]},
      {stage0_8[100]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[20],stage1_9[70],stage1_8[125],stage1_7[154]}
   );
   gpc615_5 gpc312 (
      {stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345]},
      {stage0_8[101]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[21],stage1_9[71],stage1_8[126],stage1_7[155]}
   );
   gpc615_5 gpc313 (
      {stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350]},
      {stage0_8[102]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[22],stage1_9[72],stage1_8[127],stage1_7[156]}
   );
   gpc615_5 gpc314 (
      {stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355]},
      {stage0_8[103]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[23],stage1_9[73],stage1_8[128],stage1_7[157]}
   );
   gpc615_5 gpc315 (
      {stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360]},
      {stage0_8[104]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[24],stage1_9[74],stage1_8[129],stage1_7[158]}
   );
   gpc615_5 gpc316 (
      {stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage0_8[105]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[25],stage1_9[75],stage1_8[130],stage1_7[159]}
   );
   gpc615_5 gpc317 (
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_8[106]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[26],stage1_9[76],stage1_8[131],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375]},
      {stage0_8[107]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[27],stage1_9[77],stage1_8[132],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380]},
      {stage0_8[108]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[28],stage1_9[78],stage1_8[133],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385]},
      {stage0_8[109]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[29],stage1_9[79],stage1_8[134],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390]},
      {stage0_8[110]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[30],stage1_9[80],stage1_8[135],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage0_8[111]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[31],stage1_9[81],stage1_8[136],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_8[112]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[32],stage1_9[82],stage1_8[137],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405]},
      {stage0_8[113]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[33],stage1_9[83],stage1_8[138],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410]},
      {stage0_8[114]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[34],stage1_9[84],stage1_8[139],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415]},
      {stage0_8[115]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[35],stage1_9[85],stage1_8[140],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420]},
      {stage0_8[116]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[36],stage1_9[86],stage1_8[141],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage0_8[117]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[37],stage1_9[87],stage1_8[142],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_8[118]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[38],stage1_9[88],stage1_8[143],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435]},
      {stage0_8[119]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[39],stage1_9[89],stage1_8[144],stage1_7[173]}
   );
   gpc606_5 gpc331 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[24],stage1_10[40],stage1_9[90],stage1_8[145]}
   );
   gpc606_5 gpc332 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[25],stage1_10[41],stage1_9[91],stage1_8[146]}
   );
   gpc606_5 gpc333 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[26],stage1_10[42],stage1_9[92],stage1_8[147]}
   );
   gpc606_5 gpc334 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[27],stage1_10[43],stage1_9[93],stage1_8[148]}
   );
   gpc606_5 gpc335 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[28],stage1_10[44],stage1_9[94],stage1_8[149]}
   );
   gpc606_5 gpc336 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[29],stage1_10[45],stage1_9[95],stage1_8[150]}
   );
   gpc606_5 gpc337 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[30],stage1_10[46],stage1_9[96],stage1_8[151]}
   );
   gpc606_5 gpc338 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[31],stage1_10[47],stage1_9[97],stage1_8[152]}
   );
   gpc606_5 gpc339 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[32],stage1_10[48],stage1_9[98],stage1_8[153]}
   );
   gpc606_5 gpc340 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[33],stage1_10[49],stage1_9[99],stage1_8[154]}
   );
   gpc606_5 gpc341 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[34],stage1_10[50],stage1_9[100],stage1_8[155]}
   );
   gpc606_5 gpc342 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[35],stage1_10[51],stage1_9[101],stage1_8[156]}
   );
   gpc606_5 gpc343 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[36],stage1_10[52],stage1_9[102],stage1_8[157]}
   );
   gpc606_5 gpc344 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[37],stage1_10[53],stage1_9[103],stage1_8[158]}
   );
   gpc606_5 gpc345 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[38],stage1_10[54],stage1_9[104],stage1_8[159]}
   );
   gpc606_5 gpc346 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[39],stage1_10[55],stage1_9[105],stage1_8[160]}
   );
   gpc606_5 gpc347 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[40],stage1_10[56],stage1_9[106],stage1_8[161]}
   );
   gpc606_5 gpc348 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[41],stage1_10[57],stage1_9[107],stage1_8[162]}
   );
   gpc606_5 gpc349 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[42],stage1_10[58],stage1_9[108],stage1_8[163]}
   );
   gpc606_5 gpc350 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[43],stage1_10[59],stage1_9[109],stage1_8[164]}
   );
   gpc606_5 gpc351 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[44],stage1_10[60],stage1_9[110],stage1_8[165]}
   );
   gpc606_5 gpc352 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[45],stage1_10[61],stage1_9[111],stage1_8[166]}
   );
   gpc606_5 gpc353 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[46],stage1_10[62],stage1_9[112],stage1_8[167]}
   );
   gpc606_5 gpc354 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[47],stage1_10[63],stage1_9[113],stage1_8[168]}
   );
   gpc606_5 gpc355 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[48],stage1_10[64],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc356 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[49],stage1_10[65],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc357 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[50],stage1_10[66],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc358 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[51],stage1_10[67],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc359 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[52],stage1_10[68],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc360 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[53],stage1_10[69],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc361 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[54],stage1_10[70],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc362 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[55],stage1_10[71],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc363 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[56],stage1_10[72],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc364 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[57],stage1_10[73],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc365 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[58],stage1_10[74],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc366 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[59],stage1_10[75],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc367 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[60],stage1_10[76],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc368 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[61],stage1_10[77],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc369 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[62],stage1_10[78],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc370 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[63],stage1_10[79],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc371 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[64],stage1_10[80],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc372 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[65],stage1_10[81],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc373 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[66],stage1_10[82],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc374 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[67],stage1_10[83],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc375 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[68],stage1_10[84],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc376 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[69],stage1_10[85],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc377 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[70],stage1_10[86],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc378 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[71],stage1_10[87],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc379 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[72],stage1_10[88],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc380 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[73],stage1_10[89],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc381 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[74],stage1_10[90],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc382 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[75],stage1_10[91],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc383 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[76],stage1_10[92],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc384 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[77],stage1_10[93],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc385 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[78],stage1_10[94],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc386 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[79],stage1_10[95],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc387 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[80],stage1_10[96],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc388 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[81],stage1_10[97],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc389 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[82],stage1_10[98],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc390 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[83],stage1_10[99],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc391 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[84],stage1_10[100],stage1_9[150],stage1_8[205]}
   );
   gpc117_4 gpc392 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[366]},
      {stage0_11[0]},
      {stage1_12[61],stage1_11[85],stage1_10[101],stage1_9[151]}
   );
   gpc117_4 gpc393 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156], stage0_9[157]},
      {stage0_10[367]},
      {stage0_11[1]},
      {stage1_12[62],stage1_11[86],stage1_10[102],stage1_9[152]}
   );
   gpc117_4 gpc394 (
      {stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164]},
      {stage0_10[368]},
      {stage0_11[2]},
      {stage1_12[63],stage1_11[87],stage1_10[103],stage1_9[153]}
   );
   gpc117_4 gpc395 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171]},
      {stage0_10[369]},
      {stage0_11[3]},
      {stage1_12[64],stage1_11[88],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177]},
      {stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9]},
      {stage1_13[0],stage1_12[65],stage1_11[89],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183]},
      {stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15]},
      {stage1_13[1],stage1_12[66],stage1_11[90],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189]},
      {stage0_11[16], stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21]},
      {stage1_13[2],stage1_12[67],stage1_11[91],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage1_13[3],stage1_12[68],stage1_11[92],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201]},
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33]},
      {stage1_13[4],stage1_12[69],stage1_11[93],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207]},
      {stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39]},
      {stage1_13[5],stage1_12[70],stage1_11[94],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213]},
      {stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45]},
      {stage1_13[6],stage1_12[71],stage1_11[95],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_11[46], stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51]},
      {stage1_13[7],stage1_12[72],stage1_11[96],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_11[52], stage0_11[53], stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57]},
      {stage1_13[8],stage1_12[73],stage1_11[97],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231]},
      {stage0_11[58], stage0_11[59], stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63]},
      {stage1_13[9],stage1_12[74],stage1_11[98],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237]},
      {stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69]},
      {stage1_13[10],stage1_12[75],stage1_11[99],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243]},
      {stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75]},
      {stage1_13[11],stage1_12[76],stage1_11[100],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249]},
      {stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81]},
      {stage1_13[12],stage1_12[77],stage1_11[101],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87]},
      {stage1_13[13],stage1_12[78],stage1_11[102],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261]},
      {stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93]},
      {stage1_13[14],stage1_12[79],stage1_11[103],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267]},
      {stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99]},
      {stage1_13[15],stage1_12[80],stage1_11[104],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273]},
      {stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105]},
      {stage1_13[16],stage1_12[81],stage1_11[105],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279]},
      {stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111]},
      {stage1_13[17],stage1_12[82],stage1_11[106],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117]},
      {stage1_13[18],stage1_12[83],stage1_11[107],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291]},
      {stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123]},
      {stage1_13[19],stage1_12[84],stage1_11[108],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297]},
      {stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage1_13[20],stage1_12[85],stage1_11[109],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303]},
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135]},
      {stage1_13[21],stage1_12[86],stage1_11[110],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309]},
      {stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141]},
      {stage1_13[22],stage1_12[87],stage1_11[111],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_11[142], stage0_11[143], stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147]},
      {stage1_13[23],stage1_12[88],stage1_11[112],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321]},
      {stage0_11[148], stage0_11[149], stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153]},
      {stage1_13[24],stage1_12[89],stage1_11[113],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327]},
      {stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage1_13[25],stage1_12[90],stage1_11[114],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333]},
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165]},
      {stage1_13[26],stage1_12[91],stage1_11[115],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339]},
      {stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171]},
      {stage1_13[27],stage1_12[92],stage1_11[116],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_11[172], stage0_11[173], stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177]},
      {stage1_13[28],stage1_12[93],stage1_11[117],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351]},
      {stage0_11[178], stage0_11[179], stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183]},
      {stage1_13[29],stage1_12[94],stage1_11[118],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357]},
      {stage0_11[184], stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage1_13[30],stage1_12[95],stage1_11[119],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363]},
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195]},
      {stage1_13[31],stage1_12[96],stage1_11[120],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369]},
      {stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201]},
      {stage1_13[32],stage1_12[97],stage1_11[121],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_11[202], stage0_11[203], stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207]},
      {stage1_13[33],stage1_12[98],stage1_11[122],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381]},
      {stage0_11[208], stage0_11[209], stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213]},
      {stage1_13[34],stage1_12[99],stage1_11[123],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387]},
      {stage0_11[214], stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage1_13[35],stage1_12[100],stage1_11[124],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393]},
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225]},
      {stage1_13[36],stage1_12[101],stage1_11[125],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399]},
      {stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231]},
      {stage1_13[37],stage1_12[102],stage1_11[126],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_11[232], stage0_11[233], stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237]},
      {stage1_13[38],stage1_12[103],stage1_11[127],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411]},
      {stage0_11[238], stage0_11[239], stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243]},
      {stage1_13[39],stage1_12[104],stage1_11[128],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417]},
      {stage0_11[244], stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage1_13[40],stage1_12[105],stage1_11[129],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc437 (
      {stage0_9[418], stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255]},
      {stage1_13[41],stage1_12[106],stage1_11[130],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc438 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429]},
      {stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261]},
      {stage1_13[42],stage1_12[107],stage1_11[131],stage1_10[147],stage1_9[197]}
   );
   gpc606_5 gpc439 (
      {stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_11[262], stage0_11[263], stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267]},
      {stage1_13[43],stage1_12[108],stage1_11[132],stage1_10[148],stage1_9[198]}
   );
   gpc606_5 gpc440 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441]},
      {stage0_11[268], stage0_11[269], stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273]},
      {stage1_13[44],stage1_12[109],stage1_11[133],stage1_10[149],stage1_9[199]}
   );
   gpc606_5 gpc441 (
      {stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447]},
      {stage0_11[274], stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage1_13[45],stage1_12[110],stage1_11[134],stage1_10[150],stage1_9[200]}
   );
   gpc606_5 gpc442 (
      {stage0_9[448], stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285]},
      {stage1_13[46],stage1_12[111],stage1_11[135],stage1_10[151],stage1_9[201]}
   );
   gpc606_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459]},
      {stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291]},
      {stage1_13[47],stage1_12[112],stage1_11[136],stage1_10[152],stage1_9[202]}
   );
   gpc606_5 gpc444 (
      {stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_11[292], stage0_11[293], stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297]},
      {stage1_13[48],stage1_12[113],stage1_11[137],stage1_10[153],stage1_9[203]}
   );
   gpc606_5 gpc445 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471]},
      {stage0_11[298], stage0_11[299], stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303]},
      {stage1_13[49],stage1_12[114],stage1_11[138],stage1_10[154],stage1_9[204]}
   );
   gpc606_5 gpc446 (
      {stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477]},
      {stage0_11[304], stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage1_13[50],stage1_12[115],stage1_11[139],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc447 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374]},
      {stage0_11[310]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[51],stage1_12[116],stage1_11[140],stage1_10[156]}
   );
   gpc615_5 gpc448 (
      {stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379]},
      {stage0_11[311]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[52],stage1_12[117],stage1_11[141],stage1_10[157]}
   );
   gpc615_5 gpc449 (
      {stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383], stage0_10[384]},
      {stage0_11[312]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[53],stage1_12[118],stage1_11[142],stage1_10[158]}
   );
   gpc615_5 gpc450 (
      {stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage0_11[313]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[54],stage1_12[119],stage1_11[143],stage1_10[159]}
   );
   gpc615_5 gpc451 (
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394]},
      {stage0_11[314]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[55],stage1_12[120],stage1_11[144],stage1_10[160]}
   );
   gpc615_5 gpc452 (
      {stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_11[315]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[56],stage1_12[121],stage1_11[145],stage1_10[161]}
   );
   gpc615_5 gpc453 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404]},
      {stage0_11[316]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[57],stage1_12[122],stage1_11[146],stage1_10[162]}
   );
   gpc615_5 gpc454 (
      {stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409]},
      {stage0_11[317]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[58],stage1_12[123],stage1_11[147],stage1_10[163]}
   );
   gpc615_5 gpc455 (
      {stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413], stage0_10[414]},
      {stage0_11[318]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[59],stage1_12[124],stage1_11[148],stage1_10[164]}
   );
   gpc615_5 gpc456 (
      {stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage0_11[319]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[60],stage1_12[125],stage1_11[149],stage1_10[165]}
   );
   gpc615_5 gpc457 (
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424]},
      {stage0_11[320]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[61],stage1_12[126],stage1_11[150],stage1_10[166]}
   );
   gpc615_5 gpc458 (
      {stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429]},
      {stage0_11[321]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[62],stage1_12[127],stage1_11[151],stage1_10[167]}
   );
   gpc615_5 gpc459 (
      {stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433], stage0_10[434]},
      {stage0_11[322]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[63],stage1_12[128],stage1_11[152],stage1_10[168]}
   );
   gpc615_5 gpc460 (
      {stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438], stage0_10[439]},
      {stage0_11[323]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[64],stage1_12[129],stage1_11[153],stage1_10[169]}
   );
   gpc615_5 gpc461 (
      {stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443], stage0_10[444]},
      {stage0_11[324]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[65],stage1_12[130],stage1_11[154],stage1_10[170]}
   );
   gpc615_5 gpc462 (
      {stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage0_11[325]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[66],stage1_12[131],stage1_11[155],stage1_10[171]}
   );
   gpc615_5 gpc463 (
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454]},
      {stage0_11[326]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[67],stage1_12[132],stage1_11[156],stage1_10[172]}
   );
   gpc615_5 gpc464 (
      {stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459]},
      {stage0_11[327]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[68],stage1_12[133],stage1_11[157],stage1_10[173]}
   );
   gpc615_5 gpc465 (
      {stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463], stage0_10[464]},
      {stage0_11[328]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[69],stage1_12[134],stage1_11[158],stage1_10[174]}
   );
   gpc615_5 gpc466 (
      {stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468], stage0_10[469]},
      {stage0_11[329]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[70],stage1_12[135],stage1_11[159],stage1_10[175]}
   );
   gpc615_5 gpc467 (
      {stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473], stage0_10[474]},
      {stage0_11[330]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[71],stage1_12[136],stage1_11[160],stage1_10[176]}
   );
   gpc615_5 gpc468 (
      {stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage0_12[126]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[21],stage1_13[72],stage1_12[137],stage1_11[161]}
   );
   gpc615_5 gpc469 (
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340]},
      {stage0_12[127]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[22],stage1_13[73],stage1_12[138],stage1_11[162]}
   );
   gpc615_5 gpc470 (
      {stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345]},
      {stage0_12[128]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[23],stage1_13[74],stage1_12[139],stage1_11[163]}
   );
   gpc615_5 gpc471 (
      {stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350]},
      {stage0_12[129]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[24],stage1_13[75],stage1_12[140],stage1_11[164]}
   );
   gpc615_5 gpc472 (
      {stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355]},
      {stage0_12[130]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[25],stage1_13[76],stage1_12[141],stage1_11[165]}
   );
   gpc615_5 gpc473 (
      {stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360]},
      {stage0_12[131]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[26],stage1_13[77],stage1_12[142],stage1_11[166]}
   );
   gpc615_5 gpc474 (
      {stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage0_12[132]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[27],stage1_13[78],stage1_12[143],stage1_11[167]}
   );
   gpc615_5 gpc475 (
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370]},
      {stage0_12[133]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[28],stage1_13[79],stage1_12[144],stage1_11[168]}
   );
   gpc615_5 gpc476 (
      {stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375]},
      {stage0_12[134]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[29],stage1_13[80],stage1_12[145],stage1_11[169]}
   );
   gpc615_5 gpc477 (
      {stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379], stage0_11[380]},
      {stage0_12[135]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[30],stage1_13[81],stage1_12[146],stage1_11[170]}
   );
   gpc615_5 gpc478 (
      {stage0_11[381], stage0_11[382], stage0_11[383], stage0_11[384], stage0_11[385]},
      {stage0_12[136]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[31],stage1_13[82],stage1_12[147],stage1_11[171]}
   );
   gpc615_5 gpc479 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[137]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[32],stage1_13[83],stage1_12[148],stage1_11[172]}
   );
   gpc615_5 gpc480 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[138]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[33],stage1_13[84],stage1_12[149],stage1_11[173]}
   );
   gpc615_5 gpc481 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[139]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[34],stage1_13[85],stage1_12[150],stage1_11[174]}
   );
   gpc615_5 gpc482 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[140]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[35],stage1_13[86],stage1_12[151],stage1_11[175]}
   );
   gpc615_5 gpc483 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[141]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[36],stage1_13[87],stage1_12[152],stage1_11[176]}
   );
   gpc615_5 gpc484 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[142]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[37],stage1_13[88],stage1_12[153],stage1_11[177]}
   );
   gpc615_5 gpc485 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[143]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[38],stage1_13[89],stage1_12[154],stage1_11[178]}
   );
   gpc615_5 gpc486 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[144]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[39],stage1_13[90],stage1_12[155],stage1_11[179]}
   );
   gpc615_5 gpc487 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[145]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[40],stage1_13[91],stage1_12[156],stage1_11[180]}
   );
   gpc615_5 gpc488 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[146]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[41],stage1_13[92],stage1_12[157],stage1_11[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[147]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[42],stage1_13[93],stage1_12[158],stage1_11[182]}
   );
   gpc615_5 gpc490 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[148]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[43],stage1_13[94],stage1_12[159],stage1_11[183]}
   );
   gpc615_5 gpc491 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[149]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[44],stage1_13[95],stage1_12[160],stage1_11[184]}
   );
   gpc606_5 gpc492 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[24],stage1_14[45],stage1_13[96],stage1_12[161]}
   );
   gpc606_5 gpc493 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[25],stage1_14[46],stage1_13[97],stage1_12[162]}
   );
   gpc606_5 gpc494 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[26],stage1_14[47],stage1_13[98],stage1_12[163]}
   );
   gpc606_5 gpc495 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[27],stage1_14[48],stage1_13[99],stage1_12[164]}
   );
   gpc606_5 gpc496 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[28],stage1_14[49],stage1_13[100],stage1_12[165]}
   );
   gpc606_5 gpc497 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[29],stage1_14[50],stage1_13[101],stage1_12[166]}
   );
   gpc606_5 gpc498 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[30],stage1_14[51],stage1_13[102],stage1_12[167]}
   );
   gpc606_5 gpc499 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[31],stage1_14[52],stage1_13[103],stage1_12[168]}
   );
   gpc606_5 gpc500 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[32],stage1_14[53],stage1_13[104],stage1_12[169]}
   );
   gpc606_5 gpc501 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[33],stage1_14[54],stage1_13[105],stage1_12[170]}
   );
   gpc606_5 gpc502 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[34],stage1_14[55],stage1_13[106],stage1_12[171]}
   );
   gpc606_5 gpc503 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[35],stage1_14[56],stage1_13[107],stage1_12[172]}
   );
   gpc606_5 gpc504 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[36],stage1_14[57],stage1_13[108],stage1_12[173]}
   );
   gpc606_5 gpc505 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[37],stage1_14[58],stage1_13[109],stage1_12[174]}
   );
   gpc606_5 gpc506 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[38],stage1_14[59],stage1_13[110],stage1_12[175]}
   );
   gpc606_5 gpc507 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[39],stage1_14[60],stage1_13[111],stage1_12[176]}
   );
   gpc606_5 gpc508 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[40],stage1_14[61],stage1_13[112],stage1_12[177]}
   );
   gpc606_5 gpc509 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[41],stage1_14[62],stage1_13[113],stage1_12[178]}
   );
   gpc606_5 gpc510 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[42],stage1_14[63],stage1_13[114],stage1_12[179]}
   );
   gpc606_5 gpc511 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[43],stage1_14[64],stage1_13[115],stage1_12[180]}
   );
   gpc606_5 gpc512 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[44],stage1_14[65],stage1_13[116],stage1_12[181]}
   );
   gpc606_5 gpc513 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[45],stage1_14[66],stage1_13[117],stage1_12[182]}
   );
   gpc606_5 gpc514 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[46],stage1_14[67],stage1_13[118],stage1_12[183]}
   );
   gpc606_5 gpc515 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[47],stage1_14[68],stage1_13[119],stage1_12[184]}
   );
   gpc606_5 gpc516 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[48],stage1_14[69],stage1_13[120],stage1_12[185]}
   );
   gpc606_5 gpc517 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[49],stage1_14[70],stage1_13[121],stage1_12[186]}
   );
   gpc606_5 gpc518 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[50],stage1_14[71],stage1_13[122],stage1_12[187]}
   );
   gpc606_5 gpc519 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[51],stage1_14[72],stage1_13[123],stage1_12[188]}
   );
   gpc606_5 gpc520 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[52],stage1_14[73],stage1_13[124],stage1_12[189]}
   );
   gpc606_5 gpc521 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[53],stage1_14[74],stage1_13[125],stage1_12[190]}
   );
   gpc606_5 gpc522 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[54],stage1_14[75],stage1_13[126],stage1_12[191]}
   );
   gpc606_5 gpc523 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[55],stage1_14[76],stage1_13[127],stage1_12[192]}
   );
   gpc606_5 gpc524 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[56],stage1_14[77],stage1_13[128],stage1_12[193]}
   );
   gpc606_5 gpc525 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[57],stage1_14[78],stage1_13[129],stage1_12[194]}
   );
   gpc606_5 gpc526 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[58],stage1_14[79],stage1_13[130],stage1_12[195]}
   );
   gpc606_5 gpc527 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[59],stage1_14[80],stage1_13[131],stage1_12[196]}
   );
   gpc606_5 gpc528 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[60],stage1_14[81],stage1_13[132],stage1_12[197]}
   );
   gpc606_5 gpc529 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[61],stage1_14[82],stage1_13[133],stage1_12[198]}
   );
   gpc606_5 gpc530 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[62],stage1_14[83],stage1_13[134],stage1_12[199]}
   );
   gpc606_5 gpc531 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[63],stage1_14[84],stage1_13[135],stage1_12[200]}
   );
   gpc606_5 gpc532 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[64],stage1_14[85],stage1_13[136],stage1_12[201]}
   );
   gpc606_5 gpc533 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[65],stage1_14[86],stage1_13[137],stage1_12[202]}
   );
   gpc606_5 gpc534 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[66],stage1_14[87],stage1_13[138],stage1_12[203]}
   );
   gpc606_5 gpc535 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[43],stage1_15[67],stage1_14[88],stage1_13[139]}
   );
   gpc606_5 gpc536 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[44],stage1_15[68],stage1_14[89],stage1_13[140]}
   );
   gpc606_5 gpc537 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[45],stage1_15[69],stage1_14[90],stage1_13[141]}
   );
   gpc606_5 gpc538 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[46],stage1_15[70],stage1_14[91],stage1_13[142]}
   );
   gpc606_5 gpc539 (
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[47],stage1_15[71],stage1_14[92],stage1_13[143]}
   );
   gpc606_5 gpc540 (
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[48],stage1_15[72],stage1_14[93],stage1_13[144]}
   );
   gpc606_5 gpc541 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[49],stage1_15[73],stage1_14[94],stage1_13[145]}
   );
   gpc606_5 gpc542 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[50],stage1_15[74],stage1_14[95],stage1_13[146]}
   );
   gpc606_5 gpc543 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[51],stage1_15[75],stage1_14[96],stage1_13[147]}
   );
   gpc606_5 gpc544 (
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[52],stage1_15[76],stage1_14[97],stage1_13[148]}
   );
   gpc606_5 gpc545 (
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[53],stage1_15[77],stage1_14[98],stage1_13[149]}
   );
   gpc606_5 gpc546 (
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[54],stage1_15[78],stage1_14[99],stage1_13[150]}
   );
   gpc606_5 gpc547 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[55],stage1_15[79],stage1_14[100],stage1_13[151]}
   );
   gpc606_5 gpc548 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[56],stage1_15[80],stage1_14[101],stage1_13[152]}
   );
   gpc606_5 gpc549 (
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[57],stage1_15[81],stage1_14[102],stage1_13[153]}
   );
   gpc606_5 gpc550 (
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[58],stage1_15[82],stage1_14[103],stage1_13[154]}
   );
   gpc606_5 gpc551 (
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[59],stage1_15[83],stage1_14[104],stage1_13[155]}
   );
   gpc606_5 gpc552 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[60],stage1_15[84],stage1_14[105],stage1_13[156]}
   );
   gpc606_5 gpc553 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[61],stage1_15[85],stage1_14[106],stage1_13[157]}
   );
   gpc606_5 gpc554 (
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[62],stage1_15[86],stage1_14[107],stage1_13[158]}
   );
   gpc606_5 gpc555 (
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[63],stage1_15[87],stage1_14[108],stage1_13[159]}
   );
   gpc606_5 gpc556 (
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[64],stage1_15[88],stage1_14[109],stage1_13[160]}
   );
   gpc606_5 gpc557 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[65],stage1_15[89],stage1_14[110],stage1_13[161]}
   );
   gpc606_5 gpc558 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[66],stage1_15[90],stage1_14[111],stage1_13[162]}
   );
   gpc606_5 gpc559 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[67],stage1_15[91],stage1_14[112],stage1_13[163]}
   );
   gpc606_5 gpc560 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[68],stage1_15[92],stage1_14[113],stage1_13[164]}
   );
   gpc606_5 gpc561 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[69],stage1_15[93],stage1_14[114],stage1_13[165]}
   );
   gpc606_5 gpc562 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[70],stage1_15[94],stage1_14[115],stage1_13[166]}
   );
   gpc606_5 gpc563 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[71],stage1_15[95],stage1_14[116],stage1_13[167]}
   );
   gpc606_5 gpc564 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[72],stage1_15[96],stage1_14[117],stage1_13[168]}
   );
   gpc606_5 gpc565 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[73],stage1_15[97],stage1_14[118],stage1_13[169]}
   );
   gpc606_5 gpc566 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[74],stage1_15[98],stage1_14[119],stage1_13[170]}
   );
   gpc606_5 gpc567 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[75],stage1_15[99],stage1_14[120],stage1_13[171]}
   );
   gpc606_5 gpc568 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[76],stage1_15[100],stage1_14[121],stage1_13[172]}
   );
   gpc606_5 gpc569 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[77],stage1_15[101],stage1_14[122],stage1_13[173]}
   );
   gpc606_5 gpc570 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[78],stage1_15[102],stage1_14[123],stage1_13[174]}
   );
   gpc606_5 gpc571 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[79],stage1_15[103],stage1_14[124],stage1_13[175]}
   );
   gpc606_5 gpc572 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[80],stage1_15[104],stage1_14[125],stage1_13[176]}
   );
   gpc606_5 gpc573 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[81],stage1_15[105],stage1_14[126],stage1_13[177]}
   );
   gpc606_5 gpc574 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[82],stage1_15[106],stage1_14[127],stage1_13[178]}
   );
   gpc606_5 gpc575 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[83],stage1_15[107],stage1_14[128],stage1_13[179]}
   );
   gpc606_5 gpc576 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[84],stage1_15[108],stage1_14[129],stage1_13[180]}
   );
   gpc606_5 gpc577 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[85],stage1_15[109],stage1_14[130],stage1_13[181]}
   );
   gpc606_5 gpc578 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[86],stage1_15[110],stage1_14[131],stage1_13[182]}
   );
   gpc606_5 gpc579 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[87],stage1_15[111],stage1_14[132],stage1_13[183]}
   );
   gpc606_5 gpc580 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[88],stage1_15[112],stage1_14[133],stage1_13[184]}
   );
   gpc606_5 gpc581 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[89],stage1_15[113],stage1_14[134],stage1_13[185]}
   );
   gpc606_5 gpc582 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[90],stage1_15[114],stage1_14[135],stage1_13[186]}
   );
   gpc606_5 gpc583 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[91],stage1_15[115],stage1_14[136],stage1_13[187]}
   );
   gpc606_5 gpc584 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[92],stage1_15[116],stage1_14[137],stage1_13[188]}
   );
   gpc606_5 gpc585 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[93],stage1_15[117],stage1_14[138],stage1_13[189]}
   );
   gpc606_5 gpc586 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[94],stage1_15[118],stage1_14[139],stage1_13[190]}
   );
   gpc615_5 gpc587 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[258]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[95],stage1_15[119],stage1_14[140],stage1_13[191]}
   );
   gpc615_5 gpc588 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[259]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[96],stage1_15[120],stage1_14[141],stage1_13[192]}
   );
   gpc615_5 gpc589 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[260]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[97],stage1_15[121],stage1_14[142],stage1_13[193]}
   );
   gpc615_5 gpc590 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[261]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[98],stage1_15[122],stage1_14[143],stage1_13[194]}
   );
   gpc606_5 gpc591 (
      {stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[56],stage1_16[99],stage1_15[123],stage1_14[144]}
   );
   gpc606_5 gpc592 (
      {stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[57],stage1_16[100],stage1_15[124],stage1_14[145]}
   );
   gpc606_5 gpc593 (
      {stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[58],stage1_16[101],stage1_15[125],stage1_14[146]}
   );
   gpc606_5 gpc594 (
      {stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[59],stage1_16[102],stage1_15[126],stage1_14[147]}
   );
   gpc606_5 gpc595 (
      {stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[60],stage1_16[103],stage1_15[127],stage1_14[148]}
   );
   gpc606_5 gpc596 (
      {stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[61],stage1_16[104],stage1_15[128],stage1_14[149]}
   );
   gpc606_5 gpc597 (
      {stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[62],stage1_16[105],stage1_15[129],stage1_14[150]}
   );
   gpc615_5 gpc598 (
      {stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307], stage0_14[308]},
      {stage0_15[336]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[63],stage1_16[106],stage1_15[130],stage1_14[151]}
   );
   gpc615_5 gpc599 (
      {stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage0_15[337]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[64],stage1_16[107],stage1_15[131],stage1_14[152]}
   );
   gpc615_5 gpc600 (
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318]},
      {stage0_15[338]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[65],stage1_16[108],stage1_15[132],stage1_14[153]}
   );
   gpc615_5 gpc601 (
      {stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_15[339]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[66],stage1_16[109],stage1_15[133],stage1_14[154]}
   );
   gpc615_5 gpc602 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328]},
      {stage0_15[340]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[67],stage1_16[110],stage1_15[134],stage1_14[155]}
   );
   gpc615_5 gpc603 (
      {stage0_14[329], stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333]},
      {stage0_15[341]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[68],stage1_16[111],stage1_15[135],stage1_14[156]}
   );
   gpc615_5 gpc604 (
      {stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337], stage0_14[338]},
      {stage0_15[342]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[69],stage1_16[112],stage1_15[136],stage1_14[157]}
   );
   gpc615_5 gpc605 (
      {stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage0_15[343]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[70],stage1_16[113],stage1_15[137],stage1_14[158]}
   );
   gpc615_5 gpc606 (
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348]},
      {stage0_15[344]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[71],stage1_16[114],stage1_15[138],stage1_14[159]}
   );
   gpc615_5 gpc607 (
      {stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_16[96]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[16],stage1_17[72],stage1_16[115],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354]},
      {stage0_16[97]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[17],stage1_17[73],stage1_16[116],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage0_16[98]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[18],stage1_17[74],stage1_16[117],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364]},
      {stage0_16[99]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[19],stage1_17[75],stage1_16[118],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369]},
      {stage0_16[100]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[20],stage1_17[76],stage1_16[119],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374]},
      {stage0_16[101]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[21],stage1_17[77],stage1_16[120],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379]},
      {stage0_16[102]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[22],stage1_17[78],stage1_16[121],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384]},
      {stage0_16[103]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[23],stage1_17[79],stage1_16[122],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage0_16[104]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[24],stage1_17[80],stage1_16[123],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394]},
      {stage0_16[105]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[25],stage1_17[81],stage1_16[124],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399]},
      {stage0_16[106]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[26],stage1_17[82],stage1_16[125],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404]},
      {stage0_16[107]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[27],stage1_17[83],stage1_16[126],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409]},
      {stage0_16[108]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[28],stage1_17[84],stage1_16[127],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414]},
      {stage0_16[109]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[29],stage1_17[85],stage1_16[128],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage0_16[110]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[30],stage1_17[86],stage1_16[129],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424]},
      {stage0_16[111]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[31],stage1_17[87],stage1_16[130],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429]},
      {stage0_16[112]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[32],stage1_17[88],stage1_16[131],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434]},
      {stage0_16[113]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[33],stage1_17[89],stage1_16[132],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439]},
      {stage0_16[114]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[34],stage1_17[90],stage1_16[133],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444]},
      {stage0_16[115]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[35],stage1_17[91],stage1_16[134],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage0_16[116]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[36],stage1_17[92],stage1_16[135],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454]},
      {stage0_16[117]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[37],stage1_17[93],stage1_16[136],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459]},
      {stage0_16[118]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[38],stage1_17[94],stage1_16[137],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463], stage0_15[464]},
      {stage0_16[119]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[39],stage1_17[95],stage1_16[138],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468], stage0_15[469]},
      {stage0_16[120]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[40],stage1_17[96],stage1_16[139],stage1_15[163]}
   );
   gpc615_5 gpc632 (
      {stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473], stage0_15[474]},
      {stage0_16[121]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[41],stage1_17[97],stage1_16[140],stage1_15[164]}
   );
   gpc615_5 gpc633 (
      {stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage0_16[122]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[42],stage1_17[98],stage1_16[141],stage1_15[165]}
   );
   gpc606_5 gpc634 (
      {stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127], stage0_16[128]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[27],stage1_18[43],stage1_17[99],stage1_16[142]}
   );
   gpc606_5 gpc635 (
      {stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133], stage0_16[134]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[28],stage1_18[44],stage1_17[100],stage1_16[143]}
   );
   gpc606_5 gpc636 (
      {stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139], stage0_16[140]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[29],stage1_18[45],stage1_17[101],stage1_16[144]}
   );
   gpc606_5 gpc637 (
      {stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145], stage0_16[146]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[30],stage1_18[46],stage1_17[102],stage1_16[145]}
   );
   gpc606_5 gpc638 (
      {stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[31],stage1_18[47],stage1_17[103],stage1_16[146]}
   );
   gpc606_5 gpc639 (
      {stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[32],stage1_18[48],stage1_17[104],stage1_16[147]}
   );
   gpc606_5 gpc640 (
      {stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[33],stage1_18[49],stage1_17[105],stage1_16[148]}
   );
   gpc606_5 gpc641 (
      {stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[34],stage1_18[50],stage1_17[106],stage1_16[149]}
   );
   gpc606_5 gpc642 (
      {stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[35],stage1_18[51],stage1_17[107],stage1_16[150]}
   );
   gpc606_5 gpc643 (
      {stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[36],stage1_18[52],stage1_17[108],stage1_16[151]}
   );
   gpc606_5 gpc644 (
      {stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[37],stage1_18[53],stage1_17[109],stage1_16[152]}
   );
   gpc606_5 gpc645 (
      {stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[38],stage1_18[54],stage1_17[110],stage1_16[153]}
   );
   gpc606_5 gpc646 (
      {stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[39],stage1_18[55],stage1_17[111],stage1_16[154]}
   );
   gpc606_5 gpc647 (
      {stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[40],stage1_18[56],stage1_17[112],stage1_16[155]}
   );
   gpc606_5 gpc648 (
      {stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[41],stage1_18[57],stage1_17[113],stage1_16[156]}
   );
   gpc606_5 gpc649 (
      {stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[42],stage1_18[58],stage1_17[114],stage1_16[157]}
   );
   gpc606_5 gpc650 (
      {stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[43],stage1_18[59],stage1_17[115],stage1_16[158]}
   );
   gpc606_5 gpc651 (
      {stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[44],stage1_18[60],stage1_17[116],stage1_16[159]}
   );
   gpc606_5 gpc652 (
      {stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[45],stage1_18[61],stage1_17[117],stage1_16[160]}
   );
   gpc606_5 gpc653 (
      {stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[46],stage1_18[62],stage1_17[118],stage1_16[161]}
   );
   gpc606_5 gpc654 (
      {stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[47],stage1_18[63],stage1_17[119],stage1_16[162]}
   );
   gpc606_5 gpc655 (
      {stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[48],stage1_18[64],stage1_17[120],stage1_16[163]}
   );
   gpc606_5 gpc656 (
      {stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259], stage0_16[260]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[49],stage1_18[65],stage1_17[121],stage1_16[164]}
   );
   gpc606_5 gpc657 (
      {stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265], stage0_16[266]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[50],stage1_18[66],stage1_17[122],stage1_16[165]}
   );
   gpc606_5 gpc658 (
      {stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271], stage0_16[272]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[51],stage1_18[67],stage1_17[123],stage1_16[166]}
   );
   gpc606_5 gpc659 (
      {stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277], stage0_16[278]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[52],stage1_18[68],stage1_17[124],stage1_16[167]}
   );
   gpc606_5 gpc660 (
      {stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283], stage0_16[284]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[53],stage1_18[69],stage1_17[125],stage1_16[168]}
   );
   gpc606_5 gpc661 (
      {stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289], stage0_16[290]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[54],stage1_18[70],stage1_17[126],stage1_16[169]}
   );
   gpc606_5 gpc662 (
      {stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295], stage0_16[296]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[55],stage1_18[71],stage1_17[127],stage1_16[170]}
   );
   gpc606_5 gpc663 (
      {stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301], stage0_16[302]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[56],stage1_18[72],stage1_17[128],stage1_16[171]}
   );
   gpc606_5 gpc664 (
      {stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307], stage0_16[308]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[57],stage1_18[73],stage1_17[129],stage1_16[172]}
   );
   gpc606_5 gpc665 (
      {stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313], stage0_16[314]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[58],stage1_18[74],stage1_17[130],stage1_16[173]}
   );
   gpc606_5 gpc666 (
      {stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319], stage0_16[320]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[59],stage1_18[75],stage1_17[131],stage1_16[174]}
   );
   gpc606_5 gpc667 (
      {stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325], stage0_16[326]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[60],stage1_18[76],stage1_17[132],stage1_16[175]}
   );
   gpc606_5 gpc668 (
      {stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331], stage0_16[332]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[61],stage1_18[77],stage1_17[133],stage1_16[176]}
   );
   gpc606_5 gpc669 (
      {stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337], stage0_16[338]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[62],stage1_18[78],stage1_17[134],stage1_16[177]}
   );
   gpc606_5 gpc670 (
      {stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343], stage0_16[344]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[63],stage1_18[79],stage1_17[135],stage1_16[178]}
   );
   gpc606_5 gpc671 (
      {stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349], stage0_16[350]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[64],stage1_18[80],stage1_17[136],stage1_16[179]}
   );
   gpc606_5 gpc672 (
      {stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355], stage0_16[356]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[65],stage1_18[81],stage1_17[137],stage1_16[180]}
   );
   gpc606_5 gpc673 (
      {stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361], stage0_16[362]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[66],stage1_18[82],stage1_17[138],stage1_16[181]}
   );
   gpc606_5 gpc674 (
      {stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367], stage0_16[368]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[67],stage1_18[83],stage1_17[139],stage1_16[182]}
   );
   gpc606_5 gpc675 (
      {stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373], stage0_16[374]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[68],stage1_18[84],stage1_17[140],stage1_16[183]}
   );
   gpc606_5 gpc676 (
      {stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379], stage0_16[380]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[69],stage1_18[85],stage1_17[141],stage1_16[184]}
   );
   gpc606_5 gpc677 (
      {stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385], stage0_16[386]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[70],stage1_18[86],stage1_17[142],stage1_16[185]}
   );
   gpc606_5 gpc678 (
      {stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391], stage0_16[392]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[71],stage1_18[87],stage1_17[143],stage1_16[186]}
   );
   gpc606_5 gpc679 (
      {stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397], stage0_16[398]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[72],stage1_18[88],stage1_17[144],stage1_16[187]}
   );
   gpc606_5 gpc680 (
      {stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403], stage0_16[404]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[73],stage1_18[89],stage1_17[145],stage1_16[188]}
   );
   gpc606_5 gpc681 (
      {stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409], stage0_16[410]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[74],stage1_18[90],stage1_17[146],stage1_16[189]}
   );
   gpc606_5 gpc682 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[48],stage1_19[75],stage1_18[91],stage1_17[147]}
   );
   gpc606_5 gpc683 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[49],stage1_19[76],stage1_18[92],stage1_17[148]}
   );
   gpc606_5 gpc684 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[50],stage1_19[77],stage1_18[93],stage1_17[149]}
   );
   gpc606_5 gpc685 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[51],stage1_19[78],stage1_18[94],stage1_17[150]}
   );
   gpc606_5 gpc686 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[52],stage1_19[79],stage1_18[95],stage1_17[151]}
   );
   gpc606_5 gpc687 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[53],stage1_19[80],stage1_18[96],stage1_17[152]}
   );
   gpc606_5 gpc688 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[54],stage1_19[81],stage1_18[97],stage1_17[153]}
   );
   gpc606_5 gpc689 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[55],stage1_19[82],stage1_18[98],stage1_17[154]}
   );
   gpc606_5 gpc690 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[56],stage1_19[83],stage1_18[99],stage1_17[155]}
   );
   gpc606_5 gpc691 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[57],stage1_19[84],stage1_18[100],stage1_17[156]}
   );
   gpc606_5 gpc692 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[58],stage1_19[85],stage1_18[101],stage1_17[157]}
   );
   gpc606_5 gpc693 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[59],stage1_19[86],stage1_18[102],stage1_17[158]}
   );
   gpc606_5 gpc694 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[60],stage1_19[87],stage1_18[103],stage1_17[159]}
   );
   gpc606_5 gpc695 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[61],stage1_19[88],stage1_18[104],stage1_17[160]}
   );
   gpc606_5 gpc696 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[62],stage1_19[89],stage1_18[105],stage1_17[161]}
   );
   gpc606_5 gpc697 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[63],stage1_19[90],stage1_18[106],stage1_17[162]}
   );
   gpc606_5 gpc698 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[64],stage1_19[91],stage1_18[107],stage1_17[163]}
   );
   gpc606_5 gpc699 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[65],stage1_19[92],stage1_18[108],stage1_17[164]}
   );
   gpc606_5 gpc700 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[66],stage1_19[93],stage1_18[109],stage1_17[165]}
   );
   gpc606_5 gpc701 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[67],stage1_19[94],stage1_18[110],stage1_17[166]}
   );
   gpc606_5 gpc702 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[68],stage1_19[95],stage1_18[111],stage1_17[167]}
   );
   gpc606_5 gpc703 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[69],stage1_19[96],stage1_18[112],stage1_17[168]}
   );
   gpc606_5 gpc704 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[70],stage1_19[97],stage1_18[113],stage1_17[169]}
   );
   gpc606_5 gpc705 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[71],stage1_19[98],stage1_18[114],stage1_17[170]}
   );
   gpc606_5 gpc706 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[72],stage1_19[99],stage1_18[115],stage1_17[171]}
   );
   gpc606_5 gpc707 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[73],stage1_19[100],stage1_18[116],stage1_17[172]}
   );
   gpc606_5 gpc708 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[74],stage1_19[101],stage1_18[117],stage1_17[173]}
   );
   gpc606_5 gpc709 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[75],stage1_19[102],stage1_18[118],stage1_17[174]}
   );
   gpc606_5 gpc710 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[76],stage1_19[103],stage1_18[119],stage1_17[175]}
   );
   gpc606_5 gpc711 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[77],stage1_19[104],stage1_18[120],stage1_17[176]}
   );
   gpc606_5 gpc712 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[78],stage1_19[105],stage1_18[121],stage1_17[177]}
   );
   gpc606_5 gpc713 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[79],stage1_19[106],stage1_18[122],stage1_17[178]}
   );
   gpc606_5 gpc714 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[80],stage1_19[107],stage1_18[123],stage1_17[179]}
   );
   gpc606_5 gpc715 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[81],stage1_19[108],stage1_18[124],stage1_17[180]}
   );
   gpc606_5 gpc716 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[82],stage1_19[109],stage1_18[125],stage1_17[181]}
   );
   gpc606_5 gpc717 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[83],stage1_19[110],stage1_18[126],stage1_17[182]}
   );
   gpc606_5 gpc718 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[84],stage1_19[111],stage1_18[127],stage1_17[183]}
   );
   gpc606_5 gpc719 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[85],stage1_19[112],stage1_18[128],stage1_17[184]}
   );
   gpc606_5 gpc720 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[86],stage1_19[113],stage1_18[129],stage1_17[185]}
   );
   gpc606_5 gpc721 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[87],stage1_19[114],stage1_18[130],stage1_17[186]}
   );
   gpc606_5 gpc722 (
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[40],stage1_20[88],stage1_19[115],stage1_18[131]}
   );
   gpc606_5 gpc723 (
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[41],stage1_20[89],stage1_19[116],stage1_18[132]}
   );
   gpc606_5 gpc724 (
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[42],stage1_20[90],stage1_19[117],stage1_18[133]}
   );
   gpc606_5 gpc725 (
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[43],stage1_20[91],stage1_19[118],stage1_18[134]}
   );
   gpc615_5 gpc726 (
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316]},
      {stage0_19[240]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[44],stage1_20[92],stage1_19[119],stage1_18[135]}
   );
   gpc615_5 gpc727 (
      {stage0_18[317], stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321]},
      {stage0_19[241]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[45],stage1_20[93],stage1_19[120],stage1_18[136]}
   );
   gpc615_5 gpc728 (
      {stage0_18[322], stage0_18[323], stage0_18[324], stage0_18[325], stage0_18[326]},
      {stage0_19[242]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[46],stage1_20[94],stage1_19[121],stage1_18[137]}
   );
   gpc615_5 gpc729 (
      {stage0_18[327], stage0_18[328], stage0_18[329], stage0_18[330], stage0_18[331]},
      {stage0_19[243]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[47],stage1_20[95],stage1_19[122],stage1_18[138]}
   );
   gpc615_5 gpc730 (
      {stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335], stage0_18[336]},
      {stage0_19[244]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[48],stage1_20[96],stage1_19[123],stage1_18[139]}
   );
   gpc615_5 gpc731 (
      {stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage0_19[245]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[49],stage1_20[97],stage1_19[124],stage1_18[140]}
   );
   gpc615_5 gpc732 (
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346]},
      {stage0_19[246]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[50],stage1_20[98],stage1_19[125],stage1_18[141]}
   );
   gpc615_5 gpc733 (
      {stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351]},
      {stage0_19[247]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[51],stage1_20[99],stage1_19[126],stage1_18[142]}
   );
   gpc615_5 gpc734 (
      {stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355], stage0_18[356]},
      {stage0_19[248]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[52],stage1_20[100],stage1_19[127],stage1_18[143]}
   );
   gpc615_5 gpc735 (
      {stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360], stage0_18[361]},
      {stage0_19[249]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[53],stage1_20[101],stage1_19[128],stage1_18[144]}
   );
   gpc615_5 gpc736 (
      {stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365], stage0_18[366]},
      {stage0_19[250]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[54],stage1_20[102],stage1_19[129],stage1_18[145]}
   );
   gpc615_5 gpc737 (
      {stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage0_19[251]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[55],stage1_20[103],stage1_19[130],stage1_18[146]}
   );
   gpc615_5 gpc738 (
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376]},
      {stage0_19[252]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[56],stage1_20[104],stage1_19[131],stage1_18[147]}
   );
   gpc615_5 gpc739 (
      {stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381]},
      {stage0_19[253]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[57],stage1_20[105],stage1_19[132],stage1_18[148]}
   );
   gpc615_5 gpc740 (
      {stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385], stage0_18[386]},
      {stage0_19[254]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[58],stage1_20[106],stage1_19[133],stage1_18[149]}
   );
   gpc615_5 gpc741 (
      {stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390], stage0_18[391]},
      {stage0_19[255]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[59],stage1_20[107],stage1_19[134],stage1_18[150]}
   );
   gpc615_5 gpc742 (
      {stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395], stage0_18[396]},
      {stage0_19[256]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[60],stage1_20[108],stage1_19[135],stage1_18[151]}
   );
   gpc615_5 gpc743 (
      {stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage0_19[257]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[61],stage1_20[109],stage1_19[136],stage1_18[152]}
   );
   gpc615_5 gpc744 (
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406]},
      {stage0_19[258]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[62],stage1_20[110],stage1_19[137],stage1_18[153]}
   );
   gpc615_5 gpc745 (
      {stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411]},
      {stage0_19[259]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[63],stage1_20[111],stage1_19[138],stage1_18[154]}
   );
   gpc615_5 gpc746 (
      {stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415], stage0_18[416]},
      {stage0_19[260]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[64],stage1_20[112],stage1_19[139],stage1_18[155]}
   );
   gpc615_5 gpc747 (
      {stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420], stage0_18[421]},
      {stage0_19[261]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[65],stage1_20[113],stage1_19[140],stage1_18[156]}
   );
   gpc615_5 gpc748 (
      {stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425], stage0_18[426]},
      {stage0_19[262]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[66],stage1_20[114],stage1_19[141],stage1_18[157]}
   );
   gpc615_5 gpc749 (
      {stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430], stage0_18[431]},
      {stage0_19[263]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[67],stage1_20[115],stage1_19[142],stage1_18[158]}
   );
   gpc615_5 gpc750 (
      {stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435], stage0_18[436]},
      {stage0_19[264]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[68],stage1_20[116],stage1_19[143],stage1_18[159]}
   );
   gpc615_5 gpc751 (
      {stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440], stage0_18[441]},
      {stage0_19[265]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[69],stage1_20[117],stage1_19[144],stage1_18[160]}
   );
   gpc615_5 gpc752 (
      {stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445], stage0_18[446]},
      {stage0_19[266]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[70],stage1_20[118],stage1_19[145],stage1_18[161]}
   );
   gpc606_5 gpc753 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271], stage0_19[272]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[31],stage1_21[71],stage1_20[119],stage1_19[146]}
   );
   gpc606_5 gpc754 (
      {stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276], stage0_19[277], stage0_19[278]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[32],stage1_21[72],stage1_20[120],stage1_19[147]}
   );
   gpc606_5 gpc755 (
      {stage0_19[279], stage0_19[280], stage0_19[281], stage0_19[282], stage0_19[283], stage0_19[284]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[33],stage1_21[73],stage1_20[121],stage1_19[148]}
   );
   gpc606_5 gpc756 (
      {stage0_19[285], stage0_19[286], stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[34],stage1_21[74],stage1_20[122],stage1_19[149]}
   );
   gpc606_5 gpc757 (
      {stage0_19[291], stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[35],stage1_21[75],stage1_20[123],stage1_19[150]}
   );
   gpc615_5 gpc758 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[186]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[36],stage1_21[76],stage1_20[124],stage1_19[151]}
   );
   gpc615_5 gpc759 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[187]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[37],stage1_21[77],stage1_20[125],stage1_19[152]}
   );
   gpc615_5 gpc760 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[188]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[38],stage1_21[78],stage1_20[126],stage1_19[153]}
   );
   gpc615_5 gpc761 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[189]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[39],stage1_21[79],stage1_20[127],stage1_19[154]}
   );
   gpc615_5 gpc762 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[190]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[40],stage1_21[80],stage1_20[128],stage1_19[155]}
   );
   gpc615_5 gpc763 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[191]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[41],stage1_21[81],stage1_20[129],stage1_19[156]}
   );
   gpc615_5 gpc764 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[192]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[42],stage1_21[82],stage1_20[130],stage1_19[157]}
   );
   gpc615_5 gpc765 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[193]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[43],stage1_21[83],stage1_20[131],stage1_19[158]}
   );
   gpc615_5 gpc766 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[194]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[44],stage1_21[84],stage1_20[132],stage1_19[159]}
   );
   gpc615_5 gpc767 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[195]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[45],stage1_21[85],stage1_20[133],stage1_19[160]}
   );
   gpc606_5 gpc768 (
      {stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[15],stage1_22[46],stage1_21[86],stage1_20[134]}
   );
   gpc606_5 gpc769 (
      {stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[16],stage1_22[47],stage1_21[87],stage1_20[135]}
   );
   gpc606_5 gpc770 (
      {stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[17],stage1_22[48],stage1_21[88],stage1_20[136]}
   );
   gpc606_5 gpc771 (
      {stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[18],stage1_22[49],stage1_21[89],stage1_20[137]}
   );
   gpc606_5 gpc772 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[19],stage1_22[50],stage1_21[90],stage1_20[138]}
   );
   gpc606_5 gpc773 (
      {stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[20],stage1_22[51],stage1_21[91],stage1_20[139]}
   );
   gpc606_5 gpc774 (
      {stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[21],stage1_22[52],stage1_21[92],stage1_20[140]}
   );
   gpc606_5 gpc775 (
      {stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[22],stage1_22[53],stage1_21[93],stage1_20[141]}
   );
   gpc606_5 gpc776 (
      {stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[23],stage1_22[54],stage1_21[94],stage1_20[142]}
   );
   gpc606_5 gpc777 (
      {stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[24],stage1_22[55],stage1_21[95],stage1_20[143]}
   );
   gpc606_5 gpc778 (
      {stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[25],stage1_22[56],stage1_21[96],stage1_20[144]}
   );
   gpc606_5 gpc779 (
      {stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[26],stage1_22[57],stage1_21[97],stage1_20[145]}
   );
   gpc606_5 gpc780 (
      {stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[27],stage1_22[58],stage1_21[98],stage1_20[146]}
   );
   gpc606_5 gpc781 (
      {stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[28],stage1_22[59],stage1_21[99],stage1_20[147]}
   );
   gpc606_5 gpc782 (
      {stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[29],stage1_22[60],stage1_21[100],stage1_20[148]}
   );
   gpc606_5 gpc783 (
      {stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[30],stage1_22[61],stage1_21[101],stage1_20[149]}
   );
   gpc606_5 gpc784 (
      {stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[31],stage1_22[62],stage1_21[102],stage1_20[150]}
   );
   gpc606_5 gpc785 (
      {stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[32],stage1_22[63],stage1_21[103],stage1_20[151]}
   );
   gpc606_5 gpc786 (
      {stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[33],stage1_22[64],stage1_21[104],stage1_20[152]}
   );
   gpc606_5 gpc787 (
      {stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[34],stage1_22[65],stage1_21[105],stage1_20[153]}
   );
   gpc606_5 gpc788 (
      {stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[35],stage1_22[66],stage1_21[106],stage1_20[154]}
   );
   gpc606_5 gpc789 (
      {stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[36],stage1_22[67],stage1_21[107],stage1_20[155]}
   );
   gpc606_5 gpc790 (
      {stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[37],stage1_22[68],stage1_21[108],stage1_20[156]}
   );
   gpc606_5 gpc791 (
      {stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[38],stage1_22[69],stage1_21[109],stage1_20[157]}
   );
   gpc606_5 gpc792 (
      {stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[39],stage1_22[70],stage1_21[110],stage1_20[158]}
   );
   gpc606_5 gpc793 (
      {stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[40],stage1_22[71],stage1_21[111],stage1_20[159]}
   );
   gpc606_5 gpc794 (
      {stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[41],stage1_22[72],stage1_21[112],stage1_20[160]}
   );
   gpc606_5 gpc795 (
      {stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[42],stage1_22[73],stage1_21[113],stage1_20[161]}
   );
   gpc606_5 gpc796 (
      {stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[43],stage1_22[74],stage1_21[114],stage1_20[162]}
   );
   gpc606_5 gpc797 (
      {stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[44],stage1_22[75],stage1_21[115],stage1_20[163]}
   );
   gpc606_5 gpc798 (
      {stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[45],stage1_22[76],stage1_21[116],stage1_20[164]}
   );
   gpc606_5 gpc799 (
      {stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[46],stage1_22[77],stage1_21[117],stage1_20[165]}
   );
   gpc606_5 gpc800 (
      {stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[47],stage1_22[78],stage1_21[118],stage1_20[166]}
   );
   gpc606_5 gpc801 (
      {stage0_20[394], stage0_20[395], stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[48],stage1_22[79],stage1_21[119],stage1_20[167]}
   );
   gpc606_5 gpc802 (
      {stage0_20[400], stage0_20[401], stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[49],stage1_22[80],stage1_21[120],stage1_20[168]}
   );
   gpc606_5 gpc803 (
      {stage0_20[406], stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[50],stage1_22[81],stage1_21[121],stage1_20[169]}
   );
   gpc606_5 gpc804 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[51],stage1_22[82],stage1_21[122],stage1_20[170]}
   );
   gpc606_5 gpc805 (
      {stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[52],stage1_22[83],stage1_21[123],stage1_20[171]}
   );
   gpc606_5 gpc806 (
      {stage0_20[424], stage0_20[425], stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[53],stage1_22[84],stage1_21[124],stage1_20[172]}
   );
   gpc606_5 gpc807 (
      {stage0_20[430], stage0_20[431], stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[54],stage1_22[85],stage1_21[125],stage1_20[173]}
   );
   gpc606_5 gpc808 (
      {stage0_20[436], stage0_20[437], stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[55],stage1_22[86],stage1_21[126],stage1_20[174]}
   );
   gpc606_5 gpc809 (
      {stage0_20[442], stage0_20[443], stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[56],stage1_22[87],stage1_21[127],stage1_20[175]}
   );
   gpc606_5 gpc810 (
      {stage0_20[448], stage0_20[449], stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[57],stage1_22[88],stage1_21[128],stage1_20[176]}
   );
   gpc606_5 gpc811 (
      {stage0_20[454], stage0_20[455], stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[58],stage1_22[89],stage1_21[129],stage1_20[177]}
   );
   gpc606_5 gpc812 (
      {stage0_20[460], stage0_20[461], stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[59],stage1_22[90],stage1_21[130],stage1_20[178]}
   );
   gpc606_5 gpc813 (
      {stage0_20[466], stage0_20[467], stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[60],stage1_22[91],stage1_21[131],stage1_20[179]}
   );
   gpc606_5 gpc814 (
      {stage0_20[472], stage0_20[473], stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[61],stage1_22[92],stage1_21[132],stage1_20[180]}
   );
   gpc606_5 gpc815 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[47],stage1_23[62],stage1_22[93],stage1_21[133]}
   );
   gpc606_5 gpc816 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[48],stage1_23[63],stage1_22[94],stage1_21[134]}
   );
   gpc606_5 gpc817 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[49],stage1_23[64],stage1_22[95],stage1_21[135]}
   );
   gpc606_5 gpc818 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[50],stage1_23[65],stage1_22[96],stage1_21[136]}
   );
   gpc606_5 gpc819 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[51],stage1_23[66],stage1_22[97],stage1_21[137]}
   );
   gpc606_5 gpc820 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[52],stage1_23[67],stage1_22[98],stage1_21[138]}
   );
   gpc606_5 gpc821 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[53],stage1_23[68],stage1_22[99],stage1_21[139]}
   );
   gpc606_5 gpc822 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[54],stage1_23[69],stage1_22[100],stage1_21[140]}
   );
   gpc606_5 gpc823 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[55],stage1_23[70],stage1_22[101],stage1_21[141]}
   );
   gpc606_5 gpc824 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[56],stage1_23[71],stage1_22[102],stage1_21[142]}
   );
   gpc606_5 gpc825 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[57],stage1_23[72],stage1_22[103],stage1_21[143]}
   );
   gpc606_5 gpc826 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[58],stage1_23[73],stage1_22[104],stage1_21[144]}
   );
   gpc606_5 gpc827 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[59],stage1_23[74],stage1_22[105],stage1_21[145]}
   );
   gpc606_5 gpc828 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[60],stage1_23[75],stage1_22[106],stage1_21[146]}
   );
   gpc606_5 gpc829 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[61],stage1_23[76],stage1_22[107],stage1_21[147]}
   );
   gpc606_5 gpc830 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[62],stage1_23[77],stage1_22[108],stage1_21[148]}
   );
   gpc606_5 gpc831 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[63],stage1_23[78],stage1_22[109],stage1_21[149]}
   );
   gpc606_5 gpc832 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[64],stage1_23[79],stage1_22[110],stage1_21[150]}
   );
   gpc606_5 gpc833 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[65],stage1_23[80],stage1_22[111],stage1_21[151]}
   );
   gpc606_5 gpc834 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[66],stage1_23[81],stage1_22[112],stage1_21[152]}
   );
   gpc606_5 gpc835 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[67],stage1_23[82],stage1_22[113],stage1_21[153]}
   );
   gpc606_5 gpc836 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[68],stage1_23[83],stage1_22[114],stage1_21[154]}
   );
   gpc606_5 gpc837 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[69],stage1_23[84],stage1_22[115],stage1_21[155]}
   );
   gpc606_5 gpc838 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[70],stage1_23[85],stage1_22[116],stage1_21[156]}
   );
   gpc606_5 gpc839 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[71],stage1_23[86],stage1_22[117],stage1_21[157]}
   );
   gpc606_5 gpc840 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[72],stage1_23[87],stage1_22[118],stage1_21[158]}
   );
   gpc606_5 gpc841 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[73],stage1_23[88],stage1_22[119],stage1_21[159]}
   );
   gpc606_5 gpc842 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[74],stage1_23[89],stage1_22[120],stage1_21[160]}
   );
   gpc606_5 gpc843 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[75],stage1_23[90],stage1_22[121],stage1_21[161]}
   );
   gpc606_5 gpc844 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[76],stage1_23[91],stage1_22[122],stage1_21[162]}
   );
   gpc606_5 gpc845 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[77],stage1_23[92],stage1_22[123],stage1_21[163]}
   );
   gpc606_5 gpc846 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[78],stage1_23[93],stage1_22[124],stage1_21[164]}
   );
   gpc606_5 gpc847 (
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[79],stage1_23[94],stage1_22[125],stage1_21[165]}
   );
   gpc606_5 gpc848 (
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[80],stage1_23[95],stage1_22[126],stage1_21[166]}
   );
   gpc606_5 gpc849 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[81],stage1_23[96],stage1_22[127],stage1_21[167]}
   );
   gpc606_5 gpc850 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[82],stage1_23[97],stage1_22[128],stage1_21[168]}
   );
   gpc606_5 gpc851 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[83],stage1_23[98],stage1_22[129],stage1_21[169]}
   );
   gpc606_5 gpc852 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[84],stage1_23[99],stage1_22[130],stage1_21[170]}
   );
   gpc606_5 gpc853 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[85],stage1_23[100],stage1_22[131],stage1_21[171]}
   );
   gpc606_5 gpc854 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[86],stage1_23[101],stage1_22[132],stage1_21[172]}
   );
   gpc606_5 gpc855 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[87],stage1_23[102],stage1_22[133],stage1_21[173]}
   );
   gpc606_5 gpc856 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[88],stage1_23[103],stage1_22[134],stage1_21[174]}
   );
   gpc606_5 gpc857 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[89],stage1_23[104],stage1_22[135],stage1_21[175]}
   );
   gpc606_5 gpc858 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[90],stage1_23[105],stage1_22[136],stage1_21[176]}
   );
   gpc606_5 gpc859 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[91],stage1_23[106],stage1_22[137],stage1_21[177]}
   );
   gpc606_5 gpc860 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[92],stage1_23[107],stage1_22[138],stage1_21[178]}
   );
   gpc606_5 gpc861 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[93],stage1_23[108],stage1_22[139],stage1_21[179]}
   );
   gpc606_5 gpc862 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[94],stage1_23[109],stage1_22[140],stage1_21[180]}
   );
   gpc606_5 gpc863 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[95],stage1_23[110],stage1_22[141],stage1_21[181]}
   );
   gpc606_5 gpc864 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[96],stage1_23[111],stage1_22[142],stage1_21[182]}
   );
   gpc606_5 gpc865 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[97],stage1_23[112],stage1_22[143],stage1_21[183]}
   );
   gpc606_5 gpc866 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[98],stage1_23[113],stage1_22[144],stage1_21[184]}
   );
   gpc606_5 gpc867 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[99],stage1_23[114],stage1_22[145],stage1_21[185]}
   );
   gpc606_5 gpc868 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[100],stage1_23[115],stage1_22[146],stage1_21[186]}
   );
   gpc606_5 gpc869 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[101],stage1_23[116],stage1_22[147],stage1_21[187]}
   );
   gpc606_5 gpc870 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[102],stage1_23[117],stage1_22[148],stage1_21[188]}
   );
   gpc606_5 gpc871 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[103],stage1_23[118],stage1_22[149],stage1_21[189]}
   );
   gpc606_5 gpc872 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[104],stage1_23[119],stage1_22[150],stage1_21[190]}
   );
   gpc606_5 gpc873 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[105],stage1_23[120],stage1_22[151],stage1_21[191]}
   );
   gpc606_5 gpc874 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[106],stage1_23[121],stage1_22[152],stage1_21[192]}
   );
   gpc606_5 gpc875 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[107],stage1_23[122],stage1_22[153],stage1_21[193]}
   );
   gpc606_5 gpc876 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[108],stage1_23[123],stage1_22[154],stage1_21[194]}
   );
   gpc606_5 gpc877 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[109],stage1_23[124],stage1_22[155],stage1_21[195]}
   );
   gpc606_5 gpc878 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[110],stage1_23[125],stage1_22[156],stage1_21[196]}
   );
   gpc606_5 gpc879 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[111],stage1_23[126],stage1_22[157],stage1_21[197]}
   );
   gpc606_5 gpc880 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[112],stage1_23[127],stage1_22[158],stage1_21[198]}
   );
   gpc615_5 gpc881 (
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286]},
      {stage0_23[396]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[66],stage1_24[113],stage1_23[128],stage1_22[159]}
   );
   gpc615_5 gpc882 (
      {stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291]},
      {stage0_23[397]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[67],stage1_24[114],stage1_23[129],stage1_22[160]}
   );
   gpc615_5 gpc883 (
      {stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage0_23[398]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[68],stage1_24[115],stage1_23[130],stage1_22[161]}
   );
   gpc615_5 gpc884 (
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301]},
      {stage0_23[399]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[69],stage1_24[116],stage1_23[131],stage1_22[162]}
   );
   gpc615_5 gpc885 (
      {stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306]},
      {stage0_23[400]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[70],stage1_24[117],stage1_23[132],stage1_22[163]}
   );
   gpc615_5 gpc886 (
      {stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage0_23[401]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[71],stage1_24[118],stage1_23[133],stage1_22[164]}
   );
   gpc615_5 gpc887 (
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316]},
      {stage0_23[402]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[72],stage1_24[119],stage1_23[134],stage1_22[165]}
   );
   gpc615_5 gpc888 (
      {stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321]},
      {stage0_23[403]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[73],stage1_24[120],stage1_23[135],stage1_22[166]}
   );
   gpc615_5 gpc889 (
      {stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage0_23[404]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[74],stage1_24[121],stage1_23[136],stage1_22[167]}
   );
   gpc615_5 gpc890 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331]},
      {stage0_23[405]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[75],stage1_24[122],stage1_23[137],stage1_22[168]}
   );
   gpc615_5 gpc891 (
      {stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336]},
      {stage0_23[406]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[76],stage1_24[123],stage1_23[138],stage1_22[169]}
   );
   gpc615_5 gpc892 (
      {stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage0_23[407]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[77],stage1_24[124],stage1_23[139],stage1_22[170]}
   );
   gpc615_5 gpc893 (
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346]},
      {stage0_23[408]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[78],stage1_24[125],stage1_23[140],stage1_22[171]}
   );
   gpc615_5 gpc894 (
      {stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351]},
      {stage0_23[409]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[79],stage1_24[126],stage1_23[141],stage1_22[172]}
   );
   gpc615_5 gpc895 (
      {stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_23[410]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[80],stage1_24[127],stage1_23[142],stage1_22[173]}
   );
   gpc615_5 gpc896 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361]},
      {stage0_23[411]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[81],stage1_24[128],stage1_23[143],stage1_22[174]}
   );
   gpc615_5 gpc897 (
      {stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366]},
      {stage0_23[412]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[82],stage1_24[129],stage1_23[144],stage1_22[175]}
   );
   gpc615_5 gpc898 (
      {stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage0_23[413]},
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage1_26[17],stage1_25[83],stage1_24[130],stage1_23[145],stage1_22[176]}
   );
   gpc615_5 gpc899 (
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376]},
      {stage0_23[414]},
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage1_26[18],stage1_25[84],stage1_24[131],stage1_23[146],stage1_22[177]}
   );
   gpc615_5 gpc900 (
      {stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381]},
      {stage0_23[415]},
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage1_26[19],stage1_25[85],stage1_24[132],stage1_23[147],stage1_22[178]}
   );
   gpc615_5 gpc901 (
      {stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_23[416]},
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage1_26[20],stage1_25[86],stage1_24[133],stage1_23[148],stage1_22[179]}
   );
   gpc615_5 gpc902 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[417]},
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage1_26[21],stage1_25[87],stage1_24[134],stage1_23[149],stage1_22[180]}
   );
   gpc615_5 gpc903 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[418]},
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage1_26[22],stage1_25[88],stage1_24[135],stage1_23[150],stage1_22[181]}
   );
   gpc615_5 gpc904 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[419]},
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage1_26[23],stage1_25[89],stage1_24[136],stage1_23[151],stage1_22[182]}
   );
   gpc615_5 gpc905 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[420]},
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage1_26[24],stage1_25[90],stage1_24[137],stage1_23[152],stage1_22[183]}
   );
   gpc615_5 gpc906 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[421]},
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage1_26[25],stage1_25[91],stage1_24[138],stage1_23[153],stage1_22[184]}
   );
   gpc615_5 gpc907 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[422]},
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage1_26[26],stage1_25[92],stage1_24[139],stage1_23[154],stage1_22[185]}
   );
   gpc615_5 gpc908 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[423]},
      {stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167]},
      {stage1_26[27],stage1_25[93],stage1_24[140],stage1_23[155],stage1_22[186]}
   );
   gpc615_5 gpc909 (
      {stage0_23[424], stage0_23[425], stage0_23[426], stage0_23[427], stage0_23[428]},
      {stage0_24[168]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[28],stage1_25[94],stage1_24[141],stage1_23[156]}
   );
   gpc615_5 gpc910 (
      {stage0_23[429], stage0_23[430], stage0_23[431], stage0_23[432], stage0_23[433]},
      {stage0_24[169]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[29],stage1_25[95],stage1_24[142],stage1_23[157]}
   );
   gpc615_5 gpc911 (
      {stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437], stage0_23[438]},
      {stage0_24[170]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[30],stage1_25[96],stage1_24[143],stage1_23[158]}
   );
   gpc615_5 gpc912 (
      {stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage0_24[171]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[31],stage1_25[97],stage1_24[144],stage1_23[159]}
   );
   gpc615_5 gpc913 (
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448]},
      {stage0_24[172]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[32],stage1_25[98],stage1_24[145],stage1_23[160]}
   );
   gpc615_5 gpc914 (
      {stage0_23[449], stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453]},
      {stage0_24[173]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[33],stage1_25[99],stage1_24[146],stage1_23[161]}
   );
   gpc615_5 gpc915 (
      {stage0_23[454], stage0_23[455], stage0_23[456], stage0_23[457], stage0_23[458]},
      {stage0_24[174]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[34],stage1_25[100],stage1_24[147],stage1_23[162]}
   );
   gpc615_5 gpc916 (
      {stage0_23[459], stage0_23[460], stage0_23[461], stage0_23[462], stage0_23[463]},
      {stage0_24[175]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[35],stage1_25[101],stage1_24[148],stage1_23[163]}
   );
   gpc615_5 gpc917 (
      {stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467], stage0_23[468]},
      {stage0_24[176]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[36],stage1_25[102],stage1_24[149],stage1_23[164]}
   );
   gpc615_5 gpc918 (
      {stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage0_24[177]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[37],stage1_25[103],stage1_24[150],stage1_23[165]}
   );
   gpc606_5 gpc919 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[38],stage1_25[104],stage1_24[151]}
   );
   gpc606_5 gpc920 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[39],stage1_25[105],stage1_24[152]}
   );
   gpc606_5 gpc921 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[40],stage1_25[106],stage1_24[153]}
   );
   gpc615_5 gpc922 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200]},
      {stage0_25[60]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[41],stage1_25[107],stage1_24[154]}
   );
   gpc615_5 gpc923 (
      {stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205]},
      {stage0_25[61]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[42],stage1_25[108],stage1_24[155]}
   );
   gpc615_5 gpc924 (
      {stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_25[62]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[43],stage1_25[109],stage1_24[156]}
   );
   gpc615_5 gpc925 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215]},
      {stage0_25[63]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[44],stage1_25[110],stage1_24[157]}
   );
   gpc615_5 gpc926 (
      {stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_25[64]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[45],stage1_25[111],stage1_24[158]}
   );
   gpc615_5 gpc927 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_25[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[46],stage1_25[112],stage1_24[159]}
   );
   gpc615_5 gpc928 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230]},
      {stage0_25[66]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[47],stage1_25[113],stage1_24[160]}
   );
   gpc615_5 gpc929 (
      {stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235]},
      {stage0_25[67]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[48],stage1_25[114],stage1_24[161]}
   );
   gpc615_5 gpc930 (
      {stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_25[68]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[49],stage1_25[115],stage1_24[162]}
   );
   gpc615_5 gpc931 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245]},
      {stage0_25[69]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[22],stage1_26[50],stage1_25[116],stage1_24[163]}
   );
   gpc615_5 gpc932 (
      {stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_25[70]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[23],stage1_26[51],stage1_25[117],stage1_24[164]}
   );
   gpc615_5 gpc933 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_25[71]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[24],stage1_26[52],stage1_25[118],stage1_24[165]}
   );
   gpc615_5 gpc934 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260]},
      {stage0_25[72]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[25],stage1_26[53],stage1_25[119],stage1_24[166]}
   );
   gpc615_5 gpc935 (
      {stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265]},
      {stage0_25[73]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[26],stage1_26[54],stage1_25[120],stage1_24[167]}
   );
   gpc615_5 gpc936 (
      {stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_25[74]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[27],stage1_26[55],stage1_25[121],stage1_24[168]}
   );
   gpc615_5 gpc937 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275]},
      {stage0_25[75]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[28],stage1_26[56],stage1_25[122],stage1_24[169]}
   );
   gpc615_5 gpc938 (
      {stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_25[76]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[29],stage1_26[57],stage1_25[123],stage1_24[170]}
   );
   gpc615_5 gpc939 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_25[77]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[30],stage1_26[58],stage1_25[124],stage1_24[171]}
   );
   gpc615_5 gpc940 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290]},
      {stage0_25[78]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[31],stage1_26[59],stage1_25[125],stage1_24[172]}
   );
   gpc615_5 gpc941 (
      {stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295]},
      {stage0_25[79]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[32],stage1_26[60],stage1_25[126],stage1_24[173]}
   );
   gpc615_5 gpc942 (
      {stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_25[80]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[33],stage1_26[61],stage1_25[127],stage1_24[174]}
   );
   gpc615_5 gpc943 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305]},
      {stage0_25[81]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[34],stage1_26[62],stage1_25[128],stage1_24[175]}
   );
   gpc615_5 gpc944 (
      {stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_25[82]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[35],stage1_26[63],stage1_25[129],stage1_24[176]}
   );
   gpc615_5 gpc945 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_25[83]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[36],stage1_26[64],stage1_25[130],stage1_24[177]}
   );
   gpc615_5 gpc946 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320]},
      {stage0_25[84]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[37],stage1_26[65],stage1_25[131],stage1_24[178]}
   );
   gpc615_5 gpc947 (
      {stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325]},
      {stage0_25[85]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[38],stage1_26[66],stage1_25[132],stage1_24[179]}
   );
   gpc615_5 gpc948 (
      {stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_25[86]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[39],stage1_26[67],stage1_25[133],stage1_24[180]}
   );
   gpc615_5 gpc949 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335]},
      {stage0_25[87]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[40],stage1_26[68],stage1_25[134],stage1_24[181]}
   );
   gpc615_5 gpc950 (
      {stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_25[88]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[41],stage1_26[69],stage1_25[135],stage1_24[182]}
   );
   gpc615_5 gpc951 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_25[89]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[42],stage1_26[70],stage1_25[136],stage1_24[183]}
   );
   gpc615_5 gpc952 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350]},
      {stage0_25[90]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[43],stage1_26[71],stage1_25[137],stage1_24[184]}
   );
   gpc615_5 gpc953 (
      {stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355]},
      {stage0_25[91]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[44],stage1_26[72],stage1_25[138],stage1_24[185]}
   );
   gpc615_5 gpc954 (
      {stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_25[92]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[45],stage1_26[73],stage1_25[139],stage1_24[186]}
   );
   gpc615_5 gpc955 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365]},
      {stage0_25[93]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[46],stage1_26[74],stage1_25[140],stage1_24[187]}
   );
   gpc615_5 gpc956 (
      {stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_25[94]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[47],stage1_26[75],stage1_25[141],stage1_24[188]}
   );
   gpc615_5 gpc957 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375]},
      {stage0_25[95]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[48],stage1_26[76],stage1_25[142],stage1_24[189]}
   );
   gpc615_5 gpc958 (
      {stage0_24[376], stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380]},
      {stage0_25[96]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[49],stage1_26[77],stage1_25[143],stage1_24[190]}
   );
   gpc615_5 gpc959 (
      {stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385]},
      {stage0_25[97]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[50],stage1_26[78],stage1_25[144],stage1_24[191]}
   );
   gpc615_5 gpc960 (
      {stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_25[98]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[51],stage1_26[79],stage1_25[145],stage1_24[192]}
   );
   gpc615_5 gpc961 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395]},
      {stage0_25[99]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[52],stage1_26[80],stage1_25[146],stage1_24[193]}
   );
   gpc615_5 gpc962 (
      {stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_25[100]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[53],stage1_26[81],stage1_25[147],stage1_24[194]}
   );
   gpc615_5 gpc963 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405]},
      {stage0_25[101]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[54],stage1_26[82],stage1_25[148],stage1_24[195]}
   );
   gpc615_5 gpc964 (
      {stage0_24[406], stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410]},
      {stage0_25[102]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[55],stage1_26[83],stage1_25[149],stage1_24[196]}
   );
   gpc615_5 gpc965 (
      {stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415]},
      {stage0_25[103]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[56],stage1_26[84],stage1_25[150],stage1_24[197]}
   );
   gpc615_5 gpc966 (
      {stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_25[104]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[57],stage1_26[85],stage1_25[151],stage1_24[198]}
   );
   gpc615_5 gpc967 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425]},
      {stage0_25[105]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[58],stage1_26[86],stage1_25[152],stage1_24[199]}
   );
   gpc615_5 gpc968 (
      {stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_25[106]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[59],stage1_26[87],stage1_25[153],stage1_24[200]}
   );
   gpc615_5 gpc969 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435]},
      {stage0_25[107]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[60],stage1_26[88],stage1_25[154],stage1_24[201]}
   );
   gpc615_5 gpc970 (
      {stage0_24[436], stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440]},
      {stage0_25[108]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[61],stage1_26[89],stage1_25[155],stage1_24[202]}
   );
   gpc615_5 gpc971 (
      {stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445]},
      {stage0_25[109]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[62],stage1_26[90],stage1_25[156],stage1_24[203]}
   );
   gpc615_5 gpc972 (
      {stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_25[110]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[63],stage1_26[91],stage1_25[157],stage1_24[204]}
   );
   gpc615_5 gpc973 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455]},
      {stage0_25[111]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[64],stage1_26[92],stage1_25[158],stage1_24[205]}
   );
   gpc615_5 gpc974 (
      {stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_25[112]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[65],stage1_26[93],stage1_25[159],stage1_24[206]}
   );
   gpc615_5 gpc975 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465]},
      {stage0_25[113]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[66],stage1_26[94],stage1_25[160],stage1_24[207]}
   );
   gpc615_5 gpc976 (
      {stage0_24[466], stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470]},
      {stage0_25[114]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[67],stage1_26[95],stage1_25[161],stage1_24[208]}
   );
   gpc615_5 gpc977 (
      {stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475]},
      {stage0_25[115]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[68],stage1_26[96],stage1_25[162],stage1_24[209]}
   );
   gpc615_5 gpc978 (
      {stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_25[116]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[69],stage1_26[97],stage1_25[163],stage1_24[210]}
   );
   gpc615_5 gpc979 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485]},
      {stage0_25[117]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[70],stage1_26[98],stage1_25[164],stage1_24[211]}
   );
   gpc606_5 gpc980 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[61],stage1_27[71],stage1_26[99],stage1_25[165]}
   );
   gpc606_5 gpc981 (
      {stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[62],stage1_27[72],stage1_26[100],stage1_25[166]}
   );
   gpc606_5 gpc982 (
      {stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[63],stage1_27[73],stage1_26[101],stage1_25[167]}
   );
   gpc606_5 gpc983 (
      {stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[64],stage1_27[74],stage1_26[102],stage1_25[168]}
   );
   gpc606_5 gpc984 (
      {stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[65],stage1_27[75],stage1_26[103],stage1_25[169]}
   );
   gpc606_5 gpc985 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[66],stage1_27[76],stage1_26[104],stage1_25[170]}
   );
   gpc606_5 gpc986 (
      {stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[67],stage1_27[77],stage1_26[105],stage1_25[171]}
   );
   gpc606_5 gpc987 (
      {stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[68],stage1_27[78],stage1_26[106],stage1_25[172]}
   );
   gpc606_5 gpc988 (
      {stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[69],stage1_27[79],stage1_26[107],stage1_25[173]}
   );
   gpc606_5 gpc989 (
      {stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[70],stage1_27[80],stage1_26[108],stage1_25[174]}
   );
   gpc606_5 gpc990 (
      {stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[71],stage1_27[81],stage1_26[109],stage1_25[175]}
   );
   gpc606_5 gpc991 (
      {stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[72],stage1_27[82],stage1_26[110],stage1_25[176]}
   );
   gpc606_5 gpc992 (
      {stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[73],stage1_27[83],stage1_26[111],stage1_25[177]}
   );
   gpc606_5 gpc993 (
      {stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[74],stage1_27[84],stage1_26[112],stage1_25[178]}
   );
   gpc606_5 gpc994 (
      {stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[75],stage1_27[85],stage1_26[113],stage1_25[179]}
   );
   gpc606_5 gpc995 (
      {stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[76],stage1_27[86],stage1_26[114],stage1_25[180]}
   );
   gpc606_5 gpc996 (
      {stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[77],stage1_27[87],stage1_26[115],stage1_25[181]}
   );
   gpc606_5 gpc997 (
      {stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[78],stage1_27[88],stage1_26[116],stage1_25[182]}
   );
   gpc615_5 gpc998 (
      {stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229], stage0_25[230]},
      {stage0_26[366]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[79],stage1_27[89],stage1_26[117],stage1_25[183]}
   );
   gpc615_5 gpc999 (
      {stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_26[367]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[80],stage1_27[90],stage1_26[118],stage1_25[184]}
   );
   gpc615_5 gpc1000 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240]},
      {stage0_26[368]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[81],stage1_27[91],stage1_26[119],stage1_25[185]}
   );
   gpc615_5 gpc1001 (
      {stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_26[369]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[82],stage1_27[92],stage1_26[120],stage1_25[186]}
   );
   gpc615_5 gpc1002 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[370]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[83],stage1_27[93],stage1_26[121],stage1_25[187]}
   );
   gpc615_5 gpc1003 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[371]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[84],stage1_27[94],stage1_26[122],stage1_25[188]}
   );
   gpc615_5 gpc1004 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[372]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[85],stage1_27[95],stage1_26[123],stage1_25[189]}
   );
   gpc615_5 gpc1005 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[373]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[86],stage1_27[96],stage1_26[124],stage1_25[190]}
   );
   gpc615_5 gpc1006 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[374]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[87],stage1_27[97],stage1_26[125],stage1_25[191]}
   );
   gpc615_5 gpc1007 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[375]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[88],stage1_27[98],stage1_26[126],stage1_25[192]}
   );
   gpc615_5 gpc1008 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[376]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[89],stage1_27[99],stage1_26[127],stage1_25[193]}
   );
   gpc615_5 gpc1009 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[377]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[90],stage1_27[100],stage1_26[128],stage1_25[194]}
   );
   gpc615_5 gpc1010 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[378]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[91],stage1_27[101],stage1_26[129],stage1_25[195]}
   );
   gpc615_5 gpc1011 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[379]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[92],stage1_27[102],stage1_26[130],stage1_25[196]}
   );
   gpc615_5 gpc1012 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[380]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[93],stage1_27[103],stage1_26[131],stage1_25[197]}
   );
   gpc615_5 gpc1013 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[381]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[94],stage1_27[104],stage1_26[132],stage1_25[198]}
   );
   gpc615_5 gpc1014 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[382]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[95],stage1_27[105],stage1_26[133],stage1_25[199]}
   );
   gpc615_5 gpc1015 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[383]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[96],stage1_27[106],stage1_26[134],stage1_25[200]}
   );
   gpc615_5 gpc1016 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[384]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[97],stage1_27[107],stage1_26[135],stage1_25[201]}
   );
   gpc615_5 gpc1017 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[385]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[98],stage1_27[108],stage1_26[136],stage1_25[202]}
   );
   gpc615_5 gpc1018 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[386]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[99],stage1_27[109],stage1_26[137],stage1_25[203]}
   );
   gpc615_5 gpc1019 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[387]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[100],stage1_27[110],stage1_26[138],stage1_25[204]}
   );
   gpc615_5 gpc1020 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[388]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[101],stage1_27[111],stage1_26[139],stage1_25[205]}
   );
   gpc615_5 gpc1021 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[389]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[102],stage1_27[112],stage1_26[140],stage1_25[206]}
   );
   gpc615_5 gpc1022 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[390]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[103],stage1_27[113],stage1_26[141],stage1_25[207]}
   );
   gpc615_5 gpc1023 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[391]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[104],stage1_27[114],stage1_26[142],stage1_25[208]}
   );
   gpc615_5 gpc1024 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[392]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[105],stage1_27[115],stage1_26[143],stage1_25[209]}
   );
   gpc615_5 gpc1025 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[393]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[106],stage1_27[116],stage1_26[144],stage1_25[210]}
   );
   gpc615_5 gpc1026 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[394]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[107],stage1_27[117],stage1_26[145],stage1_25[211]}
   );
   gpc615_5 gpc1027 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[395]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[108],stage1_27[118],stage1_26[146],stage1_25[212]}
   );
   gpc615_5 gpc1028 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[396]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[109],stage1_27[119],stage1_26[147],stage1_25[213]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[397]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[110],stage1_27[120],stage1_26[148],stage1_25[214]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[398]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[111],stage1_27[121],stage1_26[149],stage1_25[215]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[399]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[112],stage1_27[122],stage1_26[150],stage1_25[216]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[400]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[113],stage1_27[123],stage1_26[151],stage1_25[217]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[401]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[114],stage1_27[124],stage1_26[152],stage1_25[218]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[402]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[115],stage1_27[125],stage1_26[153],stage1_25[219]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[403]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[116],stage1_27[126],stage1_26[154],stage1_25[220]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[404]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[117],stage1_27[127],stage1_26[155],stage1_25[221]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[405]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[118],stage1_27[128],stage1_26[156],stage1_25[222]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[406]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[119],stage1_27[129],stage1_26[157],stage1_25[223]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[407]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[120],stage1_27[130],stage1_26[158],stage1_25[224]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[408]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[121],stage1_27[131],stage1_26[159],stage1_25[225]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[409]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[122],stage1_27[132],stage1_26[160],stage1_25[226]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[410]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[123],stage1_27[133],stage1_26[161],stage1_25[227]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[411]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[124],stage1_27[134],stage1_26[162],stage1_25[228]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[412]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[125],stage1_27[135],stage1_26[163],stage1_25[229]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[413]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[126],stage1_27[136],stage1_26[164],stage1_25[230]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[414]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[127],stage1_27[137],stage1_26[165],stage1_25[231]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[415]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[128],stage1_27[138],stage1_26[166],stage1_25[232]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[416]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[129],stage1_27[139],stage1_26[167],stage1_25[233]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[417]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[130],stage1_27[140],stage1_26[168],stage1_25[234]}
   );
   gpc606_5 gpc1050 (
      {stage0_26[418], stage0_26[419], stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[70],stage1_28[131],stage1_27[141],stage1_26[169]}
   );
   gpc606_5 gpc1051 (
      {stage0_26[424], stage0_26[425], stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[71],stage1_28[132],stage1_27[142],stage1_26[170]}
   );
   gpc615_5 gpc1052 (
      {stage0_26[430], stage0_26[431], stage0_26[432], stage0_26[433], stage0_26[434]},
      {stage0_27[420]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[72],stage1_28[133],stage1_27[143],stage1_26[171]}
   );
   gpc615_5 gpc1053 (
      {stage0_26[435], stage0_26[436], stage0_26[437], stage0_26[438], stage0_26[439]},
      {stage0_27[421]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[73],stage1_28[134],stage1_27[144],stage1_26[172]}
   );
   gpc615_5 gpc1054 (
      {stage0_26[440], stage0_26[441], stage0_26[442], stage0_26[443], stage0_26[444]},
      {stage0_27[422]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[74],stage1_28[135],stage1_27[145],stage1_26[173]}
   );
   gpc606_5 gpc1055 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427], stage0_27[428]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[75],stage1_28[136],stage1_27[146]}
   );
   gpc606_5 gpc1056 (
      {stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432], stage0_27[433], stage0_27[434]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[76],stage1_28[137],stage1_27[147]}
   );
   gpc606_5 gpc1057 (
      {stage0_27[435], stage0_27[436], stage0_27[437], stage0_27[438], stage0_27[439], stage0_27[440]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[77],stage1_28[138],stage1_27[148]}
   );
   gpc606_5 gpc1058 (
      {stage0_27[441], stage0_27[442], stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[78],stage1_28[139],stage1_27[149]}
   );
   gpc606_5 gpc1059 (
      {stage0_27[447], stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[79],stage1_28[140],stage1_27[150]}
   );
   gpc606_5 gpc1060 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457], stage0_27[458]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[80],stage1_28[141],stage1_27[151]}
   );
   gpc606_5 gpc1061 (
      {stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462], stage0_27[463], stage0_27[464]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[81],stage1_28[142],stage1_27[152]}
   );
   gpc606_5 gpc1062 (
      {stage0_27[465], stage0_27[466], stage0_27[467], stage0_27[468], stage0_27[469], stage0_27[470]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[82],stage1_28[143],stage1_27[153]}
   );
   gpc606_5 gpc1063 (
      {stage0_27[471], stage0_27[472], stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[83],stage1_28[144],stage1_27[154]}
   );
   gpc606_5 gpc1064 (
      {stage0_27[477], stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[84],stage1_28[145],stage1_27[155]}
   );
   gpc606_5 gpc1065 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[10],stage1_30[15],stage1_29[85],stage1_28[146]}
   );
   gpc606_5 gpc1066 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[11],stage1_30[16],stage1_29[86],stage1_28[147]}
   );
   gpc606_5 gpc1067 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[12],stage1_30[17],stage1_29[87],stage1_28[148]}
   );
   gpc606_5 gpc1068 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[13],stage1_30[18],stage1_29[88],stage1_28[149]}
   );
   gpc606_5 gpc1069 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[14],stage1_30[19],stage1_29[89],stage1_28[150]}
   );
   gpc606_5 gpc1070 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[15],stage1_30[20],stage1_29[90],stage1_28[151]}
   );
   gpc606_5 gpc1071 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[16],stage1_30[21],stage1_29[91],stage1_28[152]}
   );
   gpc606_5 gpc1072 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[17],stage1_30[22],stage1_29[92],stage1_28[153]}
   );
   gpc606_5 gpc1073 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[18],stage1_30[23],stage1_29[93],stage1_28[154]}
   );
   gpc606_5 gpc1074 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[19],stage1_30[24],stage1_29[94],stage1_28[155]}
   );
   gpc606_5 gpc1075 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[20],stage1_30[25],stage1_29[95],stage1_28[156]}
   );
   gpc606_5 gpc1076 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[21],stage1_30[26],stage1_29[96],stage1_28[157]}
   );
   gpc606_5 gpc1077 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[22],stage1_30[27],stage1_29[97],stage1_28[158]}
   );
   gpc606_5 gpc1078 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[23],stage1_30[28],stage1_29[98],stage1_28[159]}
   );
   gpc606_5 gpc1079 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[24],stage1_30[29],stage1_29[99],stage1_28[160]}
   );
   gpc606_5 gpc1080 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[25],stage1_30[30],stage1_29[100],stage1_28[161]}
   );
   gpc606_5 gpc1081 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[26],stage1_30[31],stage1_29[101],stage1_28[162]}
   );
   gpc606_5 gpc1082 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[27],stage1_30[32],stage1_29[102],stage1_28[163]}
   );
   gpc606_5 gpc1083 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[28],stage1_30[33],stage1_29[103],stage1_28[164]}
   );
   gpc606_5 gpc1084 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[29],stage1_30[34],stage1_29[104],stage1_28[165]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[30],stage1_30[35],stage1_29[105],stage1_28[166]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[31],stage1_30[36],stage1_29[106],stage1_28[167]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[32],stage1_30[37],stage1_29[107],stage1_28[168]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[33],stage1_30[38],stage1_29[108],stage1_28[169]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[34],stage1_30[39],stage1_29[109],stage1_28[170]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[35],stage1_30[40],stage1_29[110],stage1_28[171]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[36],stage1_30[41],stage1_29[111],stage1_28[172]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[37],stage1_30[42],stage1_29[112],stage1_28[173]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[38],stage1_30[43],stage1_29[113],stage1_28[174]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[39],stage1_30[44],stage1_29[114],stage1_28[175]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[40],stage1_30[45],stage1_29[115],stage1_28[176]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[41],stage1_30[46],stage1_29[116],stage1_28[177]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[42],stage1_30[47],stage1_29[117],stage1_28[178]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[43],stage1_30[48],stage1_29[118],stage1_28[179]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[44],stage1_30[49],stage1_29[119],stage1_28[180]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[240], stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[45],stage1_30[50],stage1_29[120],stage1_28[181]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[246], stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[46],stage1_30[51],stage1_29[121],stage1_28[182]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[252], stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[47],stage1_30[52],stage1_29[122],stage1_28[183]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[258], stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[48],stage1_30[53],stage1_29[123],stage1_28[184]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[264], stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[49],stage1_30[54],stage1_29[124],stage1_28[185]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[270], stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[50],stage1_30[55],stage1_29[125],stage1_28[186]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[276], stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[51],stage1_30[56],stage1_29[126],stage1_28[187]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[282], stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[52],stage1_30[57],stage1_29[127],stage1_28[188]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[288], stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[53],stage1_30[58],stage1_29[128],stage1_28[189]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[294], stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[54],stage1_30[59],stage1_29[129],stage1_28[190]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[300], stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[55],stage1_30[60],stage1_29[130],stage1_28[191]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[56],stage1_30[61],stage1_29[131],stage1_28[192]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[57],stage1_30[62],stage1_29[132],stage1_28[193]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[318], stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[58],stage1_30[63],stage1_29[133],stage1_28[194]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[324], stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[59],stage1_30[64],stage1_29[134],stage1_28[195]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[330], stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[60],stage1_30[65],stage1_29[135],stage1_28[196]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[61],stage1_30[66],stage1_29[136],stage1_28[197]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[62],stage1_30[67],stage1_29[137],stage1_28[198]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[348], stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[63],stage1_30[68],stage1_29[138],stage1_28[199]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[354], stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[64],stage1_30[69],stage1_29[139],stage1_28[200]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[360], stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[65],stage1_30[70],stage1_29[140],stage1_28[201]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[66],stage1_30[71],stage1_29[141],stage1_28[202]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[67],stage1_30[72],stage1_29[142],stage1_28[203]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[378], stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[68],stage1_30[73],stage1_29[143],stage1_28[204]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[384], stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[69],stage1_30[74],stage1_29[144],stage1_28[205]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[390], stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[70],stage1_30[75],stage1_29[145],stage1_28[206]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[71],stage1_30[76],stage1_29[146],stage1_28[207]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[72],stage1_30[77],stage1_29[147],stage1_28[208]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[408], stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[73],stage1_30[78],stage1_29[148],stage1_28[209]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[414], stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[74],stage1_30[79],stage1_29[149],stage1_28[210]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[420], stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[75],stage1_30[80],stage1_29[150],stage1_28[211]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[76],stage1_30[81],stage1_29[151],stage1_28[212]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[77],stage1_30[82],stage1_29[152],stage1_28[213]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[438], stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[78],stage1_30[83],stage1_29[153],stage1_28[214]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[444], stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[79],stage1_30[84],stage1_29[154],stage1_28[215]}
   );
   gpc606_5 gpc1135 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[70],stage1_31[80],stage1_30[85],stage1_29[155]}
   );
   gpc606_5 gpc1136 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[71],stage1_31[81],stage1_30[86],stage1_29[156]}
   );
   gpc606_5 gpc1137 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[72],stage1_31[82],stage1_30[87],stage1_29[157]}
   );
   gpc606_5 gpc1138 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[73],stage1_31[83],stage1_30[88],stage1_29[158]}
   );
   gpc606_5 gpc1139 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[74],stage1_31[84],stage1_30[89],stage1_29[159]}
   );
   gpc606_5 gpc1140 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[75],stage1_31[85],stage1_30[90],stage1_29[160]}
   );
   gpc606_5 gpc1141 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[76],stage1_31[86],stage1_30[91],stage1_29[161]}
   );
   gpc606_5 gpc1142 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[77],stage1_31[87],stage1_30[92],stage1_29[162]}
   );
   gpc606_5 gpc1143 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[78],stage1_31[88],stage1_30[93],stage1_29[163]}
   );
   gpc606_5 gpc1144 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[79],stage1_31[89],stage1_30[94],stage1_29[164]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[80],stage1_31[90],stage1_30[95],stage1_29[165]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[81],stage1_31[91],stage1_30[96],stage1_29[166]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[82],stage1_31[92],stage1_30[97],stage1_29[167]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[83],stage1_31[93],stage1_30[98],stage1_29[168]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[84],stage1_31[94],stage1_30[99],stage1_29[169]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[85],stage1_31[95],stage1_30[100],stage1_29[170]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[86],stage1_31[96],stage1_30[101],stage1_29[171]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[87],stage1_31[97],stage1_30[102],stage1_29[172]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[88],stage1_31[98],stage1_30[103],stage1_29[173]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[89],stage1_31[99],stage1_30[104],stage1_29[174]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[90],stage1_31[100],stage1_30[105],stage1_29[175]}
   );
   gpc615_5 gpc1156 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_30[420]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[91],stage1_31[101],stage1_30[106],stage1_29[176]}
   );
   gpc615_5 gpc1157 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195]},
      {stage0_30[421]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[92],stage1_31[102],stage1_30[107],stage1_29[177]}
   );
   gpc615_5 gpc1158 (
      {stage0_29[196], stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200]},
      {stage0_30[422]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[93],stage1_31[103],stage1_30[108],stage1_29[178]}
   );
   gpc615_5 gpc1159 (
      {stage0_29[201], stage0_29[202], stage0_29[203], stage0_29[204], stage0_29[205]},
      {stage0_30[423]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[94],stage1_31[104],stage1_30[109],stage1_29[179]}
   );
   gpc615_5 gpc1160 (
      {stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209], stage0_29[210]},
      {stage0_30[424]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[95],stage1_31[105],stage1_30[110],stage1_29[180]}
   );
   gpc615_5 gpc1161 (
      {stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_30[425]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[96],stage1_31[106],stage1_30[111],stage1_29[181]}
   );
   gpc615_5 gpc1162 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_30[426]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[97],stage1_31[107],stage1_30[112],stage1_29[182]}
   );
   gpc615_5 gpc1163 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225]},
      {stage0_30[427]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[98],stage1_31[108],stage1_30[113],stage1_29[183]}
   );
   gpc615_5 gpc1164 (
      {stage0_29[226], stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230]},
      {stage0_30[428]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[99],stage1_31[109],stage1_30[114],stage1_29[184]}
   );
   gpc615_5 gpc1165 (
      {stage0_29[231], stage0_29[232], stage0_29[233], stage0_29[234], stage0_29[235]},
      {stage0_30[429]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[100],stage1_31[110],stage1_30[115],stage1_29[185]}
   );
   gpc615_5 gpc1166 (
      {stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239], stage0_29[240]},
      {stage0_30[430]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[101],stage1_31[111],stage1_30[116],stage1_29[186]}
   );
   gpc615_5 gpc1167 (
      {stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_30[431]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[102],stage1_31[112],stage1_30[117],stage1_29[187]}
   );
   gpc615_5 gpc1168 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_30[432]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[103],stage1_31[113],stage1_30[118],stage1_29[188]}
   );
   gpc615_5 gpc1169 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255]},
      {stage0_30[433]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[104],stage1_31[114],stage1_30[119],stage1_29[189]}
   );
   gpc615_5 gpc1170 (
      {stage0_29[256], stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260]},
      {stage0_30[434]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[105],stage1_31[115],stage1_30[120],stage1_29[190]}
   );
   gpc615_5 gpc1171 (
      {stage0_29[261], stage0_29[262], stage0_29[263], stage0_29[264], stage0_29[265]},
      {stage0_30[435]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[106],stage1_31[116],stage1_30[121],stage1_29[191]}
   );
   gpc615_5 gpc1172 (
      {stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269], stage0_29[270]},
      {stage0_30[436]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[107],stage1_31[117],stage1_30[122],stage1_29[192]}
   );
   gpc615_5 gpc1173 (
      {stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_30[437]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[108],stage1_31[118],stage1_30[123],stage1_29[193]}
   );
   gpc615_5 gpc1174 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_30[438]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[109],stage1_31[119],stage1_30[124],stage1_29[194]}
   );
   gpc615_5 gpc1175 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285]},
      {stage0_30[439]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[110],stage1_31[120],stage1_30[125],stage1_29[195]}
   );
   gpc615_5 gpc1176 (
      {stage0_29[286], stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290]},
      {stage0_30[440]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[111],stage1_31[121],stage1_30[126],stage1_29[196]}
   );
   gpc615_5 gpc1177 (
      {stage0_29[291], stage0_29[292], stage0_29[293], stage0_29[294], stage0_29[295]},
      {stage0_30[441]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[112],stage1_31[122],stage1_30[127],stage1_29[197]}
   );
   gpc615_5 gpc1178 (
      {stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299], stage0_29[300]},
      {stage0_30[442]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[113],stage1_31[123],stage1_30[128],stage1_29[198]}
   );
   gpc615_5 gpc1179 (
      {stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_30[443]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[114],stage1_31[124],stage1_30[129],stage1_29[199]}
   );
   gpc615_5 gpc1180 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_30[444]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[115],stage1_31[125],stage1_30[130],stage1_29[200]}
   );
   gpc615_5 gpc1181 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315]},
      {stage0_30[445]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[116],stage1_31[126],stage1_30[131],stage1_29[201]}
   );
   gpc615_5 gpc1182 (
      {stage0_29[316], stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320]},
      {stage0_30[446]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[117],stage1_31[127],stage1_30[132],stage1_29[202]}
   );
   gpc615_5 gpc1183 (
      {stage0_29[321], stage0_29[322], stage0_29[323], stage0_29[324], stage0_29[325]},
      {stage0_30[447]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[118],stage1_31[128],stage1_30[133],stage1_29[203]}
   );
   gpc615_5 gpc1184 (
      {stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329], stage0_29[330]},
      {stage0_30[448]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[119],stage1_31[129],stage1_30[134],stage1_29[204]}
   );
   gpc615_5 gpc1185 (
      {stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_30[449]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[120],stage1_31[130],stage1_30[135],stage1_29[205]}
   );
   gpc615_5 gpc1186 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_30[450]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[121],stage1_31[131],stage1_30[136],stage1_29[206]}
   );
   gpc615_5 gpc1187 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345]},
      {stage0_30[451]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[122],stage1_31[132],stage1_30[137],stage1_29[207]}
   );
   gpc615_5 gpc1188 (
      {stage0_29[346], stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350]},
      {stage0_30[452]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[123],stage1_31[133],stage1_30[138],stage1_29[208]}
   );
   gpc615_5 gpc1189 (
      {stage0_29[351], stage0_29[352], stage0_29[353], stage0_29[354], stage0_29[355]},
      {stage0_30[453]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[124],stage1_31[134],stage1_30[139],stage1_29[209]}
   );
   gpc615_5 gpc1190 (
      {stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359], stage0_29[360]},
      {stage0_30[454]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[125],stage1_31[135],stage1_30[140],stage1_29[210]}
   );
   gpc615_5 gpc1191 (
      {stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_30[455]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[126],stage1_31[136],stage1_30[141],stage1_29[211]}
   );
   gpc615_5 gpc1192 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_30[456]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[127],stage1_31[137],stage1_30[142],stage1_29[212]}
   );
   gpc615_5 gpc1193 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375]},
      {stage0_30[457]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[128],stage1_31[138],stage1_30[143],stage1_29[213]}
   );
   gpc615_5 gpc1194 (
      {stage0_29[376], stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380]},
      {stage0_30[458]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[129],stage1_31[139],stage1_30[144],stage1_29[214]}
   );
   gpc615_5 gpc1195 (
      {stage0_29[381], stage0_29[382], stage0_29[383], stage0_29[384], stage0_29[385]},
      {stage0_30[459]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[130],stage1_31[140],stage1_30[145],stage1_29[215]}
   );
   gpc615_5 gpc1196 (
      {stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389], stage0_29[390]},
      {stage0_30[460]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[131],stage1_31[141],stage1_30[146],stage1_29[216]}
   );
   gpc615_5 gpc1197 (
      {stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_30[461]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[132],stage1_31[142],stage1_30[147],stage1_29[217]}
   );
   gpc615_5 gpc1198 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_30[462]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[133],stage1_31[143],stage1_30[148],stage1_29[218]}
   );
   gpc615_5 gpc1199 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405]},
      {stage0_30[463]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[134],stage1_31[144],stage1_30[149],stage1_29[219]}
   );
   gpc615_5 gpc1200 (
      {stage0_29[406], stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410]},
      {stage0_30[464]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[135],stage1_31[145],stage1_30[150],stage1_29[220]}
   );
   gpc615_5 gpc1201 (
      {stage0_29[411], stage0_29[412], stage0_29[413], stage0_29[414], stage0_29[415]},
      {stage0_30[465]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[136],stage1_31[146],stage1_30[151],stage1_29[221]}
   );
   gpc615_5 gpc1202 (
      {stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419], stage0_29[420]},
      {stage0_30[466]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[137],stage1_31[147],stage1_30[152],stage1_29[222]}
   );
   gpc615_5 gpc1203 (
      {stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_30[467]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[138],stage1_31[148],stage1_30[153],stage1_29[223]}
   );
   gpc615_5 gpc1204 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_30[468]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[139],stage1_31[149],stage1_30[154],stage1_29[224]}
   );
   gpc615_5 gpc1205 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435]},
      {stage0_30[469]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[140],stage1_31[150],stage1_30[155],stage1_29[225]}
   );
   gpc615_5 gpc1206 (
      {stage0_29[436], stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440]},
      {stage0_30[470]},
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430], stage0_31[431]},
      {stage1_33[71],stage1_32[141],stage1_31[151],stage1_30[156],stage1_29[226]}
   );
   gpc615_5 gpc1207 (
      {stage0_29[441], stage0_29[442], stage0_29[443], stage0_29[444], stage0_29[445]},
      {stage0_30[471]},
      {stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437]},
      {stage1_33[72],stage1_32[142],stage1_31[152],stage1_30[157],stage1_29[227]}
   );
   gpc615_5 gpc1208 (
      {stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449], stage0_29[450]},
      {stage0_30[472]},
      {stage0_31[438], stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage1_33[73],stage1_32[143],stage1_31[153],stage1_30[158],stage1_29[228]}
   );
   gpc615_5 gpc1209 (
      {stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_30[473]},
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449]},
      {stage1_33[74],stage1_32[144],stage1_31[154],stage1_30[159],stage1_29[229]}
   );
   gpc615_5 gpc1210 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_30[474]},
      {stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage1_33[75],stage1_32[145],stage1_31[155],stage1_30[160],stage1_29[230]}
   );
   gpc615_5 gpc1211 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465]},
      {stage0_30[475]},
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460], stage0_31[461]},
      {stage1_33[76],stage1_32[146],stage1_31[156],stage1_30[161],stage1_29[231]}
   );
   gpc615_5 gpc1212 (
      {stage0_29[466], stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470]},
      {stage0_30[476]},
      {stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467]},
      {stage1_33[77],stage1_32[147],stage1_31[157],stage1_30[162],stage1_29[232]}
   );
   gpc615_5 gpc1213 (
      {stage0_29[471], stage0_29[472], stage0_29[473], stage0_29[474], stage0_29[475]},
      {stage0_30[477]},
      {stage0_31[468], stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage1_33[78],stage1_32[148],stage1_31[158],stage1_30[163],stage1_29[233]}
   );
   gpc615_5 gpc1214 (
      {stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479], stage0_29[480]},
      {stage0_30[478]},
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478], stage0_31[479]},
      {stage1_33[79],stage1_32[149],stage1_31[159],stage1_30[164],stage1_29[234]}
   );
   gpc615_5 gpc1215 (
      {stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_30[479]},
      {stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483], stage0_31[484], stage0_31[485]},
      {stage1_33[80],stage1_32[150],stage1_31[160],stage1_30[165],stage1_29[235]}
   );
   gpc1_1 gpc1216 (
      {stage0_0[444]},
      {stage1_0[85]}
   );
   gpc1_1 gpc1217 (
      {stage0_0[445]},
      {stage1_0[86]}
   );
   gpc1_1 gpc1218 (
      {stage0_0[446]},
      {stage1_0[87]}
   );
   gpc1_1 gpc1219 (
      {stage0_0[447]},
      {stage1_0[88]}
   );
   gpc1_1 gpc1220 (
      {stage0_0[448]},
      {stage1_0[89]}
   );
   gpc1_1 gpc1221 (
      {stage0_0[449]},
      {stage1_0[90]}
   );
   gpc1_1 gpc1222 (
      {stage0_0[450]},
      {stage1_0[91]}
   );
   gpc1_1 gpc1223 (
      {stage0_0[451]},
      {stage1_0[92]}
   );
   gpc1_1 gpc1224 (
      {stage0_0[452]},
      {stage1_0[93]}
   );
   gpc1_1 gpc1225 (
      {stage0_0[453]},
      {stage1_0[94]}
   );
   gpc1_1 gpc1226 (
      {stage0_0[454]},
      {stage1_0[95]}
   );
   gpc1_1 gpc1227 (
      {stage0_0[455]},
      {stage1_0[96]}
   );
   gpc1_1 gpc1228 (
      {stage0_0[456]},
      {stage1_0[97]}
   );
   gpc1_1 gpc1229 (
      {stage0_0[457]},
      {stage1_0[98]}
   );
   gpc1_1 gpc1230 (
      {stage0_0[458]},
      {stage1_0[99]}
   );
   gpc1_1 gpc1231 (
      {stage0_0[459]},
      {stage1_0[100]}
   );
   gpc1_1 gpc1232 (
      {stage0_0[460]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1233 (
      {stage0_0[461]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1234 (
      {stage0_0[462]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1235 (
      {stage0_0[463]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1236 (
      {stage0_0[464]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1237 (
      {stage0_0[465]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1238 (
      {stage0_0[466]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1239 (
      {stage0_0[467]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1240 (
      {stage0_0[468]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1241 (
      {stage0_0[469]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1242 (
      {stage0_0[470]},
      {stage1_0[111]}
   );
   gpc1_1 gpc1243 (
      {stage0_0[471]},
      {stage1_0[112]}
   );
   gpc1_1 gpc1244 (
      {stage0_0[472]},
      {stage1_0[113]}
   );
   gpc1_1 gpc1245 (
      {stage0_0[473]},
      {stage1_0[114]}
   );
   gpc1_1 gpc1246 (
      {stage0_0[474]},
      {stage1_0[115]}
   );
   gpc1_1 gpc1247 (
      {stage0_0[475]},
      {stage1_0[116]}
   );
   gpc1_1 gpc1248 (
      {stage0_0[476]},
      {stage1_0[117]}
   );
   gpc1_1 gpc1249 (
      {stage0_0[477]},
      {stage1_0[118]}
   );
   gpc1_1 gpc1250 (
      {stage0_0[478]},
      {stage1_0[119]}
   );
   gpc1_1 gpc1251 (
      {stage0_0[479]},
      {stage1_0[120]}
   );
   gpc1_1 gpc1252 (
      {stage0_0[480]},
      {stage1_0[121]}
   );
   gpc1_1 gpc1253 (
      {stage0_0[481]},
      {stage1_0[122]}
   );
   gpc1_1 gpc1254 (
      {stage0_0[482]},
      {stage1_0[123]}
   );
   gpc1_1 gpc1255 (
      {stage0_0[483]},
      {stage1_0[124]}
   );
   gpc1_1 gpc1256 (
      {stage0_0[484]},
      {stage1_0[125]}
   );
   gpc1_1 gpc1257 (
      {stage0_0[485]},
      {stage1_0[126]}
   );
   gpc1_1 gpc1258 (
      {stage0_1[484]},
      {stage1_1[136]}
   );
   gpc1_1 gpc1259 (
      {stage0_1[485]},
      {stage1_1[137]}
   );
   gpc1_1 gpc1260 (
      {stage0_2[415]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1261 (
      {stage0_2[416]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1262 (
      {stage0_2[417]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1263 (
      {stage0_2[418]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1264 (
      {stage0_2[419]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1265 (
      {stage0_2[420]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1266 (
      {stage0_2[421]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1267 (
      {stage0_2[422]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1268 (
      {stage0_2[423]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1269 (
      {stage0_2[424]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1270 (
      {stage0_2[425]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1271 (
      {stage0_2[426]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1272 (
      {stage0_2[427]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1273 (
      {stage0_2[428]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1274 (
      {stage0_2[429]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1275 (
      {stage0_2[430]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1276 (
      {stage0_2[431]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1277 (
      {stage0_2[432]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1278 (
      {stage0_2[433]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1279 (
      {stage0_2[434]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1280 (
      {stage0_2[435]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1281 (
      {stage0_2[436]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1282 (
      {stage0_2[437]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1283 (
      {stage0_2[438]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1284 (
      {stage0_2[439]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1285 (
      {stage0_2[440]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1286 (
      {stage0_2[441]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1287 (
      {stage0_2[442]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1288 (
      {stage0_2[443]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1289 (
      {stage0_2[444]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1290 (
      {stage0_2[445]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1291 (
      {stage0_2[446]},
      {stage1_2[188]}
   );
   gpc1_1 gpc1292 (
      {stage0_2[447]},
      {stage1_2[189]}
   );
   gpc1_1 gpc1293 (
      {stage0_2[448]},
      {stage1_2[190]}
   );
   gpc1_1 gpc1294 (
      {stage0_2[449]},
      {stage1_2[191]}
   );
   gpc1_1 gpc1295 (
      {stage0_2[450]},
      {stage1_2[192]}
   );
   gpc1_1 gpc1296 (
      {stage0_2[451]},
      {stage1_2[193]}
   );
   gpc1_1 gpc1297 (
      {stage0_2[452]},
      {stage1_2[194]}
   );
   gpc1_1 gpc1298 (
      {stage0_2[453]},
      {stage1_2[195]}
   );
   gpc1_1 gpc1299 (
      {stage0_2[454]},
      {stage1_2[196]}
   );
   gpc1_1 gpc1300 (
      {stage0_2[455]},
      {stage1_2[197]}
   );
   gpc1_1 gpc1301 (
      {stage0_2[456]},
      {stage1_2[198]}
   );
   gpc1_1 gpc1302 (
      {stage0_2[457]},
      {stage1_2[199]}
   );
   gpc1_1 gpc1303 (
      {stage0_2[458]},
      {stage1_2[200]}
   );
   gpc1_1 gpc1304 (
      {stage0_2[459]},
      {stage1_2[201]}
   );
   gpc1_1 gpc1305 (
      {stage0_2[460]},
      {stage1_2[202]}
   );
   gpc1_1 gpc1306 (
      {stage0_2[461]},
      {stage1_2[203]}
   );
   gpc1_1 gpc1307 (
      {stage0_2[462]},
      {stage1_2[204]}
   );
   gpc1_1 gpc1308 (
      {stage0_2[463]},
      {stage1_2[205]}
   );
   gpc1_1 gpc1309 (
      {stage0_2[464]},
      {stage1_2[206]}
   );
   gpc1_1 gpc1310 (
      {stage0_2[465]},
      {stage1_2[207]}
   );
   gpc1_1 gpc1311 (
      {stage0_2[466]},
      {stage1_2[208]}
   );
   gpc1_1 gpc1312 (
      {stage0_2[467]},
      {stage1_2[209]}
   );
   gpc1_1 gpc1313 (
      {stage0_2[468]},
      {stage1_2[210]}
   );
   gpc1_1 gpc1314 (
      {stage0_2[469]},
      {stage1_2[211]}
   );
   gpc1_1 gpc1315 (
      {stage0_2[470]},
      {stage1_2[212]}
   );
   gpc1_1 gpc1316 (
      {stage0_2[471]},
      {stage1_2[213]}
   );
   gpc1_1 gpc1317 (
      {stage0_2[472]},
      {stage1_2[214]}
   );
   gpc1_1 gpc1318 (
      {stage0_2[473]},
      {stage1_2[215]}
   );
   gpc1_1 gpc1319 (
      {stage0_2[474]},
      {stage1_2[216]}
   );
   gpc1_1 gpc1320 (
      {stage0_2[475]},
      {stage1_2[217]}
   );
   gpc1_1 gpc1321 (
      {stage0_2[476]},
      {stage1_2[218]}
   );
   gpc1_1 gpc1322 (
      {stage0_2[477]},
      {stage1_2[219]}
   );
   gpc1_1 gpc1323 (
      {stage0_2[478]},
      {stage1_2[220]}
   );
   gpc1_1 gpc1324 (
      {stage0_2[479]},
      {stage1_2[221]}
   );
   gpc1_1 gpc1325 (
      {stage0_2[480]},
      {stage1_2[222]}
   );
   gpc1_1 gpc1326 (
      {stage0_2[481]},
      {stage1_2[223]}
   );
   gpc1_1 gpc1327 (
      {stage0_2[482]},
      {stage1_2[224]}
   );
   gpc1_1 gpc1328 (
      {stage0_2[483]},
      {stage1_2[225]}
   );
   gpc1_1 gpc1329 (
      {stage0_2[484]},
      {stage1_2[226]}
   );
   gpc1_1 gpc1330 (
      {stage0_2[485]},
      {stage1_2[227]}
   );
   gpc1_1 gpc1331 (
      {stage0_3[484]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1332 (
      {stage0_3[485]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1333 (
      {stage0_4[485]},
      {stage1_4[225]}
   );
   gpc1_1 gpc1334 (
      {stage0_5[474]},
      {stage1_5[206]}
   );
   gpc1_1 gpc1335 (
      {stage0_5[475]},
      {stage1_5[207]}
   );
   gpc1_1 gpc1336 (
      {stage0_5[476]},
      {stage1_5[208]}
   );
   gpc1_1 gpc1337 (
      {stage0_5[477]},
      {stage1_5[209]}
   );
   gpc1_1 gpc1338 (
      {stage0_5[478]},
      {stage1_5[210]}
   );
   gpc1_1 gpc1339 (
      {stage0_5[479]},
      {stage1_5[211]}
   );
   gpc1_1 gpc1340 (
      {stage0_5[480]},
      {stage1_5[212]}
   );
   gpc1_1 gpc1341 (
      {stage0_5[481]},
      {stage1_5[213]}
   );
   gpc1_1 gpc1342 (
      {stage0_5[482]},
      {stage1_5[214]}
   );
   gpc1_1 gpc1343 (
      {stage0_5[483]},
      {stage1_5[215]}
   );
   gpc1_1 gpc1344 (
      {stage0_5[484]},
      {stage1_5[216]}
   );
   gpc1_1 gpc1345 (
      {stage0_5[485]},
      {stage1_5[217]}
   );
   gpc1_1 gpc1346 (
      {stage0_6[410]},
      {stage1_6[171]}
   );
   gpc1_1 gpc1347 (
      {stage0_6[411]},
      {stage1_6[172]}
   );
   gpc1_1 gpc1348 (
      {stage0_6[412]},
      {stage1_6[173]}
   );
   gpc1_1 gpc1349 (
      {stage0_6[413]},
      {stage1_6[174]}
   );
   gpc1_1 gpc1350 (
      {stage0_6[414]},
      {stage1_6[175]}
   );
   gpc1_1 gpc1351 (
      {stage0_6[415]},
      {stage1_6[176]}
   );
   gpc1_1 gpc1352 (
      {stage0_6[416]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1353 (
      {stage0_6[417]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1354 (
      {stage0_6[418]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1355 (
      {stage0_6[419]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1356 (
      {stage0_6[420]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1357 (
      {stage0_6[421]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1358 (
      {stage0_6[422]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1359 (
      {stage0_6[423]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1360 (
      {stage0_6[424]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1361 (
      {stage0_6[425]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1362 (
      {stage0_6[426]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1363 (
      {stage0_6[427]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1364 (
      {stage0_6[428]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1365 (
      {stage0_6[429]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1366 (
      {stage0_6[430]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1367 (
      {stage0_6[431]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1368 (
      {stage0_6[432]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1369 (
      {stage0_6[433]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1370 (
      {stage0_6[434]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1371 (
      {stage0_6[435]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1372 (
      {stage0_6[436]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1373 (
      {stage0_6[437]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1374 (
      {stage0_6[438]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1375 (
      {stage0_6[439]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1376 (
      {stage0_6[440]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1377 (
      {stage0_6[441]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1378 (
      {stage0_6[442]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1379 (
      {stage0_6[443]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1380 (
      {stage0_6[444]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1381 (
      {stage0_6[445]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1382 (
      {stage0_6[446]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1383 (
      {stage0_6[447]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1384 (
      {stage0_6[448]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1385 (
      {stage0_6[449]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1386 (
      {stage0_6[450]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1387 (
      {stage0_6[451]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1388 (
      {stage0_6[452]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1389 (
      {stage0_6[453]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1390 (
      {stage0_6[454]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1391 (
      {stage0_6[455]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1392 (
      {stage0_6[456]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1393 (
      {stage0_6[457]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1394 (
      {stage0_6[458]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1395 (
      {stage0_6[459]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1396 (
      {stage0_6[460]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1397 (
      {stage0_6[461]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1398 (
      {stage0_6[462]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1399 (
      {stage0_6[463]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1400 (
      {stage0_6[464]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1401 (
      {stage0_6[465]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1402 (
      {stage0_6[466]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1403 (
      {stage0_6[467]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1404 (
      {stage0_6[468]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1405 (
      {stage0_6[469]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1406 (
      {stage0_6[470]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1407 (
      {stage0_6[471]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1408 (
      {stage0_6[472]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1409 (
      {stage0_6[473]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1410 (
      {stage0_6[474]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1411 (
      {stage0_6[475]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1412 (
      {stage0_6[476]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1413 (
      {stage0_6[477]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1414 (
      {stage0_6[478]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1415 (
      {stage0_6[479]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1416 (
      {stage0_6[480]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1417 (
      {stage0_6[481]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1418 (
      {stage0_6[482]},
      {stage1_6[243]}
   );
   gpc1_1 gpc1419 (
      {stage0_6[483]},
      {stage1_6[244]}
   );
   gpc1_1 gpc1420 (
      {stage0_6[484]},
      {stage1_6[245]}
   );
   gpc1_1 gpc1421 (
      {stage0_6[485]},
      {stage1_6[246]}
   );
   gpc1_1 gpc1422 (
      {stage0_7[436]},
      {stage1_7[174]}
   );
   gpc1_1 gpc1423 (
      {stage0_7[437]},
      {stage1_7[175]}
   );
   gpc1_1 gpc1424 (
      {stage0_7[438]},
      {stage1_7[176]}
   );
   gpc1_1 gpc1425 (
      {stage0_7[439]},
      {stage1_7[177]}
   );
   gpc1_1 gpc1426 (
      {stage0_7[440]},
      {stage1_7[178]}
   );
   gpc1_1 gpc1427 (
      {stage0_7[441]},
      {stage1_7[179]}
   );
   gpc1_1 gpc1428 (
      {stage0_7[442]},
      {stage1_7[180]}
   );
   gpc1_1 gpc1429 (
      {stage0_7[443]},
      {stage1_7[181]}
   );
   gpc1_1 gpc1430 (
      {stage0_7[444]},
      {stage1_7[182]}
   );
   gpc1_1 gpc1431 (
      {stage0_7[445]},
      {stage1_7[183]}
   );
   gpc1_1 gpc1432 (
      {stage0_7[446]},
      {stage1_7[184]}
   );
   gpc1_1 gpc1433 (
      {stage0_7[447]},
      {stage1_7[185]}
   );
   gpc1_1 gpc1434 (
      {stage0_7[448]},
      {stage1_7[186]}
   );
   gpc1_1 gpc1435 (
      {stage0_7[449]},
      {stage1_7[187]}
   );
   gpc1_1 gpc1436 (
      {stage0_7[450]},
      {stage1_7[188]}
   );
   gpc1_1 gpc1437 (
      {stage0_7[451]},
      {stage1_7[189]}
   );
   gpc1_1 gpc1438 (
      {stage0_7[452]},
      {stage1_7[190]}
   );
   gpc1_1 gpc1439 (
      {stage0_7[453]},
      {stage1_7[191]}
   );
   gpc1_1 gpc1440 (
      {stage0_7[454]},
      {stage1_7[192]}
   );
   gpc1_1 gpc1441 (
      {stage0_7[455]},
      {stage1_7[193]}
   );
   gpc1_1 gpc1442 (
      {stage0_7[456]},
      {stage1_7[194]}
   );
   gpc1_1 gpc1443 (
      {stage0_7[457]},
      {stage1_7[195]}
   );
   gpc1_1 gpc1444 (
      {stage0_7[458]},
      {stage1_7[196]}
   );
   gpc1_1 gpc1445 (
      {stage0_7[459]},
      {stage1_7[197]}
   );
   gpc1_1 gpc1446 (
      {stage0_7[460]},
      {stage1_7[198]}
   );
   gpc1_1 gpc1447 (
      {stage0_7[461]},
      {stage1_7[199]}
   );
   gpc1_1 gpc1448 (
      {stage0_7[462]},
      {stage1_7[200]}
   );
   gpc1_1 gpc1449 (
      {stage0_7[463]},
      {stage1_7[201]}
   );
   gpc1_1 gpc1450 (
      {stage0_7[464]},
      {stage1_7[202]}
   );
   gpc1_1 gpc1451 (
      {stage0_7[465]},
      {stage1_7[203]}
   );
   gpc1_1 gpc1452 (
      {stage0_7[466]},
      {stage1_7[204]}
   );
   gpc1_1 gpc1453 (
      {stage0_7[467]},
      {stage1_7[205]}
   );
   gpc1_1 gpc1454 (
      {stage0_7[468]},
      {stage1_7[206]}
   );
   gpc1_1 gpc1455 (
      {stage0_7[469]},
      {stage1_7[207]}
   );
   gpc1_1 gpc1456 (
      {stage0_7[470]},
      {stage1_7[208]}
   );
   gpc1_1 gpc1457 (
      {stage0_7[471]},
      {stage1_7[209]}
   );
   gpc1_1 gpc1458 (
      {stage0_7[472]},
      {stage1_7[210]}
   );
   gpc1_1 gpc1459 (
      {stage0_7[473]},
      {stage1_7[211]}
   );
   gpc1_1 gpc1460 (
      {stage0_7[474]},
      {stage1_7[212]}
   );
   gpc1_1 gpc1461 (
      {stage0_7[475]},
      {stage1_7[213]}
   );
   gpc1_1 gpc1462 (
      {stage0_7[476]},
      {stage1_7[214]}
   );
   gpc1_1 gpc1463 (
      {stage0_7[477]},
      {stage1_7[215]}
   );
   gpc1_1 gpc1464 (
      {stage0_7[478]},
      {stage1_7[216]}
   );
   gpc1_1 gpc1465 (
      {stage0_7[479]},
      {stage1_7[217]}
   );
   gpc1_1 gpc1466 (
      {stage0_7[480]},
      {stage1_7[218]}
   );
   gpc1_1 gpc1467 (
      {stage0_7[481]},
      {stage1_7[219]}
   );
   gpc1_1 gpc1468 (
      {stage0_7[482]},
      {stage1_7[220]}
   );
   gpc1_1 gpc1469 (
      {stage0_7[483]},
      {stage1_7[221]}
   );
   gpc1_1 gpc1470 (
      {stage0_7[484]},
      {stage1_7[222]}
   );
   gpc1_1 gpc1471 (
      {stage0_7[485]},
      {stage1_7[223]}
   );
   gpc1_1 gpc1472 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc1473 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc1474 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc1475 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1476 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1477 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1478 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc1479 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc1480 (
      {stage0_10[475]},
      {stage1_10[177]}
   );
   gpc1_1 gpc1481 (
      {stage0_10[476]},
      {stage1_10[178]}
   );
   gpc1_1 gpc1482 (
      {stage0_10[477]},
      {stage1_10[179]}
   );
   gpc1_1 gpc1483 (
      {stage0_10[478]},
      {stage1_10[180]}
   );
   gpc1_1 gpc1484 (
      {stage0_10[479]},
      {stage1_10[181]}
   );
   gpc1_1 gpc1485 (
      {stage0_10[480]},
      {stage1_10[182]}
   );
   gpc1_1 gpc1486 (
      {stage0_10[481]},
      {stage1_10[183]}
   );
   gpc1_1 gpc1487 (
      {stage0_10[482]},
      {stage1_10[184]}
   );
   gpc1_1 gpc1488 (
      {stage0_10[483]},
      {stage1_10[185]}
   );
   gpc1_1 gpc1489 (
      {stage0_10[484]},
      {stage1_10[186]}
   );
   gpc1_1 gpc1490 (
      {stage0_10[485]},
      {stage1_10[187]}
   );
   gpc1_1 gpc1491 (
      {stage0_11[451]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1492 (
      {stage0_11[452]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1493 (
      {stage0_11[453]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1494 (
      {stage0_11[454]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1495 (
      {stage0_11[455]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1496 (
      {stage0_11[456]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1497 (
      {stage0_11[457]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1498 (
      {stage0_11[458]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1499 (
      {stage0_11[459]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1500 (
      {stage0_11[460]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1501 (
      {stage0_11[461]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1502 (
      {stage0_11[462]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1503 (
      {stage0_11[463]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1504 (
      {stage0_11[464]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1505 (
      {stage0_11[465]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1506 (
      {stage0_11[466]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1507 (
      {stage0_11[467]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1508 (
      {stage0_11[468]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1509 (
      {stage0_11[469]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1510 (
      {stage0_11[470]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1511 (
      {stage0_11[471]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1512 (
      {stage0_11[472]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1513 (
      {stage0_11[473]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1514 (
      {stage0_11[474]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1515 (
      {stage0_11[475]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1516 (
      {stage0_11[476]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1517 (
      {stage0_11[477]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1518 (
      {stage0_11[478]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1519 (
      {stage0_11[479]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1520 (
      {stage0_11[480]},
      {stage1_11[214]}
   );
   gpc1_1 gpc1521 (
      {stage0_11[481]},
      {stage1_11[215]}
   );
   gpc1_1 gpc1522 (
      {stage0_11[482]},
      {stage1_11[216]}
   );
   gpc1_1 gpc1523 (
      {stage0_11[483]},
      {stage1_11[217]}
   );
   gpc1_1 gpc1524 (
      {stage0_11[484]},
      {stage1_11[218]}
   );
   gpc1_1 gpc1525 (
      {stage0_11[485]},
      {stage1_11[219]}
   );
   gpc1_1 gpc1526 (
      {stage0_12[408]},
      {stage1_12[204]}
   );
   gpc1_1 gpc1527 (
      {stage0_12[409]},
      {stage1_12[205]}
   );
   gpc1_1 gpc1528 (
      {stage0_12[410]},
      {stage1_12[206]}
   );
   gpc1_1 gpc1529 (
      {stage0_12[411]},
      {stage1_12[207]}
   );
   gpc1_1 gpc1530 (
      {stage0_12[412]},
      {stage1_12[208]}
   );
   gpc1_1 gpc1531 (
      {stage0_12[413]},
      {stage1_12[209]}
   );
   gpc1_1 gpc1532 (
      {stage0_12[414]},
      {stage1_12[210]}
   );
   gpc1_1 gpc1533 (
      {stage0_12[415]},
      {stage1_12[211]}
   );
   gpc1_1 gpc1534 (
      {stage0_12[416]},
      {stage1_12[212]}
   );
   gpc1_1 gpc1535 (
      {stage0_12[417]},
      {stage1_12[213]}
   );
   gpc1_1 gpc1536 (
      {stage0_12[418]},
      {stage1_12[214]}
   );
   gpc1_1 gpc1537 (
      {stage0_12[419]},
      {stage1_12[215]}
   );
   gpc1_1 gpc1538 (
      {stage0_12[420]},
      {stage1_12[216]}
   );
   gpc1_1 gpc1539 (
      {stage0_12[421]},
      {stage1_12[217]}
   );
   gpc1_1 gpc1540 (
      {stage0_12[422]},
      {stage1_12[218]}
   );
   gpc1_1 gpc1541 (
      {stage0_12[423]},
      {stage1_12[219]}
   );
   gpc1_1 gpc1542 (
      {stage0_12[424]},
      {stage1_12[220]}
   );
   gpc1_1 gpc1543 (
      {stage0_12[425]},
      {stage1_12[221]}
   );
   gpc1_1 gpc1544 (
      {stage0_12[426]},
      {stage1_12[222]}
   );
   gpc1_1 gpc1545 (
      {stage0_12[427]},
      {stage1_12[223]}
   );
   gpc1_1 gpc1546 (
      {stage0_12[428]},
      {stage1_12[224]}
   );
   gpc1_1 gpc1547 (
      {stage0_12[429]},
      {stage1_12[225]}
   );
   gpc1_1 gpc1548 (
      {stage0_12[430]},
      {stage1_12[226]}
   );
   gpc1_1 gpc1549 (
      {stage0_12[431]},
      {stage1_12[227]}
   );
   gpc1_1 gpc1550 (
      {stage0_12[432]},
      {stage1_12[228]}
   );
   gpc1_1 gpc1551 (
      {stage0_12[433]},
      {stage1_12[229]}
   );
   gpc1_1 gpc1552 (
      {stage0_12[434]},
      {stage1_12[230]}
   );
   gpc1_1 gpc1553 (
      {stage0_12[435]},
      {stage1_12[231]}
   );
   gpc1_1 gpc1554 (
      {stage0_12[436]},
      {stage1_12[232]}
   );
   gpc1_1 gpc1555 (
      {stage0_12[437]},
      {stage1_12[233]}
   );
   gpc1_1 gpc1556 (
      {stage0_12[438]},
      {stage1_12[234]}
   );
   gpc1_1 gpc1557 (
      {stage0_12[439]},
      {stage1_12[235]}
   );
   gpc1_1 gpc1558 (
      {stage0_12[440]},
      {stage1_12[236]}
   );
   gpc1_1 gpc1559 (
      {stage0_12[441]},
      {stage1_12[237]}
   );
   gpc1_1 gpc1560 (
      {stage0_12[442]},
      {stage1_12[238]}
   );
   gpc1_1 gpc1561 (
      {stage0_12[443]},
      {stage1_12[239]}
   );
   gpc1_1 gpc1562 (
      {stage0_12[444]},
      {stage1_12[240]}
   );
   gpc1_1 gpc1563 (
      {stage0_12[445]},
      {stage1_12[241]}
   );
   gpc1_1 gpc1564 (
      {stage0_12[446]},
      {stage1_12[242]}
   );
   gpc1_1 gpc1565 (
      {stage0_12[447]},
      {stage1_12[243]}
   );
   gpc1_1 gpc1566 (
      {stage0_12[448]},
      {stage1_12[244]}
   );
   gpc1_1 gpc1567 (
      {stage0_12[449]},
      {stage1_12[245]}
   );
   gpc1_1 gpc1568 (
      {stage0_12[450]},
      {stage1_12[246]}
   );
   gpc1_1 gpc1569 (
      {stage0_12[451]},
      {stage1_12[247]}
   );
   gpc1_1 gpc1570 (
      {stage0_12[452]},
      {stage1_12[248]}
   );
   gpc1_1 gpc1571 (
      {stage0_12[453]},
      {stage1_12[249]}
   );
   gpc1_1 gpc1572 (
      {stage0_12[454]},
      {stage1_12[250]}
   );
   gpc1_1 gpc1573 (
      {stage0_12[455]},
      {stage1_12[251]}
   );
   gpc1_1 gpc1574 (
      {stage0_12[456]},
      {stage1_12[252]}
   );
   gpc1_1 gpc1575 (
      {stage0_12[457]},
      {stage1_12[253]}
   );
   gpc1_1 gpc1576 (
      {stage0_12[458]},
      {stage1_12[254]}
   );
   gpc1_1 gpc1577 (
      {stage0_12[459]},
      {stage1_12[255]}
   );
   gpc1_1 gpc1578 (
      {stage0_12[460]},
      {stage1_12[256]}
   );
   gpc1_1 gpc1579 (
      {stage0_12[461]},
      {stage1_12[257]}
   );
   gpc1_1 gpc1580 (
      {stage0_12[462]},
      {stage1_12[258]}
   );
   gpc1_1 gpc1581 (
      {stage0_12[463]},
      {stage1_12[259]}
   );
   gpc1_1 gpc1582 (
      {stage0_12[464]},
      {stage1_12[260]}
   );
   gpc1_1 gpc1583 (
      {stage0_12[465]},
      {stage1_12[261]}
   );
   gpc1_1 gpc1584 (
      {stage0_12[466]},
      {stage1_12[262]}
   );
   gpc1_1 gpc1585 (
      {stage0_12[467]},
      {stage1_12[263]}
   );
   gpc1_1 gpc1586 (
      {stage0_12[468]},
      {stage1_12[264]}
   );
   gpc1_1 gpc1587 (
      {stage0_12[469]},
      {stage1_12[265]}
   );
   gpc1_1 gpc1588 (
      {stage0_12[470]},
      {stage1_12[266]}
   );
   gpc1_1 gpc1589 (
      {stage0_12[471]},
      {stage1_12[267]}
   );
   gpc1_1 gpc1590 (
      {stage0_12[472]},
      {stage1_12[268]}
   );
   gpc1_1 gpc1591 (
      {stage0_12[473]},
      {stage1_12[269]}
   );
   gpc1_1 gpc1592 (
      {stage0_12[474]},
      {stage1_12[270]}
   );
   gpc1_1 gpc1593 (
      {stage0_12[475]},
      {stage1_12[271]}
   );
   gpc1_1 gpc1594 (
      {stage0_12[476]},
      {stage1_12[272]}
   );
   gpc1_1 gpc1595 (
      {stage0_12[477]},
      {stage1_12[273]}
   );
   gpc1_1 gpc1596 (
      {stage0_12[478]},
      {stage1_12[274]}
   );
   gpc1_1 gpc1597 (
      {stage0_12[479]},
      {stage1_12[275]}
   );
   gpc1_1 gpc1598 (
      {stage0_12[480]},
      {stage1_12[276]}
   );
   gpc1_1 gpc1599 (
      {stage0_12[481]},
      {stage1_12[277]}
   );
   gpc1_1 gpc1600 (
      {stage0_12[482]},
      {stage1_12[278]}
   );
   gpc1_1 gpc1601 (
      {stage0_12[483]},
      {stage1_12[279]}
   );
   gpc1_1 gpc1602 (
      {stage0_12[484]},
      {stage1_12[280]}
   );
   gpc1_1 gpc1603 (
      {stage0_12[485]},
      {stage1_12[281]}
   );
   gpc1_1 gpc1604 (
      {stage0_13[476]},
      {stage1_13[195]}
   );
   gpc1_1 gpc1605 (
      {stage0_13[477]},
      {stage1_13[196]}
   );
   gpc1_1 gpc1606 (
      {stage0_13[478]},
      {stage1_13[197]}
   );
   gpc1_1 gpc1607 (
      {stage0_13[479]},
      {stage1_13[198]}
   );
   gpc1_1 gpc1608 (
      {stage0_13[480]},
      {stage1_13[199]}
   );
   gpc1_1 gpc1609 (
      {stage0_13[481]},
      {stage1_13[200]}
   );
   gpc1_1 gpc1610 (
      {stage0_13[482]},
      {stage1_13[201]}
   );
   gpc1_1 gpc1611 (
      {stage0_13[483]},
      {stage1_13[202]}
   );
   gpc1_1 gpc1612 (
      {stage0_13[484]},
      {stage1_13[203]}
   );
   gpc1_1 gpc1613 (
      {stage0_13[485]},
      {stage1_13[204]}
   );
   gpc1_1 gpc1614 (
      {stage0_14[349]},
      {stage1_14[160]}
   );
   gpc1_1 gpc1615 (
      {stage0_14[350]},
      {stage1_14[161]}
   );
   gpc1_1 gpc1616 (
      {stage0_14[351]},
      {stage1_14[162]}
   );
   gpc1_1 gpc1617 (
      {stage0_14[352]},
      {stage1_14[163]}
   );
   gpc1_1 gpc1618 (
      {stage0_14[353]},
      {stage1_14[164]}
   );
   gpc1_1 gpc1619 (
      {stage0_14[354]},
      {stage1_14[165]}
   );
   gpc1_1 gpc1620 (
      {stage0_14[355]},
      {stage1_14[166]}
   );
   gpc1_1 gpc1621 (
      {stage0_14[356]},
      {stage1_14[167]}
   );
   gpc1_1 gpc1622 (
      {stage0_14[357]},
      {stage1_14[168]}
   );
   gpc1_1 gpc1623 (
      {stage0_14[358]},
      {stage1_14[169]}
   );
   gpc1_1 gpc1624 (
      {stage0_14[359]},
      {stage1_14[170]}
   );
   gpc1_1 gpc1625 (
      {stage0_14[360]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1626 (
      {stage0_14[361]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1627 (
      {stage0_14[362]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1628 (
      {stage0_14[363]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1629 (
      {stage0_14[364]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1630 (
      {stage0_14[365]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1631 (
      {stage0_14[366]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1632 (
      {stage0_14[367]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1633 (
      {stage0_14[368]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1634 (
      {stage0_14[369]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1635 (
      {stage0_14[370]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1636 (
      {stage0_14[371]},
      {stage1_14[182]}
   );
   gpc1_1 gpc1637 (
      {stage0_14[372]},
      {stage1_14[183]}
   );
   gpc1_1 gpc1638 (
      {stage0_14[373]},
      {stage1_14[184]}
   );
   gpc1_1 gpc1639 (
      {stage0_14[374]},
      {stage1_14[185]}
   );
   gpc1_1 gpc1640 (
      {stage0_14[375]},
      {stage1_14[186]}
   );
   gpc1_1 gpc1641 (
      {stage0_14[376]},
      {stage1_14[187]}
   );
   gpc1_1 gpc1642 (
      {stage0_14[377]},
      {stage1_14[188]}
   );
   gpc1_1 gpc1643 (
      {stage0_14[378]},
      {stage1_14[189]}
   );
   gpc1_1 gpc1644 (
      {stage0_14[379]},
      {stage1_14[190]}
   );
   gpc1_1 gpc1645 (
      {stage0_14[380]},
      {stage1_14[191]}
   );
   gpc1_1 gpc1646 (
      {stage0_14[381]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1647 (
      {stage0_14[382]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1648 (
      {stage0_14[383]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1649 (
      {stage0_14[384]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1650 (
      {stage0_14[385]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1651 (
      {stage0_14[386]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1652 (
      {stage0_14[387]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1653 (
      {stage0_14[388]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1654 (
      {stage0_14[389]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1655 (
      {stage0_14[390]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1656 (
      {stage0_14[391]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1657 (
      {stage0_14[392]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1658 (
      {stage0_14[393]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1659 (
      {stage0_14[394]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1660 (
      {stage0_14[395]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1661 (
      {stage0_14[396]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1662 (
      {stage0_14[397]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1663 (
      {stage0_14[398]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1664 (
      {stage0_14[399]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1665 (
      {stage0_14[400]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1666 (
      {stage0_14[401]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1667 (
      {stage0_14[402]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1668 (
      {stage0_14[403]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1669 (
      {stage0_14[404]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1670 (
      {stage0_14[405]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1671 (
      {stage0_14[406]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1672 (
      {stage0_14[407]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1673 (
      {stage0_14[408]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1674 (
      {stage0_14[409]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1675 (
      {stage0_14[410]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1676 (
      {stage0_14[411]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1677 (
      {stage0_14[412]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1678 (
      {stage0_14[413]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1679 (
      {stage0_14[414]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1680 (
      {stage0_14[415]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1681 (
      {stage0_14[416]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1682 (
      {stage0_14[417]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1683 (
      {stage0_14[418]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1684 (
      {stage0_14[419]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1685 (
      {stage0_14[420]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1686 (
      {stage0_14[421]},
      {stage1_14[232]}
   );
   gpc1_1 gpc1687 (
      {stage0_14[422]},
      {stage1_14[233]}
   );
   gpc1_1 gpc1688 (
      {stage0_14[423]},
      {stage1_14[234]}
   );
   gpc1_1 gpc1689 (
      {stage0_14[424]},
      {stage1_14[235]}
   );
   gpc1_1 gpc1690 (
      {stage0_14[425]},
      {stage1_14[236]}
   );
   gpc1_1 gpc1691 (
      {stage0_14[426]},
      {stage1_14[237]}
   );
   gpc1_1 gpc1692 (
      {stage0_14[427]},
      {stage1_14[238]}
   );
   gpc1_1 gpc1693 (
      {stage0_14[428]},
      {stage1_14[239]}
   );
   gpc1_1 gpc1694 (
      {stage0_14[429]},
      {stage1_14[240]}
   );
   gpc1_1 gpc1695 (
      {stage0_14[430]},
      {stage1_14[241]}
   );
   gpc1_1 gpc1696 (
      {stage0_14[431]},
      {stage1_14[242]}
   );
   gpc1_1 gpc1697 (
      {stage0_14[432]},
      {stage1_14[243]}
   );
   gpc1_1 gpc1698 (
      {stage0_14[433]},
      {stage1_14[244]}
   );
   gpc1_1 gpc1699 (
      {stage0_14[434]},
      {stage1_14[245]}
   );
   gpc1_1 gpc1700 (
      {stage0_14[435]},
      {stage1_14[246]}
   );
   gpc1_1 gpc1701 (
      {stage0_14[436]},
      {stage1_14[247]}
   );
   gpc1_1 gpc1702 (
      {stage0_14[437]},
      {stage1_14[248]}
   );
   gpc1_1 gpc1703 (
      {stage0_14[438]},
      {stage1_14[249]}
   );
   gpc1_1 gpc1704 (
      {stage0_14[439]},
      {stage1_14[250]}
   );
   gpc1_1 gpc1705 (
      {stage0_14[440]},
      {stage1_14[251]}
   );
   gpc1_1 gpc1706 (
      {stage0_14[441]},
      {stage1_14[252]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[442]},
      {stage1_14[253]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[443]},
      {stage1_14[254]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[444]},
      {stage1_14[255]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[445]},
      {stage1_14[256]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[446]},
      {stage1_14[257]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[447]},
      {stage1_14[258]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[448]},
      {stage1_14[259]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[449]},
      {stage1_14[260]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[450]},
      {stage1_14[261]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[451]},
      {stage1_14[262]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[452]},
      {stage1_14[263]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[453]},
      {stage1_14[264]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[454]},
      {stage1_14[265]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[455]},
      {stage1_14[266]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[456]},
      {stage1_14[267]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[457]},
      {stage1_14[268]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[458]},
      {stage1_14[269]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[459]},
      {stage1_14[270]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[460]},
      {stage1_14[271]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[461]},
      {stage1_14[272]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[462]},
      {stage1_14[273]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[463]},
      {stage1_14[274]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[464]},
      {stage1_14[275]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[465]},
      {stage1_14[276]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[466]},
      {stage1_14[277]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[467]},
      {stage1_14[278]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[468]},
      {stage1_14[279]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[469]},
      {stage1_14[280]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[470]},
      {stage1_14[281]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[471]},
      {stage1_14[282]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[472]},
      {stage1_14[283]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[473]},
      {stage1_14[284]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[474]},
      {stage1_14[285]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[475]},
      {stage1_14[286]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[476]},
      {stage1_14[287]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[477]},
      {stage1_14[288]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[478]},
      {stage1_14[289]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[479]},
      {stage1_14[290]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[480]},
      {stage1_14[291]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[481]},
      {stage1_14[292]}
   );
   gpc1_1 gpc1747 (
      {stage0_14[482]},
      {stage1_14[293]}
   );
   gpc1_1 gpc1748 (
      {stage0_14[483]},
      {stage1_14[294]}
   );
   gpc1_1 gpc1749 (
      {stage0_14[484]},
      {stage1_14[295]}
   );
   gpc1_1 gpc1750 (
      {stage0_14[485]},
      {stage1_14[296]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[480]},
      {stage1_15[166]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[481]},
      {stage1_15[167]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[482]},
      {stage1_15[168]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[483]},
      {stage1_15[169]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[484]},
      {stage1_15[170]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[485]},
      {stage1_15[171]}
   );
   gpc1_1 gpc1757 (
      {stage0_16[411]},
      {stage1_16[190]}
   );
   gpc1_1 gpc1758 (
      {stage0_16[412]},
      {stage1_16[191]}
   );
   gpc1_1 gpc1759 (
      {stage0_16[413]},
      {stage1_16[192]}
   );
   gpc1_1 gpc1760 (
      {stage0_16[414]},
      {stage1_16[193]}
   );
   gpc1_1 gpc1761 (
      {stage0_16[415]},
      {stage1_16[194]}
   );
   gpc1_1 gpc1762 (
      {stage0_16[416]},
      {stage1_16[195]}
   );
   gpc1_1 gpc1763 (
      {stage0_16[417]},
      {stage1_16[196]}
   );
   gpc1_1 gpc1764 (
      {stage0_16[418]},
      {stage1_16[197]}
   );
   gpc1_1 gpc1765 (
      {stage0_16[419]},
      {stage1_16[198]}
   );
   gpc1_1 gpc1766 (
      {stage0_16[420]},
      {stage1_16[199]}
   );
   gpc1_1 gpc1767 (
      {stage0_16[421]},
      {stage1_16[200]}
   );
   gpc1_1 gpc1768 (
      {stage0_16[422]},
      {stage1_16[201]}
   );
   gpc1_1 gpc1769 (
      {stage0_16[423]},
      {stage1_16[202]}
   );
   gpc1_1 gpc1770 (
      {stage0_16[424]},
      {stage1_16[203]}
   );
   gpc1_1 gpc1771 (
      {stage0_16[425]},
      {stage1_16[204]}
   );
   gpc1_1 gpc1772 (
      {stage0_16[426]},
      {stage1_16[205]}
   );
   gpc1_1 gpc1773 (
      {stage0_16[427]},
      {stage1_16[206]}
   );
   gpc1_1 gpc1774 (
      {stage0_16[428]},
      {stage1_16[207]}
   );
   gpc1_1 gpc1775 (
      {stage0_16[429]},
      {stage1_16[208]}
   );
   gpc1_1 gpc1776 (
      {stage0_16[430]},
      {stage1_16[209]}
   );
   gpc1_1 gpc1777 (
      {stage0_16[431]},
      {stage1_16[210]}
   );
   gpc1_1 gpc1778 (
      {stage0_16[432]},
      {stage1_16[211]}
   );
   gpc1_1 gpc1779 (
      {stage0_16[433]},
      {stage1_16[212]}
   );
   gpc1_1 gpc1780 (
      {stage0_16[434]},
      {stage1_16[213]}
   );
   gpc1_1 gpc1781 (
      {stage0_16[435]},
      {stage1_16[214]}
   );
   gpc1_1 gpc1782 (
      {stage0_16[436]},
      {stage1_16[215]}
   );
   gpc1_1 gpc1783 (
      {stage0_16[437]},
      {stage1_16[216]}
   );
   gpc1_1 gpc1784 (
      {stage0_16[438]},
      {stage1_16[217]}
   );
   gpc1_1 gpc1785 (
      {stage0_16[439]},
      {stage1_16[218]}
   );
   gpc1_1 gpc1786 (
      {stage0_16[440]},
      {stage1_16[219]}
   );
   gpc1_1 gpc1787 (
      {stage0_16[441]},
      {stage1_16[220]}
   );
   gpc1_1 gpc1788 (
      {stage0_16[442]},
      {stage1_16[221]}
   );
   gpc1_1 gpc1789 (
      {stage0_16[443]},
      {stage1_16[222]}
   );
   gpc1_1 gpc1790 (
      {stage0_16[444]},
      {stage1_16[223]}
   );
   gpc1_1 gpc1791 (
      {stage0_16[445]},
      {stage1_16[224]}
   );
   gpc1_1 gpc1792 (
      {stage0_16[446]},
      {stage1_16[225]}
   );
   gpc1_1 gpc1793 (
      {stage0_16[447]},
      {stage1_16[226]}
   );
   gpc1_1 gpc1794 (
      {stage0_16[448]},
      {stage1_16[227]}
   );
   gpc1_1 gpc1795 (
      {stage0_16[449]},
      {stage1_16[228]}
   );
   gpc1_1 gpc1796 (
      {stage0_16[450]},
      {stage1_16[229]}
   );
   gpc1_1 gpc1797 (
      {stage0_16[451]},
      {stage1_16[230]}
   );
   gpc1_1 gpc1798 (
      {stage0_16[452]},
      {stage1_16[231]}
   );
   gpc1_1 gpc1799 (
      {stage0_16[453]},
      {stage1_16[232]}
   );
   gpc1_1 gpc1800 (
      {stage0_16[454]},
      {stage1_16[233]}
   );
   gpc1_1 gpc1801 (
      {stage0_16[455]},
      {stage1_16[234]}
   );
   gpc1_1 gpc1802 (
      {stage0_16[456]},
      {stage1_16[235]}
   );
   gpc1_1 gpc1803 (
      {stage0_16[457]},
      {stage1_16[236]}
   );
   gpc1_1 gpc1804 (
      {stage0_16[458]},
      {stage1_16[237]}
   );
   gpc1_1 gpc1805 (
      {stage0_16[459]},
      {stage1_16[238]}
   );
   gpc1_1 gpc1806 (
      {stage0_16[460]},
      {stage1_16[239]}
   );
   gpc1_1 gpc1807 (
      {stage0_16[461]},
      {stage1_16[240]}
   );
   gpc1_1 gpc1808 (
      {stage0_16[462]},
      {stage1_16[241]}
   );
   gpc1_1 gpc1809 (
      {stage0_16[463]},
      {stage1_16[242]}
   );
   gpc1_1 gpc1810 (
      {stage0_16[464]},
      {stage1_16[243]}
   );
   gpc1_1 gpc1811 (
      {stage0_16[465]},
      {stage1_16[244]}
   );
   gpc1_1 gpc1812 (
      {stage0_16[466]},
      {stage1_16[245]}
   );
   gpc1_1 gpc1813 (
      {stage0_16[467]},
      {stage1_16[246]}
   );
   gpc1_1 gpc1814 (
      {stage0_16[468]},
      {stage1_16[247]}
   );
   gpc1_1 gpc1815 (
      {stage0_16[469]},
      {stage1_16[248]}
   );
   gpc1_1 gpc1816 (
      {stage0_16[470]},
      {stage1_16[249]}
   );
   gpc1_1 gpc1817 (
      {stage0_16[471]},
      {stage1_16[250]}
   );
   gpc1_1 gpc1818 (
      {stage0_16[472]},
      {stage1_16[251]}
   );
   gpc1_1 gpc1819 (
      {stage0_16[473]},
      {stage1_16[252]}
   );
   gpc1_1 gpc1820 (
      {stage0_16[474]},
      {stage1_16[253]}
   );
   gpc1_1 gpc1821 (
      {stage0_16[475]},
      {stage1_16[254]}
   );
   gpc1_1 gpc1822 (
      {stage0_16[476]},
      {stage1_16[255]}
   );
   gpc1_1 gpc1823 (
      {stage0_16[477]},
      {stage1_16[256]}
   );
   gpc1_1 gpc1824 (
      {stage0_16[478]},
      {stage1_16[257]}
   );
   gpc1_1 gpc1825 (
      {stage0_16[479]},
      {stage1_16[258]}
   );
   gpc1_1 gpc1826 (
      {stage0_16[480]},
      {stage1_16[259]}
   );
   gpc1_1 gpc1827 (
      {stage0_16[481]},
      {stage1_16[260]}
   );
   gpc1_1 gpc1828 (
      {stage0_16[482]},
      {stage1_16[261]}
   );
   gpc1_1 gpc1829 (
      {stage0_16[483]},
      {stage1_16[262]}
   );
   gpc1_1 gpc1830 (
      {stage0_16[484]},
      {stage1_16[263]}
   );
   gpc1_1 gpc1831 (
      {stage0_16[485]},
      {stage1_16[264]}
   );
   gpc1_1 gpc1832 (
      {stage0_17[402]},
      {stage1_17[187]}
   );
   gpc1_1 gpc1833 (
      {stage0_17[403]},
      {stage1_17[188]}
   );
   gpc1_1 gpc1834 (
      {stage0_17[404]},
      {stage1_17[189]}
   );
   gpc1_1 gpc1835 (
      {stage0_17[405]},
      {stage1_17[190]}
   );
   gpc1_1 gpc1836 (
      {stage0_17[406]},
      {stage1_17[191]}
   );
   gpc1_1 gpc1837 (
      {stage0_17[407]},
      {stage1_17[192]}
   );
   gpc1_1 gpc1838 (
      {stage0_17[408]},
      {stage1_17[193]}
   );
   gpc1_1 gpc1839 (
      {stage0_17[409]},
      {stage1_17[194]}
   );
   gpc1_1 gpc1840 (
      {stage0_17[410]},
      {stage1_17[195]}
   );
   gpc1_1 gpc1841 (
      {stage0_17[411]},
      {stage1_17[196]}
   );
   gpc1_1 gpc1842 (
      {stage0_17[412]},
      {stage1_17[197]}
   );
   gpc1_1 gpc1843 (
      {stage0_17[413]},
      {stage1_17[198]}
   );
   gpc1_1 gpc1844 (
      {stage0_17[414]},
      {stage1_17[199]}
   );
   gpc1_1 gpc1845 (
      {stage0_17[415]},
      {stage1_17[200]}
   );
   gpc1_1 gpc1846 (
      {stage0_17[416]},
      {stage1_17[201]}
   );
   gpc1_1 gpc1847 (
      {stage0_17[417]},
      {stage1_17[202]}
   );
   gpc1_1 gpc1848 (
      {stage0_17[418]},
      {stage1_17[203]}
   );
   gpc1_1 gpc1849 (
      {stage0_17[419]},
      {stage1_17[204]}
   );
   gpc1_1 gpc1850 (
      {stage0_17[420]},
      {stage1_17[205]}
   );
   gpc1_1 gpc1851 (
      {stage0_17[421]},
      {stage1_17[206]}
   );
   gpc1_1 gpc1852 (
      {stage0_17[422]},
      {stage1_17[207]}
   );
   gpc1_1 gpc1853 (
      {stage0_17[423]},
      {stage1_17[208]}
   );
   gpc1_1 gpc1854 (
      {stage0_17[424]},
      {stage1_17[209]}
   );
   gpc1_1 gpc1855 (
      {stage0_17[425]},
      {stage1_17[210]}
   );
   gpc1_1 gpc1856 (
      {stage0_17[426]},
      {stage1_17[211]}
   );
   gpc1_1 gpc1857 (
      {stage0_17[427]},
      {stage1_17[212]}
   );
   gpc1_1 gpc1858 (
      {stage0_17[428]},
      {stage1_17[213]}
   );
   gpc1_1 gpc1859 (
      {stage0_17[429]},
      {stage1_17[214]}
   );
   gpc1_1 gpc1860 (
      {stage0_17[430]},
      {stage1_17[215]}
   );
   gpc1_1 gpc1861 (
      {stage0_17[431]},
      {stage1_17[216]}
   );
   gpc1_1 gpc1862 (
      {stage0_17[432]},
      {stage1_17[217]}
   );
   gpc1_1 gpc1863 (
      {stage0_17[433]},
      {stage1_17[218]}
   );
   gpc1_1 gpc1864 (
      {stage0_17[434]},
      {stage1_17[219]}
   );
   gpc1_1 gpc1865 (
      {stage0_17[435]},
      {stage1_17[220]}
   );
   gpc1_1 gpc1866 (
      {stage0_17[436]},
      {stage1_17[221]}
   );
   gpc1_1 gpc1867 (
      {stage0_17[437]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1868 (
      {stage0_17[438]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1869 (
      {stage0_17[439]},
      {stage1_17[224]}
   );
   gpc1_1 gpc1870 (
      {stage0_17[440]},
      {stage1_17[225]}
   );
   gpc1_1 gpc1871 (
      {stage0_17[441]},
      {stage1_17[226]}
   );
   gpc1_1 gpc1872 (
      {stage0_17[442]},
      {stage1_17[227]}
   );
   gpc1_1 gpc1873 (
      {stage0_17[443]},
      {stage1_17[228]}
   );
   gpc1_1 gpc1874 (
      {stage0_17[444]},
      {stage1_17[229]}
   );
   gpc1_1 gpc1875 (
      {stage0_17[445]},
      {stage1_17[230]}
   );
   gpc1_1 gpc1876 (
      {stage0_17[446]},
      {stage1_17[231]}
   );
   gpc1_1 gpc1877 (
      {stage0_17[447]},
      {stage1_17[232]}
   );
   gpc1_1 gpc1878 (
      {stage0_17[448]},
      {stage1_17[233]}
   );
   gpc1_1 gpc1879 (
      {stage0_17[449]},
      {stage1_17[234]}
   );
   gpc1_1 gpc1880 (
      {stage0_17[450]},
      {stage1_17[235]}
   );
   gpc1_1 gpc1881 (
      {stage0_17[451]},
      {stage1_17[236]}
   );
   gpc1_1 gpc1882 (
      {stage0_17[452]},
      {stage1_17[237]}
   );
   gpc1_1 gpc1883 (
      {stage0_17[453]},
      {stage1_17[238]}
   );
   gpc1_1 gpc1884 (
      {stage0_17[454]},
      {stage1_17[239]}
   );
   gpc1_1 gpc1885 (
      {stage0_17[455]},
      {stage1_17[240]}
   );
   gpc1_1 gpc1886 (
      {stage0_17[456]},
      {stage1_17[241]}
   );
   gpc1_1 gpc1887 (
      {stage0_17[457]},
      {stage1_17[242]}
   );
   gpc1_1 gpc1888 (
      {stage0_17[458]},
      {stage1_17[243]}
   );
   gpc1_1 gpc1889 (
      {stage0_17[459]},
      {stage1_17[244]}
   );
   gpc1_1 gpc1890 (
      {stage0_17[460]},
      {stage1_17[245]}
   );
   gpc1_1 gpc1891 (
      {stage0_17[461]},
      {stage1_17[246]}
   );
   gpc1_1 gpc1892 (
      {stage0_17[462]},
      {stage1_17[247]}
   );
   gpc1_1 gpc1893 (
      {stage0_17[463]},
      {stage1_17[248]}
   );
   gpc1_1 gpc1894 (
      {stage0_17[464]},
      {stage1_17[249]}
   );
   gpc1_1 gpc1895 (
      {stage0_17[465]},
      {stage1_17[250]}
   );
   gpc1_1 gpc1896 (
      {stage0_17[466]},
      {stage1_17[251]}
   );
   gpc1_1 gpc1897 (
      {stage0_17[467]},
      {stage1_17[252]}
   );
   gpc1_1 gpc1898 (
      {stage0_17[468]},
      {stage1_17[253]}
   );
   gpc1_1 gpc1899 (
      {stage0_17[469]},
      {stage1_17[254]}
   );
   gpc1_1 gpc1900 (
      {stage0_17[470]},
      {stage1_17[255]}
   );
   gpc1_1 gpc1901 (
      {stage0_17[471]},
      {stage1_17[256]}
   );
   gpc1_1 gpc1902 (
      {stage0_17[472]},
      {stage1_17[257]}
   );
   gpc1_1 gpc1903 (
      {stage0_17[473]},
      {stage1_17[258]}
   );
   gpc1_1 gpc1904 (
      {stage0_17[474]},
      {stage1_17[259]}
   );
   gpc1_1 gpc1905 (
      {stage0_17[475]},
      {stage1_17[260]}
   );
   gpc1_1 gpc1906 (
      {stage0_17[476]},
      {stage1_17[261]}
   );
   gpc1_1 gpc1907 (
      {stage0_17[477]},
      {stage1_17[262]}
   );
   gpc1_1 gpc1908 (
      {stage0_17[478]},
      {stage1_17[263]}
   );
   gpc1_1 gpc1909 (
      {stage0_17[479]},
      {stage1_17[264]}
   );
   gpc1_1 gpc1910 (
      {stage0_17[480]},
      {stage1_17[265]}
   );
   gpc1_1 gpc1911 (
      {stage0_17[481]},
      {stage1_17[266]}
   );
   gpc1_1 gpc1912 (
      {stage0_17[482]},
      {stage1_17[267]}
   );
   gpc1_1 gpc1913 (
      {stage0_17[483]},
      {stage1_17[268]}
   );
   gpc1_1 gpc1914 (
      {stage0_17[484]},
      {stage1_17[269]}
   );
   gpc1_1 gpc1915 (
      {stage0_17[485]},
      {stage1_17[270]}
   );
   gpc1_1 gpc1916 (
      {stage0_18[447]},
      {stage1_18[162]}
   );
   gpc1_1 gpc1917 (
      {stage0_18[448]},
      {stage1_18[163]}
   );
   gpc1_1 gpc1918 (
      {stage0_18[449]},
      {stage1_18[164]}
   );
   gpc1_1 gpc1919 (
      {stage0_18[450]},
      {stage1_18[165]}
   );
   gpc1_1 gpc1920 (
      {stage0_18[451]},
      {stage1_18[166]}
   );
   gpc1_1 gpc1921 (
      {stage0_18[452]},
      {stage1_18[167]}
   );
   gpc1_1 gpc1922 (
      {stage0_18[453]},
      {stage1_18[168]}
   );
   gpc1_1 gpc1923 (
      {stage0_18[454]},
      {stage1_18[169]}
   );
   gpc1_1 gpc1924 (
      {stage0_18[455]},
      {stage1_18[170]}
   );
   gpc1_1 gpc1925 (
      {stage0_18[456]},
      {stage1_18[171]}
   );
   gpc1_1 gpc1926 (
      {stage0_18[457]},
      {stage1_18[172]}
   );
   gpc1_1 gpc1927 (
      {stage0_18[458]},
      {stage1_18[173]}
   );
   gpc1_1 gpc1928 (
      {stage0_18[459]},
      {stage1_18[174]}
   );
   gpc1_1 gpc1929 (
      {stage0_18[460]},
      {stage1_18[175]}
   );
   gpc1_1 gpc1930 (
      {stage0_18[461]},
      {stage1_18[176]}
   );
   gpc1_1 gpc1931 (
      {stage0_18[462]},
      {stage1_18[177]}
   );
   gpc1_1 gpc1932 (
      {stage0_18[463]},
      {stage1_18[178]}
   );
   gpc1_1 gpc1933 (
      {stage0_18[464]},
      {stage1_18[179]}
   );
   gpc1_1 gpc1934 (
      {stage0_18[465]},
      {stage1_18[180]}
   );
   gpc1_1 gpc1935 (
      {stage0_18[466]},
      {stage1_18[181]}
   );
   gpc1_1 gpc1936 (
      {stage0_18[467]},
      {stage1_18[182]}
   );
   gpc1_1 gpc1937 (
      {stage0_18[468]},
      {stage1_18[183]}
   );
   gpc1_1 gpc1938 (
      {stage0_18[469]},
      {stage1_18[184]}
   );
   gpc1_1 gpc1939 (
      {stage0_18[470]},
      {stage1_18[185]}
   );
   gpc1_1 gpc1940 (
      {stage0_18[471]},
      {stage1_18[186]}
   );
   gpc1_1 gpc1941 (
      {stage0_18[472]},
      {stage1_18[187]}
   );
   gpc1_1 gpc1942 (
      {stage0_18[473]},
      {stage1_18[188]}
   );
   gpc1_1 gpc1943 (
      {stage0_18[474]},
      {stage1_18[189]}
   );
   gpc1_1 gpc1944 (
      {stage0_18[475]},
      {stage1_18[190]}
   );
   gpc1_1 gpc1945 (
      {stage0_18[476]},
      {stage1_18[191]}
   );
   gpc1_1 gpc1946 (
      {stage0_18[477]},
      {stage1_18[192]}
   );
   gpc1_1 gpc1947 (
      {stage0_18[478]},
      {stage1_18[193]}
   );
   gpc1_1 gpc1948 (
      {stage0_18[479]},
      {stage1_18[194]}
   );
   gpc1_1 gpc1949 (
      {stage0_18[480]},
      {stage1_18[195]}
   );
   gpc1_1 gpc1950 (
      {stage0_18[481]},
      {stage1_18[196]}
   );
   gpc1_1 gpc1951 (
      {stage0_18[482]},
      {stage1_18[197]}
   );
   gpc1_1 gpc1952 (
      {stage0_18[483]},
      {stage1_18[198]}
   );
   gpc1_1 gpc1953 (
      {stage0_18[484]},
      {stage1_18[199]}
   );
   gpc1_1 gpc1954 (
      {stage0_18[485]},
      {stage1_18[200]}
   );
   gpc1_1 gpc1955 (
      {stage0_19[347]},
      {stage1_19[161]}
   );
   gpc1_1 gpc1956 (
      {stage0_19[348]},
      {stage1_19[162]}
   );
   gpc1_1 gpc1957 (
      {stage0_19[349]},
      {stage1_19[163]}
   );
   gpc1_1 gpc1958 (
      {stage0_19[350]},
      {stage1_19[164]}
   );
   gpc1_1 gpc1959 (
      {stage0_19[351]},
      {stage1_19[165]}
   );
   gpc1_1 gpc1960 (
      {stage0_19[352]},
      {stage1_19[166]}
   );
   gpc1_1 gpc1961 (
      {stage0_19[353]},
      {stage1_19[167]}
   );
   gpc1_1 gpc1962 (
      {stage0_19[354]},
      {stage1_19[168]}
   );
   gpc1_1 gpc1963 (
      {stage0_19[355]},
      {stage1_19[169]}
   );
   gpc1_1 gpc1964 (
      {stage0_19[356]},
      {stage1_19[170]}
   );
   gpc1_1 gpc1965 (
      {stage0_19[357]},
      {stage1_19[171]}
   );
   gpc1_1 gpc1966 (
      {stage0_19[358]},
      {stage1_19[172]}
   );
   gpc1_1 gpc1967 (
      {stage0_19[359]},
      {stage1_19[173]}
   );
   gpc1_1 gpc1968 (
      {stage0_19[360]},
      {stage1_19[174]}
   );
   gpc1_1 gpc1969 (
      {stage0_19[361]},
      {stage1_19[175]}
   );
   gpc1_1 gpc1970 (
      {stage0_19[362]},
      {stage1_19[176]}
   );
   gpc1_1 gpc1971 (
      {stage0_19[363]},
      {stage1_19[177]}
   );
   gpc1_1 gpc1972 (
      {stage0_19[364]},
      {stage1_19[178]}
   );
   gpc1_1 gpc1973 (
      {stage0_19[365]},
      {stage1_19[179]}
   );
   gpc1_1 gpc1974 (
      {stage0_19[366]},
      {stage1_19[180]}
   );
   gpc1_1 gpc1975 (
      {stage0_19[367]},
      {stage1_19[181]}
   );
   gpc1_1 gpc1976 (
      {stage0_19[368]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1977 (
      {stage0_19[369]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1978 (
      {stage0_19[370]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1979 (
      {stage0_19[371]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1980 (
      {stage0_19[372]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1981 (
      {stage0_19[373]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1982 (
      {stage0_19[374]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1983 (
      {stage0_19[375]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1984 (
      {stage0_19[376]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1985 (
      {stage0_19[377]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1986 (
      {stage0_19[378]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1987 (
      {stage0_19[379]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1988 (
      {stage0_19[380]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1989 (
      {stage0_19[381]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1990 (
      {stage0_19[382]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1991 (
      {stage0_19[383]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1992 (
      {stage0_19[384]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1993 (
      {stage0_19[385]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1994 (
      {stage0_19[386]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1995 (
      {stage0_19[387]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1996 (
      {stage0_19[388]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1997 (
      {stage0_19[389]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1998 (
      {stage0_19[390]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1999 (
      {stage0_19[391]},
      {stage1_19[205]}
   );
   gpc1_1 gpc2000 (
      {stage0_19[392]},
      {stage1_19[206]}
   );
   gpc1_1 gpc2001 (
      {stage0_19[393]},
      {stage1_19[207]}
   );
   gpc1_1 gpc2002 (
      {stage0_19[394]},
      {stage1_19[208]}
   );
   gpc1_1 gpc2003 (
      {stage0_19[395]},
      {stage1_19[209]}
   );
   gpc1_1 gpc2004 (
      {stage0_19[396]},
      {stage1_19[210]}
   );
   gpc1_1 gpc2005 (
      {stage0_19[397]},
      {stage1_19[211]}
   );
   gpc1_1 gpc2006 (
      {stage0_19[398]},
      {stage1_19[212]}
   );
   gpc1_1 gpc2007 (
      {stage0_19[399]},
      {stage1_19[213]}
   );
   gpc1_1 gpc2008 (
      {stage0_19[400]},
      {stage1_19[214]}
   );
   gpc1_1 gpc2009 (
      {stage0_19[401]},
      {stage1_19[215]}
   );
   gpc1_1 gpc2010 (
      {stage0_19[402]},
      {stage1_19[216]}
   );
   gpc1_1 gpc2011 (
      {stage0_19[403]},
      {stage1_19[217]}
   );
   gpc1_1 gpc2012 (
      {stage0_19[404]},
      {stage1_19[218]}
   );
   gpc1_1 gpc2013 (
      {stage0_19[405]},
      {stage1_19[219]}
   );
   gpc1_1 gpc2014 (
      {stage0_19[406]},
      {stage1_19[220]}
   );
   gpc1_1 gpc2015 (
      {stage0_19[407]},
      {stage1_19[221]}
   );
   gpc1_1 gpc2016 (
      {stage0_19[408]},
      {stage1_19[222]}
   );
   gpc1_1 gpc2017 (
      {stage0_19[409]},
      {stage1_19[223]}
   );
   gpc1_1 gpc2018 (
      {stage0_19[410]},
      {stage1_19[224]}
   );
   gpc1_1 gpc2019 (
      {stage0_19[411]},
      {stage1_19[225]}
   );
   gpc1_1 gpc2020 (
      {stage0_19[412]},
      {stage1_19[226]}
   );
   gpc1_1 gpc2021 (
      {stage0_19[413]},
      {stage1_19[227]}
   );
   gpc1_1 gpc2022 (
      {stage0_19[414]},
      {stage1_19[228]}
   );
   gpc1_1 gpc2023 (
      {stage0_19[415]},
      {stage1_19[229]}
   );
   gpc1_1 gpc2024 (
      {stage0_19[416]},
      {stage1_19[230]}
   );
   gpc1_1 gpc2025 (
      {stage0_19[417]},
      {stage1_19[231]}
   );
   gpc1_1 gpc2026 (
      {stage0_19[418]},
      {stage1_19[232]}
   );
   gpc1_1 gpc2027 (
      {stage0_19[419]},
      {stage1_19[233]}
   );
   gpc1_1 gpc2028 (
      {stage0_19[420]},
      {stage1_19[234]}
   );
   gpc1_1 gpc2029 (
      {stage0_19[421]},
      {stage1_19[235]}
   );
   gpc1_1 gpc2030 (
      {stage0_19[422]},
      {stage1_19[236]}
   );
   gpc1_1 gpc2031 (
      {stage0_19[423]},
      {stage1_19[237]}
   );
   gpc1_1 gpc2032 (
      {stage0_19[424]},
      {stage1_19[238]}
   );
   gpc1_1 gpc2033 (
      {stage0_19[425]},
      {stage1_19[239]}
   );
   gpc1_1 gpc2034 (
      {stage0_19[426]},
      {stage1_19[240]}
   );
   gpc1_1 gpc2035 (
      {stage0_19[427]},
      {stage1_19[241]}
   );
   gpc1_1 gpc2036 (
      {stage0_19[428]},
      {stage1_19[242]}
   );
   gpc1_1 gpc2037 (
      {stage0_19[429]},
      {stage1_19[243]}
   );
   gpc1_1 gpc2038 (
      {stage0_19[430]},
      {stage1_19[244]}
   );
   gpc1_1 gpc2039 (
      {stage0_19[431]},
      {stage1_19[245]}
   );
   gpc1_1 gpc2040 (
      {stage0_19[432]},
      {stage1_19[246]}
   );
   gpc1_1 gpc2041 (
      {stage0_19[433]},
      {stage1_19[247]}
   );
   gpc1_1 gpc2042 (
      {stage0_19[434]},
      {stage1_19[248]}
   );
   gpc1_1 gpc2043 (
      {stage0_19[435]},
      {stage1_19[249]}
   );
   gpc1_1 gpc2044 (
      {stage0_19[436]},
      {stage1_19[250]}
   );
   gpc1_1 gpc2045 (
      {stage0_19[437]},
      {stage1_19[251]}
   );
   gpc1_1 gpc2046 (
      {stage0_19[438]},
      {stage1_19[252]}
   );
   gpc1_1 gpc2047 (
      {stage0_19[439]},
      {stage1_19[253]}
   );
   gpc1_1 gpc2048 (
      {stage0_19[440]},
      {stage1_19[254]}
   );
   gpc1_1 gpc2049 (
      {stage0_19[441]},
      {stage1_19[255]}
   );
   gpc1_1 gpc2050 (
      {stage0_19[442]},
      {stage1_19[256]}
   );
   gpc1_1 gpc2051 (
      {stage0_19[443]},
      {stage1_19[257]}
   );
   gpc1_1 gpc2052 (
      {stage0_19[444]},
      {stage1_19[258]}
   );
   gpc1_1 gpc2053 (
      {stage0_19[445]},
      {stage1_19[259]}
   );
   gpc1_1 gpc2054 (
      {stage0_19[446]},
      {stage1_19[260]}
   );
   gpc1_1 gpc2055 (
      {stage0_19[447]},
      {stage1_19[261]}
   );
   gpc1_1 gpc2056 (
      {stage0_19[448]},
      {stage1_19[262]}
   );
   gpc1_1 gpc2057 (
      {stage0_19[449]},
      {stage1_19[263]}
   );
   gpc1_1 gpc2058 (
      {stage0_19[450]},
      {stage1_19[264]}
   );
   gpc1_1 gpc2059 (
      {stage0_19[451]},
      {stage1_19[265]}
   );
   gpc1_1 gpc2060 (
      {stage0_19[452]},
      {stage1_19[266]}
   );
   gpc1_1 gpc2061 (
      {stage0_19[453]},
      {stage1_19[267]}
   );
   gpc1_1 gpc2062 (
      {stage0_19[454]},
      {stage1_19[268]}
   );
   gpc1_1 gpc2063 (
      {stage0_19[455]},
      {stage1_19[269]}
   );
   gpc1_1 gpc2064 (
      {stage0_19[456]},
      {stage1_19[270]}
   );
   gpc1_1 gpc2065 (
      {stage0_19[457]},
      {stage1_19[271]}
   );
   gpc1_1 gpc2066 (
      {stage0_19[458]},
      {stage1_19[272]}
   );
   gpc1_1 gpc2067 (
      {stage0_19[459]},
      {stage1_19[273]}
   );
   gpc1_1 gpc2068 (
      {stage0_19[460]},
      {stage1_19[274]}
   );
   gpc1_1 gpc2069 (
      {stage0_19[461]},
      {stage1_19[275]}
   );
   gpc1_1 gpc2070 (
      {stage0_19[462]},
      {stage1_19[276]}
   );
   gpc1_1 gpc2071 (
      {stage0_19[463]},
      {stage1_19[277]}
   );
   gpc1_1 gpc2072 (
      {stage0_19[464]},
      {stage1_19[278]}
   );
   gpc1_1 gpc2073 (
      {stage0_19[465]},
      {stage1_19[279]}
   );
   gpc1_1 gpc2074 (
      {stage0_19[466]},
      {stage1_19[280]}
   );
   gpc1_1 gpc2075 (
      {stage0_19[467]},
      {stage1_19[281]}
   );
   gpc1_1 gpc2076 (
      {stage0_19[468]},
      {stage1_19[282]}
   );
   gpc1_1 gpc2077 (
      {stage0_19[469]},
      {stage1_19[283]}
   );
   gpc1_1 gpc2078 (
      {stage0_19[470]},
      {stage1_19[284]}
   );
   gpc1_1 gpc2079 (
      {stage0_19[471]},
      {stage1_19[285]}
   );
   gpc1_1 gpc2080 (
      {stage0_19[472]},
      {stage1_19[286]}
   );
   gpc1_1 gpc2081 (
      {stage0_19[473]},
      {stage1_19[287]}
   );
   gpc1_1 gpc2082 (
      {stage0_19[474]},
      {stage1_19[288]}
   );
   gpc1_1 gpc2083 (
      {stage0_19[475]},
      {stage1_19[289]}
   );
   gpc1_1 gpc2084 (
      {stage0_19[476]},
      {stage1_19[290]}
   );
   gpc1_1 gpc2085 (
      {stage0_19[477]},
      {stage1_19[291]}
   );
   gpc1_1 gpc2086 (
      {stage0_19[478]},
      {stage1_19[292]}
   );
   gpc1_1 gpc2087 (
      {stage0_19[479]},
      {stage1_19[293]}
   );
   gpc1_1 gpc2088 (
      {stage0_19[480]},
      {stage1_19[294]}
   );
   gpc1_1 gpc2089 (
      {stage0_19[481]},
      {stage1_19[295]}
   );
   gpc1_1 gpc2090 (
      {stage0_19[482]},
      {stage1_19[296]}
   );
   gpc1_1 gpc2091 (
      {stage0_19[483]},
      {stage1_19[297]}
   );
   gpc1_1 gpc2092 (
      {stage0_19[484]},
      {stage1_19[298]}
   );
   gpc1_1 gpc2093 (
      {stage0_19[485]},
      {stage1_19[299]}
   );
   gpc1_1 gpc2094 (
      {stage0_20[478]},
      {stage1_20[181]}
   );
   gpc1_1 gpc2095 (
      {stage0_20[479]},
      {stage1_20[182]}
   );
   gpc1_1 gpc2096 (
      {stage0_20[480]},
      {stage1_20[183]}
   );
   gpc1_1 gpc2097 (
      {stage0_20[481]},
      {stage1_20[184]}
   );
   gpc1_1 gpc2098 (
      {stage0_20[482]},
      {stage1_20[185]}
   );
   gpc1_1 gpc2099 (
      {stage0_20[483]},
      {stage1_20[186]}
   );
   gpc1_1 gpc2100 (
      {stage0_20[484]},
      {stage1_20[187]}
   );
   gpc1_1 gpc2101 (
      {stage0_20[485]},
      {stage1_20[188]}
   );
   gpc1_1 gpc2102 (
      {stage0_22[422]},
      {stage1_22[187]}
   );
   gpc1_1 gpc2103 (
      {stage0_22[423]},
      {stage1_22[188]}
   );
   gpc1_1 gpc2104 (
      {stage0_22[424]},
      {stage1_22[189]}
   );
   gpc1_1 gpc2105 (
      {stage0_22[425]},
      {stage1_22[190]}
   );
   gpc1_1 gpc2106 (
      {stage0_22[426]},
      {stage1_22[191]}
   );
   gpc1_1 gpc2107 (
      {stage0_22[427]},
      {stage1_22[192]}
   );
   gpc1_1 gpc2108 (
      {stage0_22[428]},
      {stage1_22[193]}
   );
   gpc1_1 gpc2109 (
      {stage0_22[429]},
      {stage1_22[194]}
   );
   gpc1_1 gpc2110 (
      {stage0_22[430]},
      {stage1_22[195]}
   );
   gpc1_1 gpc2111 (
      {stage0_22[431]},
      {stage1_22[196]}
   );
   gpc1_1 gpc2112 (
      {stage0_22[432]},
      {stage1_22[197]}
   );
   gpc1_1 gpc2113 (
      {stage0_22[433]},
      {stage1_22[198]}
   );
   gpc1_1 gpc2114 (
      {stage0_22[434]},
      {stage1_22[199]}
   );
   gpc1_1 gpc2115 (
      {stage0_22[435]},
      {stage1_22[200]}
   );
   gpc1_1 gpc2116 (
      {stage0_22[436]},
      {stage1_22[201]}
   );
   gpc1_1 gpc2117 (
      {stage0_22[437]},
      {stage1_22[202]}
   );
   gpc1_1 gpc2118 (
      {stage0_22[438]},
      {stage1_22[203]}
   );
   gpc1_1 gpc2119 (
      {stage0_22[439]},
      {stage1_22[204]}
   );
   gpc1_1 gpc2120 (
      {stage0_22[440]},
      {stage1_22[205]}
   );
   gpc1_1 gpc2121 (
      {stage0_22[441]},
      {stage1_22[206]}
   );
   gpc1_1 gpc2122 (
      {stage0_22[442]},
      {stage1_22[207]}
   );
   gpc1_1 gpc2123 (
      {stage0_22[443]},
      {stage1_22[208]}
   );
   gpc1_1 gpc2124 (
      {stage0_22[444]},
      {stage1_22[209]}
   );
   gpc1_1 gpc2125 (
      {stage0_22[445]},
      {stage1_22[210]}
   );
   gpc1_1 gpc2126 (
      {stage0_22[446]},
      {stage1_22[211]}
   );
   gpc1_1 gpc2127 (
      {stage0_22[447]},
      {stage1_22[212]}
   );
   gpc1_1 gpc2128 (
      {stage0_22[448]},
      {stage1_22[213]}
   );
   gpc1_1 gpc2129 (
      {stage0_22[449]},
      {stage1_22[214]}
   );
   gpc1_1 gpc2130 (
      {stage0_22[450]},
      {stage1_22[215]}
   );
   gpc1_1 gpc2131 (
      {stage0_22[451]},
      {stage1_22[216]}
   );
   gpc1_1 gpc2132 (
      {stage0_22[452]},
      {stage1_22[217]}
   );
   gpc1_1 gpc2133 (
      {stage0_22[453]},
      {stage1_22[218]}
   );
   gpc1_1 gpc2134 (
      {stage0_22[454]},
      {stage1_22[219]}
   );
   gpc1_1 gpc2135 (
      {stage0_22[455]},
      {stage1_22[220]}
   );
   gpc1_1 gpc2136 (
      {stage0_22[456]},
      {stage1_22[221]}
   );
   gpc1_1 gpc2137 (
      {stage0_22[457]},
      {stage1_22[222]}
   );
   gpc1_1 gpc2138 (
      {stage0_22[458]},
      {stage1_22[223]}
   );
   gpc1_1 gpc2139 (
      {stage0_22[459]},
      {stage1_22[224]}
   );
   gpc1_1 gpc2140 (
      {stage0_22[460]},
      {stage1_22[225]}
   );
   gpc1_1 gpc2141 (
      {stage0_22[461]},
      {stage1_22[226]}
   );
   gpc1_1 gpc2142 (
      {stage0_22[462]},
      {stage1_22[227]}
   );
   gpc1_1 gpc2143 (
      {stage0_22[463]},
      {stage1_22[228]}
   );
   gpc1_1 gpc2144 (
      {stage0_22[464]},
      {stage1_22[229]}
   );
   gpc1_1 gpc2145 (
      {stage0_22[465]},
      {stage1_22[230]}
   );
   gpc1_1 gpc2146 (
      {stage0_22[466]},
      {stage1_22[231]}
   );
   gpc1_1 gpc2147 (
      {stage0_22[467]},
      {stage1_22[232]}
   );
   gpc1_1 gpc2148 (
      {stage0_22[468]},
      {stage1_22[233]}
   );
   gpc1_1 gpc2149 (
      {stage0_22[469]},
      {stage1_22[234]}
   );
   gpc1_1 gpc2150 (
      {stage0_22[470]},
      {stage1_22[235]}
   );
   gpc1_1 gpc2151 (
      {stage0_22[471]},
      {stage1_22[236]}
   );
   gpc1_1 gpc2152 (
      {stage0_22[472]},
      {stage1_22[237]}
   );
   gpc1_1 gpc2153 (
      {stage0_22[473]},
      {stage1_22[238]}
   );
   gpc1_1 gpc2154 (
      {stage0_22[474]},
      {stage1_22[239]}
   );
   gpc1_1 gpc2155 (
      {stage0_22[475]},
      {stage1_22[240]}
   );
   gpc1_1 gpc2156 (
      {stage0_22[476]},
      {stage1_22[241]}
   );
   gpc1_1 gpc2157 (
      {stage0_22[477]},
      {stage1_22[242]}
   );
   gpc1_1 gpc2158 (
      {stage0_22[478]},
      {stage1_22[243]}
   );
   gpc1_1 gpc2159 (
      {stage0_22[479]},
      {stage1_22[244]}
   );
   gpc1_1 gpc2160 (
      {stage0_22[480]},
      {stage1_22[245]}
   );
   gpc1_1 gpc2161 (
      {stage0_22[481]},
      {stage1_22[246]}
   );
   gpc1_1 gpc2162 (
      {stage0_22[482]},
      {stage1_22[247]}
   );
   gpc1_1 gpc2163 (
      {stage0_22[483]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2164 (
      {stage0_22[484]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2165 (
      {stage0_22[485]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2166 (
      {stage0_23[474]},
      {stage1_23[166]}
   );
   gpc1_1 gpc2167 (
      {stage0_23[475]},
      {stage1_23[167]}
   );
   gpc1_1 gpc2168 (
      {stage0_23[476]},
      {stage1_23[168]}
   );
   gpc1_1 gpc2169 (
      {stage0_23[477]},
      {stage1_23[169]}
   );
   gpc1_1 gpc2170 (
      {stage0_23[478]},
      {stage1_23[170]}
   );
   gpc1_1 gpc2171 (
      {stage0_23[479]},
      {stage1_23[171]}
   );
   gpc1_1 gpc2172 (
      {stage0_23[480]},
      {stage1_23[172]}
   );
   gpc1_1 gpc2173 (
      {stage0_23[481]},
      {stage1_23[173]}
   );
   gpc1_1 gpc2174 (
      {stage0_23[482]},
      {stage1_23[174]}
   );
   gpc1_1 gpc2175 (
      {stage0_23[483]},
      {stage1_23[175]}
   );
   gpc1_1 gpc2176 (
      {stage0_23[484]},
      {stage1_23[176]}
   );
   gpc1_1 gpc2177 (
      {stage0_23[485]},
      {stage1_23[177]}
   );
   gpc1_1 gpc2178 (
      {stage0_26[445]},
      {stage1_26[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_26[446]},
      {stage1_26[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_26[447]},
      {stage1_26[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_26[448]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_26[449]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_26[450]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_26[451]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_26[452]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_26[453]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_26[454]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_26[455]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_26[456]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_26[457]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_26[458]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_26[459]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_26[460]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_26[461]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_26[462]},
      {stage1_26[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_26[463]},
      {stage1_26[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_26[464]},
      {stage1_26[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_26[465]},
      {stage1_26[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_26[466]},
      {stage1_26[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_26[467]},
      {stage1_26[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_26[468]},
      {stage1_26[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_26[469]},
      {stage1_26[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_26[470]},
      {stage1_26[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_26[471]},
      {stage1_26[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_26[472]},
      {stage1_26[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_26[473]},
      {stage1_26[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_26[474]},
      {stage1_26[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_26[475]},
      {stage1_26[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_26[476]},
      {stage1_26[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_26[477]},
      {stage1_26[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_26[478]},
      {stage1_26[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_26[479]},
      {stage1_26[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_26[480]},
      {stage1_26[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_26[481]},
      {stage1_26[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_26[482]},
      {stage1_26[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_26[483]},
      {stage1_26[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_26[484]},
      {stage1_26[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_26[485]},
      {stage1_26[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_27[483]},
      {stage1_27[156]}
   );
   gpc1_1 gpc2220 (
      {stage0_27[484]},
      {stage1_27[157]}
   );
   gpc1_1 gpc2221 (
      {stage0_27[485]},
      {stage1_27[158]}
   );
   gpc1_1 gpc2222 (
      {stage0_28[450]},
      {stage1_28[216]}
   );
   gpc1_1 gpc2223 (
      {stage0_28[451]},
      {stage1_28[217]}
   );
   gpc1_1 gpc2224 (
      {stage0_28[452]},
      {stage1_28[218]}
   );
   gpc1_1 gpc2225 (
      {stage0_28[453]},
      {stage1_28[219]}
   );
   gpc1_1 gpc2226 (
      {stage0_28[454]},
      {stage1_28[220]}
   );
   gpc1_1 gpc2227 (
      {stage0_28[455]},
      {stage1_28[221]}
   );
   gpc1_1 gpc2228 (
      {stage0_28[456]},
      {stage1_28[222]}
   );
   gpc1_1 gpc2229 (
      {stage0_28[457]},
      {stage1_28[223]}
   );
   gpc1_1 gpc2230 (
      {stage0_28[458]},
      {stage1_28[224]}
   );
   gpc1_1 gpc2231 (
      {stage0_28[459]},
      {stage1_28[225]}
   );
   gpc1_1 gpc2232 (
      {stage0_28[460]},
      {stage1_28[226]}
   );
   gpc1_1 gpc2233 (
      {stage0_28[461]},
      {stage1_28[227]}
   );
   gpc1_1 gpc2234 (
      {stage0_28[462]},
      {stage1_28[228]}
   );
   gpc1_1 gpc2235 (
      {stage0_28[463]},
      {stage1_28[229]}
   );
   gpc1_1 gpc2236 (
      {stage0_28[464]},
      {stage1_28[230]}
   );
   gpc1_1 gpc2237 (
      {stage0_28[465]},
      {stage1_28[231]}
   );
   gpc1_1 gpc2238 (
      {stage0_28[466]},
      {stage1_28[232]}
   );
   gpc1_1 gpc2239 (
      {stage0_28[467]},
      {stage1_28[233]}
   );
   gpc1_1 gpc2240 (
      {stage0_28[468]},
      {stage1_28[234]}
   );
   gpc1_1 gpc2241 (
      {stage0_28[469]},
      {stage1_28[235]}
   );
   gpc1_1 gpc2242 (
      {stage0_28[470]},
      {stage1_28[236]}
   );
   gpc1_1 gpc2243 (
      {stage0_28[471]},
      {stage1_28[237]}
   );
   gpc1_1 gpc2244 (
      {stage0_28[472]},
      {stage1_28[238]}
   );
   gpc1_1 gpc2245 (
      {stage0_28[473]},
      {stage1_28[239]}
   );
   gpc1_1 gpc2246 (
      {stage0_28[474]},
      {stage1_28[240]}
   );
   gpc1_1 gpc2247 (
      {stage0_28[475]},
      {stage1_28[241]}
   );
   gpc1_1 gpc2248 (
      {stage0_28[476]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2249 (
      {stage0_28[477]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2250 (
      {stage0_28[478]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2251 (
      {stage0_28[479]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2252 (
      {stage0_28[480]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2253 (
      {stage0_28[481]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2254 (
      {stage0_28[482]},
      {stage1_28[248]}
   );
   gpc1_1 gpc2255 (
      {stage0_28[483]},
      {stage1_28[249]}
   );
   gpc1_1 gpc2256 (
      {stage0_28[484]},
      {stage1_28[250]}
   );
   gpc1_1 gpc2257 (
      {stage0_28[485]},
      {stage1_28[251]}
   );
   gpc1_1 gpc2258 (
      {stage0_30[480]},
      {stage1_30[166]}
   );
   gpc1_1 gpc2259 (
      {stage0_30[481]},
      {stage1_30[167]}
   );
   gpc1_1 gpc2260 (
      {stage0_30[482]},
      {stage1_30[168]}
   );
   gpc1_1 gpc2261 (
      {stage0_30[483]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2262 (
      {stage0_30[484]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2263 (
      {stage0_30[485]},
      {stage1_30[171]}
   );
   gpc1163_5 gpc2264 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc2265 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc2266 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2267 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2268 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc2269 (
      {stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc2270 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2271 (
      {stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc2272 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc2273 (
      {stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc2274 (
      {stage1_0[57], stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc2275 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67], stage1_0[68]},
      {stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2276 (
      {stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72], stage1_0[73], stage1_0[74]},
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc2277 (
      {stage1_0[75], stage1_0[76], stage1_0[77], stage1_0[78], stage1_0[79], stage1_0[80]},
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc2278 (
      {stage1_0[81], stage1_0[82], stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86]},
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83], stage1_2[84]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc2279 (
      {stage1_0[87], stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc2280 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97], stage1_0[98]},
      {stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc2281 (
      {stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102], stage1_0[103], stage1_0[104]},
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc2282 (
      {stage1_0[105], stage1_0[106], stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110]},
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107], stage1_2[108]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc2283 (
      {stage1_0[111], stage1_0[112], stage1_0[113], stage1_0[114], stage1_0[115], stage1_0[116]},
      {stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113], stage1_2[114]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc2284 (
      {stage1_0[117], stage1_0[118], stage1_0[119], stage1_0[120], stage1_0[121]},
      {stage1_1[6]},
      {stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc615_5 gpc2285 (
      {stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125], stage1_0[126]},
      {stage1_1[7]},
      {stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc2286 (
      {stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2287 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage2_5[1],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2288 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18]},
      {stage2_5[2],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2289 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage2_5[3],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2290 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30]},
      {stage2_5[4],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2291 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage2_5[5],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2292 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage2_5[6],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2293 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage2_5[7],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2294 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54]},
      {stage2_5[8],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2295 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[9],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc606_5 gpc2296 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137], stage1_2[138]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[10],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc606_5 gpc2297 (
      {stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143], stage1_2[144]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[11],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc606_5 gpc2298 (
      {stage1_2[145], stage1_2[146], stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[12],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc606_5 gpc2299 (
      {stage1_2[151], stage1_2[152], stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[13],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc606_5 gpc2300 (
      {stage1_2[157], stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[14],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc606_5 gpc2301 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167], stage1_2[168]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[15],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc606_5 gpc2302 (
      {stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172], stage1_2[173], stage1_2[174]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[16],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc606_5 gpc2303 (
      {stage1_2[175], stage1_2[176], stage1_2[177], stage1_2[178], stage1_2[179], stage1_2[180]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[17],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc2304 (
      {stage1_2[181], stage1_2[182], stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[18],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc2305 (
      {stage1_2[187], stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[19],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc2306 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197], stage1_2[198]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[20],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc2307 (
      {stage1_2[199], stage1_2[200], stage1_2[201], stage1_2[202], stage1_2[203], stage1_2[204]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[21],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2308 (
      {stage1_2[205], stage1_2[206], stage1_2[207], stage1_2[208], stage1_2[209]},
      {stage1_3[55]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[22],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2309 (
      {stage1_2[210], stage1_2[211], stage1_2[212], stage1_2[213], stage1_2[214]},
      {stage1_3[56]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[23],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2310 (
      {stage1_2[215], stage1_2[216], stage1_2[217], stage1_2[218], stage1_2[219]},
      {stage1_3[57]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[24],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2311 (
      {stage1_2[220], stage1_2[221], stage1_2[222], stage1_2[223], stage1_2[224]},
      {stage1_3[58]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[25],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc2312 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[17],stage2_5[26],stage2_4[48],stage2_3[48]}
   );
   gpc606_5 gpc2313 (
      {stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[18],stage2_5[27],stage2_4[49],stage2_3[49]}
   );
   gpc606_5 gpc2314 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[19],stage2_5[28],stage2_4[50],stage2_3[50]}
   );
   gpc606_5 gpc2315 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[20],stage2_5[29],stage2_4[51],stage2_3[51]}
   );
   gpc606_5 gpc2316 (
      {stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[21],stage2_5[30],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93]},
      {stage1_4[102]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[22],stage2_5[31],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97], stage1_3[98]},
      {stage1_4[103]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[23],stage2_5[32],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage1_4[104]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[24],stage2_5[33],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108]},
      {stage1_4[105]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[25],stage2_5[34],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage1_4[106]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[26],stage2_5[35],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118]},
      {stage1_4[107]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[27],stage2_5[36],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123]},
      {stage1_4[108]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[28],stage2_5[37],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2324 (
      {stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127], stage1_3[128]},
      {stage1_4[109]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[29],stage2_5[38],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2325 (
      {stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage1_4[110]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[30],stage2_5[39],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2326 (
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[111]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[31],stage2_5[40],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2327 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[112]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[32],stage2_5[41],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2328 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[113]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[33],stage2_5[42],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2329 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[114]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[34],stage2_5[43],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2330 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[115]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[35],stage2_5[44],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2331 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[116]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[36],stage2_5[45],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2332 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[117]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[37],stage2_5[46],stage2_4[68],stage2_3[68]}
   );
   gpc1163_5 gpc2333 (
      {stage1_4[118], stage1_4[119], stage1_4[120]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[21],stage2_6[38],stage2_5[47],stage2_4[69]}
   );
   gpc615_5 gpc2334 (
      {stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage1_5[132]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[22],stage2_6[39],stage2_5[48],stage2_4[70]}
   );
   gpc615_5 gpc2335 (
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130]},
      {stage1_5[133]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[23],stage2_6[40],stage2_5[49],stage2_4[71]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_5[134]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[24],stage2_6[41],stage2_5[50],stage2_4[72]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[135]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[25],stage2_6[42],stage2_5[51],stage2_4[73]}
   );
   gpc615_5 gpc2338 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145]},
      {stage1_5[136]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[26],stage2_6[43],stage2_5[52],stage2_4[74]}
   );
   gpc615_5 gpc2339 (
      {stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_5[137]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[27],stage2_6[44],stage2_5[53],stage2_4[75]}
   );
   gpc615_5 gpc2340 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage1_5[138]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[28],stage2_6[45],stage2_5[54],stage2_4[76]}
   );
   gpc615_5 gpc2341 (
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160]},
      {stage1_5[139]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[29],stage2_6[46],stage2_5[55],stage2_4[77]}
   );
   gpc615_5 gpc2342 (
      {stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_5[140]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[30],stage2_6[47],stage2_5[56],stage2_4[78]}
   );
   gpc615_5 gpc2343 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_5[141]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[31],stage2_6[48],stage2_5[57],stage2_4[79]}
   );
   gpc615_5 gpc2344 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175]},
      {stage1_5[142]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[32],stage2_6[49],stage2_5[58],stage2_4[80]}
   );
   gpc615_5 gpc2345 (
      {stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_5[143]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[33],stage2_6[50],stage2_5[59],stage2_4[81]}
   );
   gpc615_5 gpc2346 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage1_5[144]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[34],stage2_6[51],stage2_5[60],stage2_4[82]}
   );
   gpc615_5 gpc2347 (
      {stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190]},
      {stage1_5[145]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[35],stage2_6[52],stage2_5[61],stage2_4[83]}
   );
   gpc615_5 gpc2348 (
      {stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_5[146]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[36],stage2_6[53],stage2_5[62],stage2_4[84]}
   );
   gpc615_5 gpc2349 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_5[147]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[37],stage2_6[54],stage2_5[63],stage2_4[85]}
   );
   gpc615_5 gpc2350 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205]},
      {stage1_5[148]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[38],stage2_6[55],stage2_5[64],stage2_4[86]}
   );
   gpc615_5 gpc2351 (
      {stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_5[149]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[39],stage2_6[56],stage2_5[65],stage2_4[87]}
   );
   gpc615_5 gpc2352 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215]},
      {stage1_5[150]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[40],stage2_6[57],stage2_5[66],stage2_4[88]}
   );
   gpc615_5 gpc2353 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220]},
      {stage1_5[151]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[41],stage2_6[58],stage2_5[67],stage2_4[89]}
   );
   gpc615_5 gpc2354 (
      {stage1_4[221], stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225]},
      {stage1_5[152]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[42],stage2_6[59],stage2_5[68],stage2_4[90]}
   );
   gpc606_5 gpc2355 (
      {stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157], stage1_5[158]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[22],stage2_7[43],stage2_6[60],stage2_5[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163], stage1_5[164]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[23],stage2_7[44],stage2_6[61],stage2_5[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169], stage1_5[170]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[24],stage2_7[45],stage2_6[62],stage2_5[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175], stage1_5[176]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[25],stage2_7[46],stage2_6[63],stage2_5[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181], stage1_5[182]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[26],stage2_7[47],stage2_6[64],stage2_5[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187], stage1_5[188]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[27],stage2_7[48],stage2_6[65],stage2_5[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193], stage1_5[194]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[28],stage2_7[49],stage2_6[66],stage2_5[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199], stage1_5[200]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[29],stage2_7[50],stage2_6[67],stage2_5[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205], stage1_5[206]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[30],stage2_7[51],stage2_6[68],stage2_5[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_5[207], stage1_5[208], stage1_5[209], stage1_5[210], stage1_5[211], stage1_5[212]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[31],stage2_7[52],stage2_6[69],stage2_5[78]}
   );
   gpc615_5 gpc2365 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_7[61]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[10],stage2_8[32],stage2_7[53],stage2_6[70]}
   );
   gpc615_5 gpc2366 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136]},
      {stage1_7[62]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[11],stage2_8[33],stage2_7[54],stage2_6[71]}
   );
   gpc615_5 gpc2367 (
      {stage1_6[137], stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141]},
      {stage1_7[63]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[12],stage2_8[34],stage2_7[55],stage2_6[72]}
   );
   gpc615_5 gpc2368 (
      {stage1_6[142], stage1_6[143], stage1_6[144], stage1_6[145], stage1_6[146]},
      {stage1_7[64]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[13],stage2_8[35],stage2_7[56],stage2_6[73]}
   );
   gpc615_5 gpc2369 (
      {stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150], stage1_6[151]},
      {stage1_7[65]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[14],stage2_8[36],stage2_7[57],stage2_6[74]}
   );
   gpc615_5 gpc2370 (
      {stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_7[66]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[15],stage2_8[37],stage2_7[58],stage2_6[75]}
   );
   gpc615_5 gpc2371 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_7[67]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[16],stage2_8[38],stage2_7[59],stage2_6[76]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166]},
      {stage1_7[68]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[17],stage2_8[39],stage2_7[60],stage2_6[77]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[167], stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171]},
      {stage1_7[69]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[18],stage2_8[40],stage2_7[61],stage2_6[78]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[172], stage1_6[173], stage1_6[174], stage1_6[175], stage1_6[176]},
      {stage1_7[70]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[19],stage2_8[41],stage2_7[62],stage2_6[79]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180], stage1_6[181]},
      {stage1_7[71]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[20],stage2_8[42],stage2_7[63],stage2_6[80]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_7[72]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[21],stage2_8[43],stage2_7[64],stage2_6[81]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_7[73]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[22],stage2_8[44],stage2_7[65],stage2_6[82]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[74]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[23],stage2_8[45],stage2_7[66],stage2_6[83]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[197], stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201]},
      {stage1_7[75]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[24],stage2_8[46],stage2_7[67],stage2_6[84]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[202], stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206]},
      {stage1_7[76]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[25],stage2_8[47],stage2_7[68],stage2_6[85]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[207], stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211]},
      {stage1_7[77]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[26],stage2_8[48],stage2_7[69],stage2_6[86]}
   );
   gpc615_5 gpc2382 (
      {stage1_6[212], stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216]},
      {stage1_7[78]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[27],stage2_8[49],stage2_7[70],stage2_6[87]}
   );
   gpc615_5 gpc2383 (
      {stage1_6[217], stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221]},
      {stage1_7[79]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[28],stage2_8[50],stage2_7[71],stage2_6[88]}
   );
   gpc615_5 gpc2384 (
      {stage1_6[222], stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226]},
      {stage1_7[80]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[29],stage2_8[51],stage2_7[72],stage2_6[89]}
   );
   gpc615_5 gpc2385 (
      {stage1_6[227], stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231]},
      {stage1_7[81]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[30],stage2_8[52],stage2_7[73],stage2_6[90]}
   );
   gpc615_5 gpc2386 (
      {stage1_6[232], stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236]},
      {stage1_7[82]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[31],stage2_8[53],stage2_7[74],stage2_6[91]}
   );
   gpc615_5 gpc2387 (
      {stage1_6[237], stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241]},
      {stage1_7[83]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[32],stage2_8[54],stage2_7[75],stage2_6[92]}
   );
   gpc615_5 gpc2388 (
      {stage1_6[242], stage1_6[243], stage1_6[244], stage1_6[245], stage1_6[246]},
      {stage1_7[84]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[33],stage2_8[55],stage2_7[76],stage2_6[93]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage1_8[144]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[24],stage2_9[34],stage2_8[56],stage2_7[77]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94]},
      {stage1_8[145]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[25],stage2_9[35],stage2_8[57],stage2_7[78]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[95], stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99]},
      {stage1_8[146]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[26],stage2_9[36],stage2_8[58],stage2_7[79]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104]},
      {stage1_8[147]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[27],stage2_9[37],stage2_8[59],stage2_7[80]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage1_8[148]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[28],stage2_9[38],stage2_8[60],stage2_7[81]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_8[149]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[29],stage2_9[39],stage2_8[61],stage2_7[82]}
   );
   gpc615_5 gpc2395 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage1_8[150]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[30],stage2_9[40],stage2_8[62],stage2_7[83]}
   );
   gpc615_5 gpc2396 (
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124]},
      {stage1_8[151]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[31],stage2_9[41],stage2_8[63],stage2_7[84]}
   );
   gpc615_5 gpc2397 (
      {stage1_7[125], stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129]},
      {stage1_8[152]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[32],stage2_9[42],stage2_8[64],stage2_7[85]}
   );
   gpc615_5 gpc2398 (
      {stage1_7[130], stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134]},
      {stage1_8[153]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[33],stage2_9[43],stage2_8[65],stage2_7[86]}
   );
   gpc615_5 gpc2399 (
      {stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139]},
      {stage1_8[154]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[34],stage2_9[44],stage2_8[66],stage2_7[87]}
   );
   gpc615_5 gpc2400 (
      {stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_8[155]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[35],stage2_9[45],stage2_8[67],stage2_7[88]}
   );
   gpc615_5 gpc2401 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149]},
      {stage1_8[156]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[36],stage2_9[46],stage2_8[68],stage2_7[89]}
   );
   gpc615_5 gpc2402 (
      {stage1_7[150], stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154]},
      {stage1_8[157]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[37],stage2_9[47],stage2_8[69],stage2_7[90]}
   );
   gpc615_5 gpc2403 (
      {stage1_7[155], stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159]},
      {stage1_8[158]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[38],stage2_9[48],stage2_8[70],stage2_7[91]}
   );
   gpc615_5 gpc2404 (
      {stage1_7[160], stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164]},
      {stage1_8[159]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[39],stage2_9[49],stage2_8[71],stage2_7[92]}
   );
   gpc615_5 gpc2405 (
      {stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169]},
      {stage1_8[160]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[40],stage2_9[50],stage2_8[72],stage2_7[93]}
   );
   gpc615_5 gpc2406 (
      {stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_8[161]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[41],stage2_9[51],stage2_8[73],stage2_7[94]}
   );
   gpc615_5 gpc2407 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179]},
      {stage1_8[162]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[42],stage2_9[52],stage2_8[74],stage2_7[95]}
   );
   gpc615_5 gpc2408 (
      {stage1_7[180], stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184]},
      {stage1_8[163]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[43],stage2_9[53],stage2_8[75],stage2_7[96]}
   );
   gpc615_5 gpc2409 (
      {stage1_7[185], stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189]},
      {stage1_8[164]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[44],stage2_9[54],stage2_8[76],stage2_7[97]}
   );
   gpc615_5 gpc2410 (
      {stage1_7[190], stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194]},
      {stage1_8[165]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[45],stage2_9[55],stage2_8[77],stage2_7[98]}
   );
   gpc615_5 gpc2411 (
      {stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199]},
      {stage1_8[166]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[46],stage2_9[56],stage2_8[78],stage2_7[99]}
   );
   gpc615_5 gpc2412 (
      {stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_8[167]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[47],stage2_9[57],stage2_8[79],stage2_7[100]}
   );
   gpc615_5 gpc2413 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209]},
      {stage1_8[168]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[48],stage2_9[58],stage2_8[80],stage2_7[101]}
   );
   gpc615_5 gpc2414 (
      {stage1_7[210], stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214]},
      {stage1_8[169]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[49],stage2_9[59],stage2_8[81],stage2_7[102]}
   );
   gpc623_5 gpc2415 (
      {stage1_7[215], stage1_7[216], stage1_7[217]},
      {stage1_8[170], stage1_8[171]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[50],stage2_9[60],stage2_8[82],stage2_7[103]}
   );
   gpc1415_5 gpc2416 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176]},
      {stage1_9[162]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[27],stage2_10[51],stage2_9[61],stage2_8[83]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[177], stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9]},
      {stage2_12[1],stage2_11[28],stage2_10[52],stage2_9[62],stage2_8[84]}
   );
   gpc606_5 gpc2418 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[29],stage2_10[53],stage2_9[63]}
   );
   gpc606_5 gpc2419 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[30],stage2_10[54],stage2_9[64]}
   );
   gpc606_5 gpc2420 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[31],stage2_10[55],stage2_9[65]}
   );
   gpc615_5 gpc2421 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_10[10]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[3],stage2_12[5],stage2_11[32],stage2_10[56],stage2_9[66]}
   );
   gpc615_5 gpc2422 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190]},
      {stage1_10[11]},
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage2_13[4],stage2_12[6],stage2_11[33],stage2_10[57],stage2_9[67]}
   );
   gpc615_5 gpc2423 (
      {stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_10[12]},
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage2_13[5],stage2_12[7],stage2_11[34],stage2_10[58],stage2_9[68]}
   );
   gpc615_5 gpc2424 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200]},
      {stage1_10[13]},
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage2_13[6],stage2_12[8],stage2_11[35],stage2_10[59],stage2_9[69]}
   );
   gpc615_5 gpc2425 (
      {stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205]},
      {stage1_10[14]},
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage2_13[7],stage2_12[9],stage2_11[36],stage2_10[60],stage2_9[70]}
   );
   gpc615_5 gpc2426 (
      {stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_10[15]},
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage2_13[8],stage2_12[10],stage2_11[37],stage2_10[61],stage2_9[71]}
   );
   gpc117_4 gpc2427 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[55]},
      {stage1_12[0]},
      {stage2_13[9],stage2_12[11],stage2_11[38],stage2_10[62]}
   );
   gpc117_4 gpc2428 (
      {stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_11[56]},
      {stage1_12[1]},
      {stage2_13[10],stage2_12[12],stage2_11[39],stage2_10[63]}
   );
   gpc117_4 gpc2429 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[57]},
      {stage1_12[2]},
      {stage2_13[11],stage2_12[13],stage2_11[40],stage2_10[64]}
   );
   gpc117_4 gpc2430 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage1_11[58]},
      {stage1_12[3]},
      {stage2_13[12],stage2_12[14],stage2_11[41],stage2_10[65]}
   );
   gpc117_4 gpc2431 (
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[59]},
      {stage1_12[4]},
      {stage2_13[13],stage2_12[15],stage2_11[42],stage2_10[66]}
   );
   gpc117_4 gpc2432 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57]},
      {stage1_11[60]},
      {stage1_12[5]},
      {stage2_13[14],stage2_12[16],stage2_11[43],stage2_10[67]}
   );
   gpc117_4 gpc2433 (
      {stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64]},
      {stage1_11[61]},
      {stage1_12[6]},
      {stage2_13[15],stage2_12[17],stage2_11[44],stage2_10[68]}
   );
   gpc117_4 gpc2434 (
      {stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_11[62]},
      {stage1_12[7]},
      {stage2_13[16],stage2_12[18],stage2_11[45],stage2_10[69]}
   );
   gpc117_4 gpc2435 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[63]},
      {stage1_12[8]},
      {stage2_13[17],stage2_12[19],stage2_11[46],stage2_10[70]}
   );
   gpc117_4 gpc2436 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage1_11[64]},
      {stage1_12[9]},
      {stage2_13[18],stage2_12[20],stage2_11[47],stage2_10[71]}
   );
   gpc117_4 gpc2437 (
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92]},
      {stage1_11[65]},
      {stage1_12[10]},
      {stage2_13[19],stage2_12[21],stage2_11[48],stage2_10[72]}
   );
   gpc117_4 gpc2438 (
      {stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99]},
      {stage1_11[66]},
      {stage1_12[11]},
      {stage2_13[20],stage2_12[22],stage2_11[49],stage2_10[73]}
   );
   gpc117_4 gpc2439 (
      {stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[67]},
      {stage1_12[12]},
      {stage2_13[21],stage2_12[23],stage2_11[50],stage2_10[74]}
   );
   gpc117_4 gpc2440 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_11[68]},
      {stage1_12[13]},
      {stage2_13[22],stage2_12[24],stage2_11[51],stage2_10[75]}
   );
   gpc117_4 gpc2441 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120]},
      {stage1_11[69]},
      {stage1_12[14]},
      {stage2_13[23],stage2_12[25],stage2_11[52],stage2_10[76]}
   );
   gpc117_4 gpc2442 (
      {stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125], stage1_10[126], stage1_10[127]},
      {stage1_11[70]},
      {stage1_12[15]},
      {stage2_13[24],stage2_12[26],stage2_11[53],stage2_10[77]}
   );
   gpc117_4 gpc2443 (
      {stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[71]},
      {stage1_12[16]},
      {stage2_13[25],stage2_12[27],stage2_11[54],stage2_10[78]}
   );
   gpc117_4 gpc2444 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141]},
      {stage1_11[72]},
      {stage1_12[17]},
      {stage2_13[26],stage2_12[28],stage2_11[55],stage2_10[79]}
   );
   gpc117_4 gpc2445 (
      {stage1_10[142], stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_11[73]},
      {stage1_12[18]},
      {stage2_13[27],stage2_12[29],stage2_11[56],stage2_10[80]}
   );
   gpc117_4 gpc2446 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_11[74]},
      {stage1_12[19]},
      {stage2_13[28],stage2_12[30],stage2_11[57],stage2_10[81]}
   );
   gpc606_5 gpc2447 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[0],stage2_13[29],stage2_12[31],stage2_11[58],stage2_10[82]}
   );
   gpc606_5 gpc2448 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[1],stage2_13[30],stage2_12[32],stage2_11[59],stage2_10[83]}
   );
   gpc606_5 gpc2449 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37]},
      {stage2_14[2],stage2_13[31],stage2_12[33],stage2_11[60],stage2_10[84]}
   );
   gpc606_5 gpc2450 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43]},
      {stage2_14[3],stage2_13[32],stage2_12[34],stage2_11[61],stage2_10[85]}
   );
   gpc606_5 gpc2451 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage2_14[4],stage2_13[33],stage2_12[35],stage2_11[62],stage2_10[86]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78], stage1_11[79]},
      {stage1_12[50]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[34],stage2_12[36],stage2_11[63]}
   );
   gpc615_5 gpc2453 (
      {stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_12[51]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[35],stage2_12[37],stage2_11[64]}
   );
   gpc615_5 gpc2454 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage1_12[52]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[36],stage2_12[38],stage2_11[65]}
   );
   gpc615_5 gpc2455 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[53]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[8],stage2_13[37],stage2_12[39],stage2_11[66]}
   );
   gpc615_5 gpc2456 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[54]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[9],stage2_13[38],stage2_12[40],stage2_11[67]}
   );
   gpc615_5 gpc2457 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[55]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[10],stage2_13[39],stage2_12[41],stage2_11[68]}
   );
   gpc615_5 gpc2458 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[56]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[11],stage2_13[40],stage2_12[42],stage2_11[69]}
   );
   gpc615_5 gpc2459 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[57]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[12],stage2_13[41],stage2_12[43],stage2_11[70]}
   );
   gpc615_5 gpc2460 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[58]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[13],stage2_13[42],stage2_12[44],stage2_11[71]}
   );
   gpc615_5 gpc2461 (
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124]},
      {stage1_12[59]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[14],stage2_13[43],stage2_12[45],stage2_11[72]}
   );
   gpc615_5 gpc2462 (
      {stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[60]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[15],stage2_13[44],stage2_12[46],stage2_11[73]}
   );
   gpc615_5 gpc2463 (
      {stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133], stage1_11[134]},
      {stage1_12[61]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[16],stage2_13[45],stage2_12[47],stage2_11[74]}
   );
   gpc615_5 gpc2464 (
      {stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139]},
      {stage1_12[62]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[17],stage2_13[46],stage2_12[48],stage2_11[75]}
   );
   gpc615_5 gpc2465 (
      {stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[63]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[18],stage2_13[47],stage2_12[49],stage2_11[76]}
   );
   gpc615_5 gpc2466 (
      {stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149]},
      {stage1_12[64]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[19],stage2_13[48],stage2_12[50],stage2_11[77]}
   );
   gpc615_5 gpc2467 (
      {stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154]},
      {stage1_12[65]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[20],stage2_13[49],stage2_12[51],stage2_11[78]}
   );
   gpc615_5 gpc2468 (
      {stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[66]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[21],stage2_13[50],stage2_12[52],stage2_11[79]}
   );
   gpc615_5 gpc2469 (
      {stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163], stage1_11[164]},
      {stage1_12[67]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[22],stage2_13[51],stage2_12[53],stage2_11[80]}
   );
   gpc615_5 gpc2470 (
      {stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168], stage1_11[169]},
      {stage1_12[68]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[23],stage2_13[52],stage2_12[54],stage2_11[81]}
   );
   gpc615_5 gpc2471 (
      {stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173], stage1_11[174]},
      {stage1_12[69]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[24],stage2_13[53],stage2_12[55],stage2_11[82]}
   );
   gpc615_5 gpc2472 (
      {stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178], stage1_11[179]},
      {stage1_12[70]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[25],stage2_13[54],stage2_12[56],stage2_11[83]}
   );
   gpc615_5 gpc2473 (
      {stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183], stage1_11[184]},
      {stage1_12[71]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[26],stage2_13[55],stage2_12[57],stage2_11[84]}
   );
   gpc615_5 gpc2474 (
      {stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188], stage1_11[189]},
      {stage1_12[72]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[27],stage2_13[56],stage2_12[58],stage2_11[85]}
   );
   gpc615_5 gpc2475 (
      {stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193], stage1_11[194]},
      {stage1_12[73]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[28],stage2_13[57],stage2_12[59],stage2_11[86]}
   );
   gpc615_5 gpc2476 (
      {stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198], stage1_11[199]},
      {stage1_12[74]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[29],stage2_13[58],stage2_12[60],stage2_11[87]}
   );
   gpc615_5 gpc2477 (
      {stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203], stage1_11[204]},
      {stage1_12[75]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[30],stage2_13[59],stage2_12[61],stage2_11[88]}
   );
   gpc615_5 gpc2478 (
      {stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208], stage1_11[209]},
      {stage1_12[76]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[31],stage2_13[60],stage2_12[62],stage2_11[89]}
   );
   gpc615_5 gpc2479 (
      {stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213], stage1_11[214]},
      {stage1_12[77]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[32],stage2_13[61],stage2_12[63],stage2_11[90]}
   );
   gpc615_5 gpc2480 (
      {stage1_11[215], stage1_11[216], stage1_11[217], stage1_11[218], stage1_11[219]},
      {stage1_12[78]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[33],stage2_13[62],stage2_12[64],stage2_11[91]}
   );
   gpc606_5 gpc2481 (
      {stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[29],stage2_14[34],stage2_13[63],stage2_12[65]}
   );
   gpc606_5 gpc2482 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89], stage1_12[90]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[30],stage2_14[35],stage2_13[64],stage2_12[66]}
   );
   gpc606_5 gpc2483 (
      {stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95], stage1_12[96]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[31],stage2_14[36],stage2_13[65],stage2_12[67]}
   );
   gpc606_5 gpc2484 (
      {stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[32],stage2_14[37],stage2_13[66],stage2_12[68]}
   );
   gpc606_5 gpc2485 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[33],stage2_14[38],stage2_13[67],stage2_12[69]}
   );
   gpc606_5 gpc2486 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[34],stage2_14[39],stage2_13[68],stage2_12[70]}
   );
   gpc606_5 gpc2487 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[35],stage2_14[40],stage2_13[69],stage2_12[71]}
   );
   gpc606_5 gpc2488 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[36],stage2_14[41],stage2_13[70],stage2_12[72]}
   );
   gpc606_5 gpc2489 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[37],stage2_14[42],stage2_13[71],stage2_12[73]}
   );
   gpc606_5 gpc2490 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[38],stage2_14[43],stage2_13[72],stage2_12[74]}
   );
   gpc606_5 gpc2491 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[39],stage2_14[44],stage2_13[73],stage2_12[75]}
   );
   gpc606_5 gpc2492 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[40],stage2_14[45],stage2_13[74],stage2_12[76]}
   );
   gpc606_5 gpc2493 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[41],stage2_14[46],stage2_13[75],stage2_12[77]}
   );
   gpc606_5 gpc2494 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[42],stage2_14[47],stage2_13[76],stage2_12[78]}
   );
   gpc606_5 gpc2495 (
      {stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[43],stage2_14[48],stage2_13[77],stage2_12[79]}
   );
   gpc606_5 gpc2496 (
      {stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[44],stage2_14[49],stage2_13[78],stage2_12[80]}
   );
   gpc606_5 gpc2497 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[45],stage2_14[50],stage2_13[79],stage2_12[81]}
   );
   gpc606_5 gpc2498 (
      {stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[46],stage2_14[51],stage2_13[80],stage2_12[82]}
   );
   gpc606_5 gpc2499 (
      {stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[47],stage2_14[52],stage2_13[81],stage2_12[83]}
   );
   gpc606_5 gpc2500 (
      {stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[48],stage2_14[53],stage2_13[82],stage2_12[84]}
   );
   gpc606_5 gpc2501 (
      {stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[49],stage2_14[54],stage2_13[83],stage2_12[85]}
   );
   gpc606_5 gpc2502 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209], stage1_12[210]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[50],stage2_14[55],stage2_13[84],stage2_12[86]}
   );
   gpc606_5 gpc2503 (
      {stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214], stage1_12[215], stage1_12[216]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[51],stage2_14[56],stage2_13[85],stage2_12[87]}
   );
   gpc606_5 gpc2504 (
      {stage1_12[217], stage1_12[218], stage1_12[219], stage1_12[220], stage1_12[221], stage1_12[222]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[52],stage2_14[57],stage2_13[86],stage2_12[88]}
   );
   gpc606_5 gpc2505 (
      {stage1_12[223], stage1_12[224], stage1_12[225], stage1_12[226], stage1_12[227], stage1_12[228]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[53],stage2_14[58],stage2_13[87],stage2_12[89]}
   );
   gpc606_5 gpc2506 (
      {stage1_12[229], stage1_12[230], stage1_12[231], stage1_12[232], stage1_12[233], stage1_12[234]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[54],stage2_14[59],stage2_13[88],stage2_12[90]}
   );
   gpc606_5 gpc2507 (
      {stage1_12[235], stage1_12[236], stage1_12[237], stage1_12[238], stage1_12[239], stage1_12[240]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[55],stage2_14[60],stage2_13[89],stage2_12[91]}
   );
   gpc606_5 gpc2508 (
      {stage1_12[241], stage1_12[242], stage1_12[243], stage1_12[244], stage1_12[245], stage1_12[246]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[56],stage2_14[61],stage2_13[90],stage2_12[92]}
   );
   gpc606_5 gpc2509 (
      {stage1_12[247], stage1_12[248], stage1_12[249], stage1_12[250], stage1_12[251], stage1_12[252]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[57],stage2_14[62],stage2_13[91],stage2_12[93]}
   );
   gpc606_5 gpc2510 (
      {stage1_12[253], stage1_12[254], stage1_12[255], stage1_12[256], stage1_12[257], stage1_12[258]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[58],stage2_14[63],stage2_13[92],stage2_12[94]}
   );
   gpc606_5 gpc2511 (
      {stage1_12[259], stage1_12[260], stage1_12[261], stage1_12[262], stage1_12[263], stage1_12[264]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[59],stage2_14[64],stage2_13[93],stage2_12[95]}
   );
   gpc606_5 gpc2512 (
      {stage1_12[265], stage1_12[266], stage1_12[267], stage1_12[268], stage1_12[269], stage1_12[270]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[60],stage2_14[65],stage2_13[94],stage2_12[96]}
   );
   gpc606_5 gpc2513 (
      {stage1_12[271], stage1_12[272], stage1_12[273], stage1_12[274], stage1_12[275], stage1_12[276]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[61],stage2_14[66],stage2_13[95],stage2_12[97]}
   );
   gpc606_5 gpc2514 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[33],stage2_15[62],stage2_14[67],stage2_13[96]}
   );
   gpc615_5 gpc2515 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[198]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[34],stage2_15[63],stage2_14[68],stage2_13[97]}
   );
   gpc615_5 gpc2516 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[199]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[35],stage2_15[64],stage2_14[69],stage2_13[98]}
   );
   gpc615_5 gpc2517 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[200]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[36],stage2_15[65],stage2_14[70],stage2_13[99]}
   );
   gpc615_5 gpc2518 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[201]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[37],stage2_15[66],stage2_14[71],stage2_13[100]}
   );
   gpc615_5 gpc2519 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[202]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[38],stage2_15[67],stage2_14[72],stage2_13[101]}
   );
   gpc615_5 gpc2520 (
      {stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207]},
      {stage1_15[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[6],stage2_16[39],stage2_15[68],stage2_14[73]}
   );
   gpc615_5 gpc2521 (
      {stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211], stage1_14[212]},
      {stage1_15[37]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[7],stage2_16[40],stage2_15[69],stage2_14[74]}
   );
   gpc615_5 gpc2522 (
      {stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216], stage1_14[217]},
      {stage1_15[38]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[8],stage2_16[41],stage2_15[70],stage2_14[75]}
   );
   gpc615_5 gpc2523 (
      {stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221], stage1_14[222]},
      {stage1_15[39]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[9],stage2_16[42],stage2_15[71],stage2_14[76]}
   );
   gpc615_5 gpc2524 (
      {stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226], stage1_14[227]},
      {stage1_15[40]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[10],stage2_16[43],stage2_15[72],stage2_14[77]}
   );
   gpc615_5 gpc2525 (
      {stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231], stage1_14[232]},
      {stage1_15[41]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[11],stage2_16[44],stage2_15[73],stage2_14[78]}
   );
   gpc615_5 gpc2526 (
      {stage1_14[233], stage1_14[234], stage1_14[235], stage1_14[236], stage1_14[237]},
      {stage1_15[42]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[12],stage2_16[45],stage2_15[74],stage2_14[79]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[42]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[46],stage2_15[75]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52]},
      {stage1_16[43]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[47],stage2_15[76]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[53], stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57]},
      {stage1_16[44]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[48],stage2_15[77]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62]},
      {stage1_16[45]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[49],stage2_15[78]}
   );
   gpc615_5 gpc2531 (
      {stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_16[46]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[50],stage2_15[79]}
   );
   gpc615_5 gpc2532 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72]},
      {stage1_16[47]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[51],stage2_15[80]}
   );
   gpc615_5 gpc2533 (
      {stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[48]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[52],stage2_15[81]}
   );
   gpc615_5 gpc2534 (
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82]},
      {stage1_16[49]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[53],stage2_15[82]}
   );
   gpc615_5 gpc2535 (
      {stage1_15[83], stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87]},
      {stage1_16[50]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[54],stage2_15[83]}
   );
   gpc615_5 gpc2536 (
      {stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91], stage1_15[92]},
      {stage1_16[51]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[55],stage2_15[84]}
   );
   gpc615_5 gpc2537 (
      {stage1_15[93], stage1_15[94], stage1_15[95], stage1_15[96], stage1_15[97]},
      {stage1_16[52]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[56],stage2_15[85]}
   );
   gpc615_5 gpc2538 (
      {stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101], stage1_15[102]},
      {stage1_16[53]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[57],stage2_15[86]}
   );
   gpc615_5 gpc2539 (
      {stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[54]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[19],stage2_17[25],stage2_16[58],stage2_15[87]}
   );
   gpc615_5 gpc2540 (
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112]},
      {stage1_16[55]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[20],stage2_17[26],stage2_16[59],stage2_15[88]}
   );
   gpc615_5 gpc2541 (
      {stage1_15[113], stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117]},
      {stage1_16[56]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[21],stage2_17[27],stage2_16[60],stage2_15[89]}
   );
   gpc615_5 gpc2542 (
      {stage1_15[118], stage1_15[119], stage1_15[120], stage1_15[121], stage1_15[122]},
      {stage1_16[57]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[22],stage2_17[28],stage2_16[61],stage2_15[90]}
   );
   gpc615_5 gpc2543 (
      {stage1_15[123], stage1_15[124], stage1_15[125], stage1_15[126], stage1_15[127]},
      {stage1_16[58]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[23],stage2_17[29],stage2_16[62],stage2_15[91]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[59], stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[24],stage2_17[30],stage2_16[63]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[25],stage2_17[31],stage2_16[64]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[26],stage2_17[32],stage2_16[65]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[27],stage2_17[33],stage2_16[66]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[28],stage2_17[34],stage2_16[67]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[89], stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[29],stage2_17[35],stage2_16[68]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[95], stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[30],stage2_17[36],stage2_16[69]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[101], stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[31],stage2_17[37],stage2_16[70]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[107], stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[32],stage2_17[38],stage2_16[71]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[113], stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[33],stage2_17[39],stage2_16[72]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[119], stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[34],stage2_17[40],stage2_16[73]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[125], stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[35],stage2_17[41],stage2_16[74]}
   );
   gpc606_5 gpc2556 (
      {stage1_16[131], stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[36],stage2_17[42],stage2_16[75]}
   );
   gpc606_5 gpc2557 (
      {stage1_16[137], stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[37],stage2_17[43],stage2_16[76]}
   );
   gpc606_5 gpc2558 (
      {stage1_16[143], stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[38],stage2_17[44],stage2_16[77]}
   );
   gpc606_5 gpc2559 (
      {stage1_16[149], stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[39],stage2_17[45],stage2_16[78]}
   );
   gpc606_5 gpc2560 (
      {stage1_16[155], stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[40],stage2_17[46],stage2_16[79]}
   );
   gpc606_5 gpc2561 (
      {stage1_16[161], stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[41],stage2_17[47],stage2_16[80]}
   );
   gpc606_5 gpc2562 (
      {stage1_16[167], stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[42],stage2_17[48],stage2_16[81]}
   );
   gpc606_5 gpc2563 (
      {stage1_16[173], stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[43],stage2_17[49],stage2_16[82]}
   );
   gpc606_5 gpc2564 (
      {stage1_16[179], stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[44],stage2_17[50],stage2_16[83]}
   );
   gpc606_5 gpc2565 (
      {stage1_16[185], stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[45],stage2_17[51],stage2_16[84]}
   );
   gpc606_5 gpc2566 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[46],stage2_17[52],stage2_16[85]}
   );
   gpc606_5 gpc2567 (
      {stage1_16[197], stage1_16[198], stage1_16[199], stage1_16[200], stage1_16[201], stage1_16[202]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[47],stage2_17[53],stage2_16[86]}
   );
   gpc606_5 gpc2568 (
      {stage1_16[203], stage1_16[204], stage1_16[205], stage1_16[206], stage1_16[207], stage1_16[208]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[48],stage2_17[54],stage2_16[87]}
   );
   gpc606_5 gpc2569 (
      {stage1_16[209], stage1_16[210], stage1_16[211], stage1_16[212], stage1_16[213], stage1_16[214]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[49],stage2_17[55],stage2_16[88]}
   );
   gpc606_5 gpc2570 (
      {stage1_16[215], stage1_16[216], stage1_16[217], stage1_16[218], stage1_16[219], stage1_16[220]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[50],stage2_17[56],stage2_16[89]}
   );
   gpc606_5 gpc2571 (
      {stage1_16[221], stage1_16[222], stage1_16[223], stage1_16[224], stage1_16[225], stage1_16[226]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[51],stage2_17[57],stage2_16[90]}
   );
   gpc606_5 gpc2572 (
      {stage1_16[227], stage1_16[228], stage1_16[229], stage1_16[230], stage1_16[231], stage1_16[232]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[52],stage2_17[58],stage2_16[91]}
   );
   gpc606_5 gpc2573 (
      {stage1_16[233], stage1_16[234], stage1_16[235], stage1_16[236], stage1_16[237], stage1_16[238]},
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage2_20[29],stage2_19[46],stage2_18[53],stage2_17[59],stage2_16[92]}
   );
   gpc606_5 gpc2574 (
      {stage1_16[239], stage1_16[240], stage1_16[241], stage1_16[242], stage1_16[243], stage1_16[244]},
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage2_20[30],stage2_19[47],stage2_18[54],stage2_17[60],stage2_16[93]}
   );
   gpc606_5 gpc2575 (
      {stage1_16[245], stage1_16[246], stage1_16[247], stage1_16[248], stage1_16[249], stage1_16[250]},
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190], stage1_18[191]},
      {stage2_20[31],stage2_19[48],stage2_18[55],stage2_17[61],stage2_16[94]}
   );
   gpc606_5 gpc2576 (
      {stage1_16[251], stage1_16[252], stage1_16[253], stage1_16[254], stage1_16[255], stage1_16[256]},
      {stage1_18[192], stage1_18[193], stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197]},
      {stage2_20[32],stage2_19[49],stage2_18[56],stage2_17[62],stage2_16[95]}
   );
   gpc606_5 gpc2577 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[33],stage2_19[50],stage2_18[57],stage2_17[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[34],stage2_19[51],stage2_18[58],stage2_17[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[35],stage2_19[52],stage2_18[59],stage2_17[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[36],stage2_19[53],stage2_18[60],stage2_17[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[37],stage2_19[54],stage2_18[61],stage2_17[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[38],stage2_19[55],stage2_18[62],stage2_17[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[39],stage2_19[56],stage2_18[63],stage2_17[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[40],stage2_19[57],stage2_18[64],stage2_17[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[41],stage2_19[58],stage2_18[65],stage2_17[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[42],stage2_19[59],stage2_18[66],stage2_17[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[43],stage2_19[60],stage2_18[67],stage2_17[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[44],stage2_19[61],stage2_18[68],stage2_17[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[45],stage2_19[62],stage2_18[69],stage2_17[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[46],stage2_19[63],stage2_18[70],stage2_17[76]}
   );
   gpc606_5 gpc2591 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[47],stage2_19[64],stage2_18[71],stage2_17[77]}
   );
   gpc606_5 gpc2592 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[48],stage2_19[65],stage2_18[72],stage2_17[78]}
   );
   gpc606_5 gpc2593 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[49],stage2_19[66],stage2_18[73],stage2_17[79]}
   );
   gpc606_5 gpc2594 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[50],stage2_19[67],stage2_18[74],stage2_17[80]}
   );
   gpc606_5 gpc2595 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[51],stage2_19[68],stage2_18[75],stage2_17[81]}
   );
   gpc606_5 gpc2596 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[52],stage2_19[69],stage2_18[76],stage2_17[82]}
   );
   gpc606_5 gpc2597 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[53],stage2_19[70],stage2_18[77],stage2_17[83]}
   );
   gpc606_5 gpc2598 (
      {stage1_17[228], stage1_17[229], stage1_17[230], stage1_17[231], stage1_17[232], stage1_17[233]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[54],stage2_19[71],stage2_18[78],stage2_17[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[22],stage2_20[55],stage2_19[72]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[23],stage2_20[56],stage2_19[73]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[24],stage2_20[57],stage2_19[74]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[147], stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[25],stage2_20[58],stage2_19[75]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155], stage1_19[156]},
      {stage1_20[4]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[26],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage1_20[5]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[27],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166]},
      {stage1_20[6]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[6],stage2_21[28],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171]},
      {stage1_20[7]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[7],stage2_21[29],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175], stage1_19[176]},
      {stage1_20[8]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[8],stage2_21[30],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180], stage1_19[181]},
      {stage1_20[9]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[9],stage2_21[31],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185], stage1_19[186]},
      {stage1_20[10]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[10],stage2_21[32],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2610 (
      {stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage1_20[11]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[11],stage2_21[33],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2611 (
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196]},
      {stage1_20[12]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[12],stage2_21[34],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2612 (
      {stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201]},
      {stage1_20[13]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[13],stage2_21[35],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2613 (
      {stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205], stage1_19[206]},
      {stage1_20[14]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[14],stage2_21[36],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2614 (
      {stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210], stage1_19[211]},
      {stage1_20[15]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[15],stage2_21[37],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2615 (
      {stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215], stage1_19[216]},
      {stage1_20[16]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[16],stage2_21[38],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2616 (
      {stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage1_20[17]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[17],stage2_21[39],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2617 (
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226]},
      {stage1_20[18]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[18],stage2_21[40],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2618 (
      {stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230], stage1_19[231]},
      {stage1_20[19]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[19],stage2_21[41],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2619 (
      {stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235], stage1_19[236]},
      {stage1_20[20]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[20],stage2_21[42],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2620 (
      {stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240], stage1_19[241]},
      {stage1_20[21]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[21],stage2_21[43],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2621 (
      {stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245], stage1_19[246]},
      {stage1_20[22]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[22],stage2_21[44],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2622 (
      {stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250], stage1_19[251]},
      {stage1_20[23]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[23],stage2_21[45],stage2_20[78],stage2_19[95]}
   );
   gpc615_5 gpc2623 (
      {stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255], stage1_19[256]},
      {stage1_20[24]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[24],stage2_21[46],stage2_20[79],stage2_19[96]}
   );
   gpc615_5 gpc2624 (
      {stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260], stage1_19[261]},
      {stage1_20[25]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[25],stage2_21[47],stage2_20[80],stage2_19[97]}
   );
   gpc615_5 gpc2625 (
      {stage1_19[262], stage1_19[263], stage1_19[264], stage1_19[265], stage1_19[266]},
      {stage1_20[26]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[26],stage2_21[48],stage2_20[81],stage2_19[98]}
   );
   gpc615_5 gpc2626 (
      {stage1_19[267], stage1_19[268], stage1_19[269], stage1_19[270], stage1_19[271]},
      {stage1_20[27]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[27],stage2_21[49],stage2_20[82],stage2_19[99]}
   );
   gpc615_5 gpc2627 (
      {stage1_19[272], stage1_19[273], stage1_19[274], stage1_19[275], stage1_19[276]},
      {stage1_20[28]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[28],stage2_21[50],stage2_20[83],stage2_19[100]}
   );
   gpc615_5 gpc2628 (
      {stage1_19[277], stage1_19[278], stage1_19[279], stage1_19[280], stage1_19[281]},
      {stage1_20[29]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[29],stage2_21[51],stage2_20[84],stage2_19[101]}
   );
   gpc615_5 gpc2629 (
      {stage1_19[282], stage1_19[283], stage1_19[284], stage1_19[285], stage1_19[286]},
      {stage1_20[30]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[30],stage2_21[52],stage2_20[85],stage2_19[102]}
   );
   gpc615_5 gpc2630 (
      {stage1_19[287], stage1_19[288], stage1_19[289], stage1_19[290], stage1_19[291]},
      {stage1_20[31]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[31],stage2_21[53],stage2_20[86],stage2_19[103]}
   );
   gpc623_5 gpc2631 (
      {stage1_19[292], stage1_19[293], stage1_19[294]},
      {stage1_20[32], stage1_20[33]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[32],stage2_21[54],stage2_20[87],stage2_19[104]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[34], stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[33],stage2_22[33],stage2_21[55],stage2_20[88]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[40], stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[34],stage2_22[34],stage2_21[56],stage2_20[89]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[46], stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[35],stage2_22[35],stage2_21[57],stage2_20[90]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[52], stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[36],stage2_22[36],stage2_21[58],stage2_20[91]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[58], stage1_20[59], stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[37],stage2_22[37],stage2_21[59],stage2_20[92]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[64], stage1_20[65], stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[38],stage2_22[38],stage2_21[60],stage2_20[93]}
   );
   gpc606_5 gpc2638 (
      {stage1_20[70], stage1_20[71], stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[39],stage2_22[39],stage2_21[61],stage2_20[94]}
   );
   gpc606_5 gpc2639 (
      {stage1_20[76], stage1_20[77], stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[40],stage2_22[40],stage2_21[62],stage2_20[95]}
   );
   gpc606_5 gpc2640 (
      {stage1_20[82], stage1_20[83], stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[41],stage2_22[41],stage2_21[63],stage2_20[96]}
   );
   gpc606_5 gpc2641 (
      {stage1_20[88], stage1_20[89], stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[42],stage2_22[42],stage2_21[64],stage2_20[97]}
   );
   gpc606_5 gpc2642 (
      {stage1_20[94], stage1_20[95], stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[43],stage2_22[43],stage2_21[65],stage2_20[98]}
   );
   gpc606_5 gpc2643 (
      {stage1_20[100], stage1_20[101], stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[44],stage2_22[44],stage2_21[66],stage2_20[99]}
   );
   gpc606_5 gpc2644 (
      {stage1_20[106], stage1_20[107], stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[45],stage2_22[45],stage2_21[67],stage2_20[100]}
   );
   gpc606_5 gpc2645 (
      {stage1_20[112], stage1_20[113], stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[46],stage2_22[46],stage2_21[68],stage2_20[101]}
   );
   gpc606_5 gpc2646 (
      {stage1_20[118], stage1_20[119], stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[47],stage2_22[47],stage2_21[69],stage2_20[102]}
   );
   gpc606_5 gpc2647 (
      {stage1_20[124], stage1_20[125], stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[48],stage2_22[48],stage2_21[70],stage2_20[103]}
   );
   gpc606_5 gpc2648 (
      {stage1_20[130], stage1_20[131], stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[49],stage2_22[49],stage2_21[71],stage2_20[104]}
   );
   gpc606_5 gpc2649 (
      {stage1_20[136], stage1_20[137], stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[50],stage2_22[50],stage2_21[72],stage2_20[105]}
   );
   gpc606_5 gpc2650 (
      {stage1_20[142], stage1_20[143], stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[51],stage2_22[51],stage2_21[73],stage2_20[106]}
   );
   gpc606_5 gpc2651 (
      {stage1_20[148], stage1_20[149], stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[52],stage2_22[52],stage2_21[74],stage2_20[107]}
   );
   gpc606_5 gpc2652 (
      {stage1_20[154], stage1_20[155], stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[53],stage2_22[53],stage2_21[75],stage2_20[108]}
   );
   gpc606_5 gpc2653 (
      {stage1_20[160], stage1_20[161], stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[54],stage2_22[54],stage2_21[76],stage2_20[109]}
   );
   gpc606_5 gpc2654 (
      {stage1_20[166], stage1_20[167], stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[55],stage2_22[55],stage2_21[77],stage2_20[110]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142]},
      {stage1_23[0]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[0],stage2_24[23],stage2_23[56],stage2_22[56]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[143], stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147]},
      {stage1_23[1]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[1],stage2_24[24],stage2_23[57],stage2_22[57]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[148], stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152]},
      {stage1_23[2]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[2],stage2_24[25],stage2_23[58],stage2_22[58]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[153], stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157]},
      {stage1_23[3]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[3],stage2_24[26],stage2_23[59],stage2_22[59]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162]},
      {stage1_23[4]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[4],stage2_24[27],stage2_23[60],stage2_22[60]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage1_23[5]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[5],stage2_24[28],stage2_23[61],stage2_22[61]}
   );
   gpc615_5 gpc2661 (
      {stage1_22[168], stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172]},
      {stage1_23[6]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[6],stage2_24[29],stage2_23[62],stage2_22[62]}
   );
   gpc615_5 gpc2662 (
      {stage1_22[173], stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177]},
      {stage1_23[7]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[7],stage2_24[30],stage2_23[63],stage2_22[63]}
   );
   gpc615_5 gpc2663 (
      {stage1_22[178], stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182]},
      {stage1_23[8]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[8],stage2_24[31],stage2_23[64],stage2_22[64]}
   );
   gpc615_5 gpc2664 (
      {stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187]},
      {stage1_23[9]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[9],stage2_24[32],stage2_23[65],stage2_22[65]}
   );
   gpc615_5 gpc2665 (
      {stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_23[10]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[10],stage2_24[33],stage2_23[66],stage2_22[66]}
   );
   gpc615_5 gpc2666 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[11]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[11],stage2_24[34],stage2_23[67],stage2_22[67]}
   );
   gpc615_5 gpc2667 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[12]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[12],stage2_24[35],stage2_23[68],stage2_22[68]}
   );
   gpc615_5 gpc2668 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[13]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[13],stage2_24[36],stage2_23[69],stage2_22[69]}
   );
   gpc615_5 gpc2669 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[14]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[14],stage2_24[37],stage2_23[70],stage2_22[70]}
   );
   gpc615_5 gpc2670 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[15]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[15],stage2_24[38],stage2_23[71],stage2_22[71]}
   );
   gpc615_5 gpc2671 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[16]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[16],stage2_24[39],stage2_23[72],stage2_22[72]}
   );
   gpc615_5 gpc2672 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[17]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[17],stage2_24[40],stage2_23[73],stage2_22[73]}
   );
   gpc615_5 gpc2673 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[18]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[18],stage2_24[41],stage2_23[74],stage2_22[74]}
   );
   gpc615_5 gpc2674 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[19]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[19],stage2_24[42],stage2_23[75],stage2_22[75]}
   );
   gpc615_5 gpc2675 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[20]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[20],stage2_24[43],stage2_23[76],stage2_22[76]}
   );
   gpc615_5 gpc2676 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[21]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[21],stage2_24[44],stage2_23[77],stage2_22[77]}
   );
   gpc615_5 gpc2677 (
      {stage1_22[248], stage1_22[249], stage1_22[250], 1'b0, 1'b0},
      {stage1_23[22]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[22],stage2_24[45],stage2_23[78],stage2_22[78]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[23], stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27]},
      {stage1_24[138]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[23],stage2_25[23],stage2_24[46],stage2_23[79]}
   );
   gpc615_5 gpc2679 (
      {stage1_23[28], stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32]},
      {stage1_24[139]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[24],stage2_25[24],stage2_24[47],stage2_23[80]}
   );
   gpc615_5 gpc2680 (
      {stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36], stage1_23[37]},
      {stage1_24[140]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[25],stage2_25[25],stage2_24[48],stage2_23[81]}
   );
   gpc615_5 gpc2681 (
      {stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_24[141]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[26],stage2_25[26],stage2_24[49],stage2_23[82]}
   );
   gpc615_5 gpc2682 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[142]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[27],stage2_25[27],stage2_24[50],stage2_23[83]}
   );
   gpc615_5 gpc2683 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52]},
      {stage1_24[143]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[28],stage2_25[28],stage2_24[51],stage2_23[84]}
   );
   gpc615_5 gpc2684 (
      {stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57]},
      {stage1_24[144]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[29],stage2_25[29],stage2_24[52],stage2_23[85]}
   );
   gpc615_5 gpc2685 (
      {stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_24[145]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[30],stage2_25[30],stage2_24[53],stage2_23[86]}
   );
   gpc615_5 gpc2686 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67]},
      {stage1_24[146]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[31],stage2_25[31],stage2_24[54],stage2_23[87]}
   );
   gpc615_5 gpc2687 (
      {stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_24[147]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[32],stage2_25[32],stage2_24[55],stage2_23[88]}
   );
   gpc615_5 gpc2688 (
      {stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_24[148]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[33],stage2_25[33],stage2_24[56],stage2_23[89]}
   );
   gpc615_5 gpc2689 (
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82]},
      {stage1_24[149]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[34],stage2_25[34],stage2_24[57],stage2_23[90]}
   );
   gpc615_5 gpc2690 (
      {stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87]},
      {stage1_24[150]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[35],stage2_25[35],stage2_24[58],stage2_23[91]}
   );
   gpc615_5 gpc2691 (
      {stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_24[151]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[36],stage2_25[36],stage2_24[59],stage2_23[92]}
   );
   gpc615_5 gpc2692 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97]},
      {stage1_24[152]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[37],stage2_25[37],stage2_24[60],stage2_23[93]}
   );
   gpc615_5 gpc2693 (
      {stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_24[153]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[38],stage2_25[38],stage2_24[61],stage2_23[94]}
   );
   gpc615_5 gpc2694 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage1_24[154]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[39],stage2_25[39],stage2_24[62],stage2_23[95]}
   );
   gpc615_5 gpc2695 (
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112]},
      {stage1_24[155]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[40],stage2_25[40],stage2_24[63],stage2_23[96]}
   );
   gpc615_5 gpc2696 (
      {stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117]},
      {stage1_24[156]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[41],stage2_25[41],stage2_24[64],stage2_23[97]}
   );
   gpc615_5 gpc2697 (
      {stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_24[157]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[42],stage2_25[42],stage2_24[65],stage2_23[98]}
   );
   gpc615_5 gpc2698 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127]},
      {stage1_24[158]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[43],stage2_25[43],stage2_24[66],stage2_23[99]}
   );
   gpc615_5 gpc2699 (
      {stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132]},
      {stage1_24[159]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[44],stage2_25[44],stage2_24[67],stage2_23[100]}
   );
   gpc615_5 gpc2700 (
      {stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage1_24[160]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[45],stage2_25[45],stage2_24[68],stage2_23[101]}
   );
   gpc615_5 gpc2701 (
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142]},
      {stage1_24[161]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[46],stage2_25[46],stage2_24[69],stage2_23[102]}
   );
   gpc615_5 gpc2702 (
      {stage1_23[143], stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147]},
      {stage1_24[162]},
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage2_27[24],stage2_26[47],stage2_25[47],stage2_24[70],stage2_23[103]}
   );
   gpc615_5 gpc2703 (
      {stage1_23[148], stage1_23[149], stage1_23[150], stage1_23[151], stage1_23[152]},
      {stage1_24[163]},
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage2_27[25],stage2_26[48],stage2_25[48],stage2_24[71],stage2_23[104]}
   );
   gpc615_5 gpc2704 (
      {stage1_23[153], stage1_23[154], stage1_23[155], stage1_23[156], stage1_23[157]},
      {stage1_24[164]},
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage2_27[26],stage2_26[49],stage2_25[49],stage2_24[72],stage2_23[105]}
   );
   gpc615_5 gpc2705 (
      {stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161], stage1_23[162]},
      {stage1_24[165]},
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage2_27[27],stage2_26[50],stage2_25[50],stage2_24[73],stage2_23[106]}
   );
   gpc615_5 gpc2706 (
      {stage1_23[163], stage1_23[164], stage1_23[165], stage1_23[166], stage1_23[167]},
      {stage1_24[166]},
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage2_27[28],stage2_26[51],stage2_25[51],stage2_24[74],stage2_23[107]}
   );
   gpc615_5 gpc2707 (
      {stage1_23[168], stage1_23[169], stage1_23[170], stage1_23[171], stage1_23[172]},
      {stage1_24[167]},
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage2_27[29],stage2_26[52],stage2_25[52],stage2_24[75],stage2_23[108]}
   );
   gpc615_5 gpc2708 (
      {stage1_23[173], stage1_23[174], stage1_23[175], stage1_23[176], stage1_23[177]},
      {stage1_24[168]},
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage2_27[30],stage2_26[53],stage2_25[53],stage2_24[76],stage2_23[109]}
   );
   gpc615_5 gpc2709 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[186]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[31],stage2_26[54],stage2_25[54],stage2_24[77]}
   );
   gpc615_5 gpc2710 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[187]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[32],stage2_26[55],stage2_25[55],stage2_24[78]}
   );
   gpc615_5 gpc2711 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[188]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[33],stage2_26[56],stage2_25[56],stage2_24[79]}
   );
   gpc615_5 gpc2712 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[189]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[34],stage2_26[57],stage2_25[57],stage2_24[80]}
   );
   gpc615_5 gpc2713 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[190]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[35],stage2_26[58],stage2_25[58],stage2_24[81]}
   );
   gpc606_5 gpc2714 (
      {stage1_25[191], stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[5],stage2_27[36],stage2_26[59],stage2_25[59]}
   );
   gpc606_5 gpc2715 (
      {stage1_25[197], stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[6],stage2_27[37],stage2_26[60],stage2_25[60]}
   );
   gpc606_5 gpc2716 (
      {stage1_25[203], stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[7],stage2_27[38],stage2_26[61],stage2_25[61]}
   );
   gpc615_5 gpc2717 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34]},
      {stage1_27[18]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[3],stage2_28[8],stage2_27[39],stage2_26[62]}
   );
   gpc615_5 gpc2718 (
      {stage1_26[35], stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39]},
      {stage1_27[19]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[4],stage2_28[9],stage2_27[40],stage2_26[63]}
   );
   gpc615_5 gpc2719 (
      {stage1_26[40], stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44]},
      {stage1_27[20]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[5],stage2_28[10],stage2_27[41],stage2_26[64]}
   );
   gpc615_5 gpc2720 (
      {stage1_26[45], stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49]},
      {stage1_27[21]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[6],stage2_28[11],stage2_27[42],stage2_26[65]}
   );
   gpc615_5 gpc2721 (
      {stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54]},
      {stage1_27[22]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[7],stage2_28[12],stage2_27[43],stage2_26[66]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage1_27[23]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[8],stage2_28[13],stage2_27[44],stage2_26[67]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64]},
      {stage1_27[24]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[9],stage2_28[14],stage2_27[45],stage2_26[68]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69]},
      {stage1_27[25]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[10],stage2_28[15],stage2_27[46],stage2_26[69]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74]},
      {stage1_27[26]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[11],stage2_28[16],stage2_27[47],stage2_26[70]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[75], stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79]},
      {stage1_27[27]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[12],stage2_28[17],stage2_27[48],stage2_26[71]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84]},
      {stage1_27[28]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[13],stage2_28[18],stage2_27[49],stage2_26[72]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage1_27[29]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[14],stage2_28[19],stage2_27[50],stage2_26[73]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94]},
      {stage1_27[30]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[15],stage2_28[20],stage2_27[51],stage2_26[74]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[95], stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99]},
      {stage1_27[31]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[16],stage2_28[21],stage2_27[52],stage2_26[75]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[100], stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104]},
      {stage1_27[32]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[17],stage2_28[22],stage2_27[53],stage2_26[76]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[105], stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109]},
      {stage1_27[33]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[18],stage2_28[23],stage2_27[54],stage2_26[77]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114]},
      {stage1_27[34]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[19],stage2_28[24],stage2_27[55],stage2_26[78]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage1_27[35]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[20],stage2_28[25],stage2_27[56],stage2_26[79]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124]},
      {stage1_27[36]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[21],stage2_28[26],stage2_27[57],stage2_26[80]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[125], stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129]},
      {stage1_27[37]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[22],stage2_28[27],stage2_27[58],stage2_26[81]}
   );
   gpc615_5 gpc2737 (
      {stage1_26[130], stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134]},
      {stage1_27[38]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[23],stage2_28[28],stage2_27[59],stage2_26[82]}
   );
   gpc615_5 gpc2738 (
      {stage1_26[135], stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139]},
      {stage1_27[39]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[24],stage2_28[29],stage2_27[60],stage2_26[83]}
   );
   gpc615_5 gpc2739 (
      {stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144]},
      {stage1_27[40]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[25],stage2_28[30],stage2_27[61],stage2_26[84]}
   );
   gpc615_5 gpc2740 (
      {stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage1_27[41]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[26],stage2_28[31],stage2_27[62],stage2_26[85]}
   );
   gpc615_5 gpc2741 (
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154]},
      {stage1_27[42]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[27],stage2_28[32],stage2_27[63],stage2_26[86]}
   );
   gpc615_5 gpc2742 (
      {stage1_26[155], stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159]},
      {stage1_27[43]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[28],stage2_28[33],stage2_27[64],stage2_26[87]}
   );
   gpc615_5 gpc2743 (
      {stage1_26[160], stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164]},
      {stage1_27[44]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[29],stage2_28[34],stage2_27[65],stage2_26[88]}
   );
   gpc615_5 gpc2744 (
      {stage1_26[165], stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169]},
      {stage1_27[45]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[30],stage2_28[35],stage2_27[66],stage2_26[89]}
   );
   gpc615_5 gpc2745 (
      {stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174]},
      {stage1_27[46]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[31],stage2_28[36],stage2_27[67],stage2_26[90]}
   );
   gpc615_5 gpc2746 (
      {stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage1_27[47]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[32],stage2_28[37],stage2_27[68],stage2_26[91]}
   );
   gpc615_5 gpc2747 (
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184]},
      {stage1_27[48]},
      {stage1_28[180], stage1_28[181], stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185]},
      {stage2_30[30],stage2_29[33],stage2_28[38],stage2_27[69],stage2_26[92]}
   );
   gpc615_5 gpc2748 (
      {stage1_26[185], stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189]},
      {stage1_27[49]},
      {stage1_28[186], stage1_28[187], stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191]},
      {stage2_30[31],stage2_29[34],stage2_28[39],stage2_27[70],stage2_26[93]}
   );
   gpc615_5 gpc2749 (
      {stage1_26[190], stage1_26[191], stage1_26[192], stage1_26[193], stage1_26[194]},
      {stage1_27[50]},
      {stage1_28[192], stage1_28[193], stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197]},
      {stage2_30[32],stage2_29[35],stage2_28[40],stage2_27[71],stage2_26[94]}
   );
   gpc615_5 gpc2750 (
      {stage1_26[195], stage1_26[196], stage1_26[197], stage1_26[198], stage1_26[199]},
      {stage1_27[51]},
      {stage1_28[198], stage1_28[199], stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203]},
      {stage2_30[33],stage2_29[36],stage2_28[41],stage2_27[72],stage2_26[95]}
   );
   gpc615_5 gpc2751 (
      {stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203], stage1_26[204]},
      {stage1_27[52]},
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage2_30[34],stage2_29[37],stage2_28[42],stage2_27[73],stage2_26[96]}
   );
   gpc615_5 gpc2752 (
      {stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208], stage1_26[209]},
      {stage1_27[53]},
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage2_30[35],stage2_29[38],stage2_28[43],stage2_27[74],stage2_26[97]}
   );
   gpc615_5 gpc2753 (
      {stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213], stage1_26[214]},
      {stage1_27[54]},
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage2_30[36],stage2_29[39],stage2_28[44],stage2_27[75],stage2_26[98]}
   );
   gpc615_5 gpc2754 (
      {stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage1_28[222]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[37],stage2_29[40],stage2_28[45],stage2_27[76]}
   );
   gpc615_5 gpc2755 (
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64]},
      {stage1_28[223]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[38],stage2_29[41],stage2_28[46],stage2_27[77]}
   );
   gpc615_5 gpc2756 (
      {stage1_27[65], stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69]},
      {stage1_28[224]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[39],stage2_29[42],stage2_28[47],stage2_27[78]}
   );
   gpc615_5 gpc2757 (
      {stage1_27[70], stage1_27[71], stage1_27[72], stage1_27[73], stage1_27[74]},
      {stage1_28[225]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[40],stage2_29[43],stage2_28[48],stage2_27[79]}
   );
   gpc615_5 gpc2758 (
      {stage1_27[75], stage1_27[76], stage1_27[77], stage1_27[78], stage1_27[79]},
      {stage1_28[226]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[41],stage2_29[44],stage2_28[49],stage2_27[80]}
   );
   gpc615_5 gpc2759 (
      {stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83], stage1_27[84]},
      {stage1_28[227]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[42],stage2_29[45],stage2_28[50],stage2_27[81]}
   );
   gpc615_5 gpc2760 (
      {stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage1_28[228]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[43],stage2_29[46],stage2_28[51],stage2_27[82]}
   );
   gpc615_5 gpc2761 (
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94]},
      {stage1_28[229]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[44],stage2_29[47],stage2_28[52],stage2_27[83]}
   );
   gpc615_5 gpc2762 (
      {stage1_27[95], stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99]},
      {stage1_28[230]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[45],stage2_29[48],stage2_28[53],stage2_27[84]}
   );
   gpc615_5 gpc2763 (
      {stage1_27[100], stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104]},
      {stage1_28[231]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[46],stage2_29[49],stage2_28[54],stage2_27[85]}
   );
   gpc615_5 gpc2764 (
      {stage1_27[105], stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109]},
      {stage1_28[232]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[47],stage2_29[50],stage2_28[55],stage2_27[86]}
   );
   gpc615_5 gpc2765 (
      {stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114]},
      {stage1_28[233]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[48],stage2_29[51],stage2_28[56],stage2_27[87]}
   );
   gpc615_5 gpc2766 (
      {stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage1_28[234]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[49],stage2_29[52],stage2_28[57],stage2_27[88]}
   );
   gpc615_5 gpc2767 (
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124]},
      {stage1_28[235]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[50],stage2_29[53],stage2_28[58],stage2_27[89]}
   );
   gpc615_5 gpc2768 (
      {stage1_27[125], stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129]},
      {stage1_28[236]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[51],stage2_29[54],stage2_28[59],stage2_27[90]}
   );
   gpc615_5 gpc2769 (
      {stage1_27[130], stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134]},
      {stage1_28[237]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[52],stage2_29[55],stage2_28[60],stage2_27[91]}
   );
   gpc615_5 gpc2770 (
      {stage1_27[135], stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139]},
      {stage1_28[238]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[53],stage2_29[56],stage2_28[61],stage2_27[92]}
   );
   gpc615_5 gpc2771 (
      {stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144]},
      {stage1_28[239]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[54],stage2_29[57],stage2_28[62],stage2_27[93]}
   );
   gpc615_5 gpc2772 (
      {stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage1_28[240]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[55],stage2_29[58],stage2_28[63],stage2_27[94]}
   );
   gpc615_5 gpc2773 (
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154]},
      {stage1_28[241]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[56],stage2_29[59],stage2_28[64],stage2_27[95]}
   );
   gpc615_5 gpc2774 (
      {stage1_27[155], stage1_27[156], stage1_27[157], stage1_27[158], 1'b0},
      {stage1_28[242]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[57],stage2_29[60],stage2_28[65],stage2_27[96]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[0],stage2_31[21],stage2_30[58],stage2_29[61]}
   );
   gpc606_5 gpc2776 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[1],stage2_31[22],stage2_30[59],stage2_29[62]}
   );
   gpc606_5 gpc2777 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[2],stage2_31[23],stage2_30[60],stage2_29[63]}
   );
   gpc606_5 gpc2778 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[3],stage2_31[24],stage2_30[61],stage2_29[64]}
   );
   gpc606_5 gpc2779 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[4],stage2_31[25],stage2_30[62],stage2_29[65]}
   );
   gpc606_5 gpc2780 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[5],stage2_31[26],stage2_30[63],stage2_29[66]}
   );
   gpc606_5 gpc2781 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[6],stage2_31[27],stage2_30[64],stage2_29[67]}
   );
   gpc606_5 gpc2782 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[7],stage2_31[28],stage2_30[65],stage2_29[68]}
   );
   gpc606_5 gpc2783 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[8],stage2_31[29],stage2_30[66],stage2_29[69]}
   );
   gpc606_5 gpc2784 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[9],stage2_31[30],stage2_30[67],stage2_29[70]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[10],stage2_32[10],stage2_31[31],stage2_30[68]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[11],stage2_32[11],stage2_31[32],stage2_30[69]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[12],stage2_32[12],stage2_31[33],stage2_30[70]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[13],stage2_32[13],stage2_31[34],stage2_30[71]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[14],stage2_32[14],stage2_31[35],stage2_30[72]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[15],stage2_32[15],stage2_31[36],stage2_30[73]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[16],stage2_32[16],stage2_31[37],stage2_30[74]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[17],stage2_32[17],stage2_31[38],stage2_30[75]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[18],stage2_32[18],stage2_31[39],stage2_30[76]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[19],stage2_32[19],stage2_31[40],stage2_30[77]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[20],stage2_32[20],stage2_31[41],stage2_30[78]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[21],stage2_32[21],stage2_31[42],stage2_30[79]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[22],stage2_32[22],stage2_31[43],stage2_30[80]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[23],stage2_32[23],stage2_31[44],stage2_30[81]}
   );
   gpc606_5 gpc2799 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[24],stage2_32[24],stage2_31[45],stage2_30[82]}
   );
   gpc606_5 gpc2800 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[25],stage2_32[25],stage2_31[46],stage2_30[83]}
   );
   gpc606_5 gpc2801 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[26],stage2_32[26],stage2_31[47],stage2_30[84]}
   );
   gpc606_5 gpc2802 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[27],stage2_32[27],stage2_31[48],stage2_30[85]}
   );
   gpc606_5 gpc2803 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[28],stage2_32[28],stage2_31[49],stage2_30[86]}
   );
   gpc606_5 gpc2804 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[29],stage2_32[29],stage2_31[50],stage2_30[87]}
   );
   gpc606_5 gpc2805 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[30],stage2_32[30],stage2_31[51],stage2_30[88]}
   );
   gpc606_5 gpc2806 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[31],stage2_32[31],stage2_31[52],stage2_30[89]}
   );
   gpc606_5 gpc2807 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[22],stage2_33[32],stage2_32[32],stage2_31[53]}
   );
   gpc606_5 gpc2808 (
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[23],stage2_33[33],stage2_32[33],stage2_31[54]}
   );
   gpc606_5 gpc2809 (
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[24],stage2_33[34],stage2_32[34],stage2_31[55]}
   );
   gpc606_5 gpc2810 (
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[25],stage2_33[35],stage2_32[35],stage2_31[56]}
   );
   gpc606_5 gpc2811 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[26],stage2_33[36],stage2_32[36],stage2_31[57]}
   );
   gpc606_5 gpc2812 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[27],stage2_33[37],stage2_32[37],stage2_31[58]}
   );
   gpc606_5 gpc2813 (
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[28],stage2_33[38],stage2_32[38],stage2_31[59]}
   );
   gpc606_5 gpc2814 (
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[29],stage2_33[39],stage2_32[39],stage2_31[60]}
   );
   gpc606_5 gpc2815 (
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[30],stage2_33[40],stage2_32[40],stage2_31[61]}
   );
   gpc606_5 gpc2816 (
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[31],stage2_33[41],stage2_32[41],stage2_31[62]}
   );
   gpc606_5 gpc2817 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[32],stage2_33[42],stage2_32[42],stage2_31[63]}
   );
   gpc606_5 gpc2818 (
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[33],stage2_33[43],stage2_32[43],stage2_31[64]}
   );
   gpc606_5 gpc2819 (
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[34],stage2_33[44],stage2_32[44],stage2_31[65]}
   );
   gpc606_5 gpc2820 (
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage1_33[78], stage1_33[79], stage1_33[80], 1'b0, 1'b0, 1'b0},
      {stage2_35[13],stage2_34[35],stage2_33[45],stage2_32[45],stage2_31[66]}
   );
   gpc1_1 gpc2821 (
      {stage1_1[62]},
      {stage2_1[31]}
   );
   gpc1_1 gpc2822 (
      {stage1_1[63]},
      {stage2_1[32]}
   );
   gpc1_1 gpc2823 (
      {stage1_1[64]},
      {stage2_1[33]}
   );
   gpc1_1 gpc2824 (
      {stage1_1[65]},
      {stage2_1[34]}
   );
   gpc1_1 gpc2825 (
      {stage1_1[66]},
      {stage2_1[35]}
   );
   gpc1_1 gpc2826 (
      {stage1_1[67]},
      {stage2_1[36]}
   );
   gpc1_1 gpc2827 (
      {stage1_1[68]},
      {stage2_1[37]}
   );
   gpc1_1 gpc2828 (
      {stage1_1[69]},
      {stage2_1[38]}
   );
   gpc1_1 gpc2829 (
      {stage1_1[70]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2830 (
      {stage1_1[71]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2831 (
      {stage1_1[72]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2832 (
      {stage1_1[73]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2833 (
      {stage1_1[74]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2834 (
      {stage1_1[75]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2835 (
      {stage1_1[76]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2836 (
      {stage1_1[77]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2837 (
      {stage1_1[78]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2838 (
      {stage1_1[79]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2839 (
      {stage1_1[80]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2840 (
      {stage1_1[81]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2841 (
      {stage1_1[82]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2842 (
      {stage1_1[83]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2843 (
      {stage1_1[84]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2844 (
      {stage1_1[85]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2845 (
      {stage1_1[86]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2846 (
      {stage1_1[87]},
      {stage2_1[56]}
   );
   gpc1_1 gpc2847 (
      {stage1_1[88]},
      {stage2_1[57]}
   );
   gpc1_1 gpc2848 (
      {stage1_1[89]},
      {stage2_1[58]}
   );
   gpc1_1 gpc2849 (
      {stage1_1[90]},
      {stage2_1[59]}
   );
   gpc1_1 gpc2850 (
      {stage1_1[91]},
      {stage2_1[60]}
   );
   gpc1_1 gpc2851 (
      {stage1_1[92]},
      {stage2_1[61]}
   );
   gpc1_1 gpc2852 (
      {stage1_1[93]},
      {stage2_1[62]}
   );
   gpc1_1 gpc2853 (
      {stage1_1[94]},
      {stage2_1[63]}
   );
   gpc1_1 gpc2854 (
      {stage1_1[95]},
      {stage2_1[64]}
   );
   gpc1_1 gpc2855 (
      {stage1_1[96]},
      {stage2_1[65]}
   );
   gpc1_1 gpc2856 (
      {stage1_1[97]},
      {stage2_1[66]}
   );
   gpc1_1 gpc2857 (
      {stage1_1[98]},
      {stage2_1[67]}
   );
   gpc1_1 gpc2858 (
      {stage1_1[99]},
      {stage2_1[68]}
   );
   gpc1_1 gpc2859 (
      {stage1_1[100]},
      {stage2_1[69]}
   );
   gpc1_1 gpc2860 (
      {stage1_1[101]},
      {stage2_1[70]}
   );
   gpc1_1 gpc2861 (
      {stage1_1[102]},
      {stage2_1[71]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[103]},
      {stage2_1[72]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[104]},
      {stage2_1[73]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[105]},
      {stage2_1[74]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[106]},
      {stage2_1[75]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[107]},
      {stage2_1[76]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[108]},
      {stage2_1[77]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[109]},
      {stage2_1[78]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[110]},
      {stage2_1[79]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[111]},
      {stage2_1[80]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[112]},
      {stage2_1[81]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[113]},
      {stage2_1[82]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[114]},
      {stage2_1[83]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[115]},
      {stage2_1[84]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[116]},
      {stage2_1[85]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[117]},
      {stage2_1[86]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[118]},
      {stage2_1[87]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[119]},
      {stage2_1[88]}
   );
   gpc1_1 gpc2879 (
      {stage1_1[120]},
      {stage2_1[89]}
   );
   gpc1_1 gpc2880 (
      {stage1_1[121]},
      {stage2_1[90]}
   );
   gpc1_1 gpc2881 (
      {stage1_1[122]},
      {stage2_1[91]}
   );
   gpc1_1 gpc2882 (
      {stage1_1[123]},
      {stage2_1[92]}
   );
   gpc1_1 gpc2883 (
      {stage1_1[124]},
      {stage2_1[93]}
   );
   gpc1_1 gpc2884 (
      {stage1_1[125]},
      {stage2_1[94]}
   );
   gpc1_1 gpc2885 (
      {stage1_1[126]},
      {stage2_1[95]}
   );
   gpc1_1 gpc2886 (
      {stage1_1[127]},
      {stage2_1[96]}
   );
   gpc1_1 gpc2887 (
      {stage1_1[128]},
      {stage2_1[97]}
   );
   gpc1_1 gpc2888 (
      {stage1_1[129]},
      {stage2_1[98]}
   );
   gpc1_1 gpc2889 (
      {stage1_1[130]},
      {stage2_1[99]}
   );
   gpc1_1 gpc2890 (
      {stage1_1[131]},
      {stage2_1[100]}
   );
   gpc1_1 gpc2891 (
      {stage1_1[132]},
      {stage2_1[101]}
   );
   gpc1_1 gpc2892 (
      {stage1_1[133]},
      {stage2_1[102]}
   );
   gpc1_1 gpc2893 (
      {stage1_1[134]},
      {stage2_1[103]}
   );
   gpc1_1 gpc2894 (
      {stage1_1[135]},
      {stage2_1[104]}
   );
   gpc1_1 gpc2895 (
      {stage1_1[136]},
      {stage2_1[105]}
   );
   gpc1_1 gpc2896 (
      {stage1_1[137]},
      {stage2_1[106]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[225]},
      {stage2_2[48]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[226]},
      {stage2_2[49]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[227]},
      {stage2_2[50]}
   );
   gpc1_1 gpc2900 (
      {stage1_3[169]},
      {stage2_3[69]}
   );
   gpc1_1 gpc2901 (
      {stage1_3[170]},
      {stage2_3[70]}
   );
   gpc1_1 gpc2902 (
      {stage1_3[171]},
      {stage2_3[71]}
   );
   gpc1_1 gpc2903 (
      {stage1_3[172]},
      {stage2_3[72]}
   );
   gpc1_1 gpc2904 (
      {stage1_3[173]},
      {stage2_3[73]}
   );
   gpc1_1 gpc2905 (
      {stage1_3[174]},
      {stage2_3[74]}
   );
   gpc1_1 gpc2906 (
      {stage1_3[175]},
      {stage2_3[75]}
   );
   gpc1_1 gpc2907 (
      {stage1_3[176]},
      {stage2_3[76]}
   );
   gpc1_1 gpc2908 (
      {stage1_3[177]},
      {stage2_3[77]}
   );
   gpc1_1 gpc2909 (
      {stage1_3[178]},
      {stage2_3[78]}
   );
   gpc1_1 gpc2910 (
      {stage1_3[179]},
      {stage2_3[79]}
   );
   gpc1_1 gpc2911 (
      {stage1_3[180]},
      {stage2_3[80]}
   );
   gpc1_1 gpc2912 (
      {stage1_3[181]},
      {stage2_3[81]}
   );
   gpc1_1 gpc2913 (
      {stage1_3[182]},
      {stage2_3[82]}
   );
   gpc1_1 gpc2914 (
      {stage1_3[183]},
      {stage2_3[83]}
   );
   gpc1_1 gpc2915 (
      {stage1_3[184]},
      {stage2_3[84]}
   );
   gpc1_1 gpc2916 (
      {stage1_3[185]},
      {stage2_3[85]}
   );
   gpc1_1 gpc2917 (
      {stage1_3[186]},
      {stage2_3[86]}
   );
   gpc1_1 gpc2918 (
      {stage1_3[187]},
      {stage2_3[87]}
   );
   gpc1_1 gpc2919 (
      {stage1_5[213]},
      {stage2_5[79]}
   );
   gpc1_1 gpc2920 (
      {stage1_5[214]},
      {stage2_5[80]}
   );
   gpc1_1 gpc2921 (
      {stage1_5[215]},
      {stage2_5[81]}
   );
   gpc1_1 gpc2922 (
      {stage1_5[216]},
      {stage2_5[82]}
   );
   gpc1_1 gpc2923 (
      {stage1_5[217]},
      {stage2_5[83]}
   );
   gpc1_1 gpc2924 (
      {stage1_7[218]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2925 (
      {stage1_7[219]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2926 (
      {stage1_7[220]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2927 (
      {stage1_7[221]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2928 (
      {stage1_7[222]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2929 (
      {stage1_7[223]},
      {stage2_7[109]}
   );
   gpc1_1 gpc2930 (
      {stage1_8[183]},
      {stage2_8[85]}
   );
   gpc1_1 gpc2931 (
      {stage1_8[184]},
      {stage2_8[86]}
   );
   gpc1_1 gpc2932 (
      {stage1_8[185]},
      {stage2_8[87]}
   );
   gpc1_1 gpc2933 (
      {stage1_8[186]},
      {stage2_8[88]}
   );
   gpc1_1 gpc2934 (
      {stage1_8[187]},
      {stage2_8[89]}
   );
   gpc1_1 gpc2935 (
      {stage1_8[188]},
      {stage2_8[90]}
   );
   gpc1_1 gpc2936 (
      {stage1_8[189]},
      {stage2_8[91]}
   );
   gpc1_1 gpc2937 (
      {stage1_8[190]},
      {stage2_8[92]}
   );
   gpc1_1 gpc2938 (
      {stage1_8[191]},
      {stage2_8[93]}
   );
   gpc1_1 gpc2939 (
      {stage1_8[192]},
      {stage2_8[94]}
   );
   gpc1_1 gpc2940 (
      {stage1_8[193]},
      {stage2_8[95]}
   );
   gpc1_1 gpc2941 (
      {stage1_8[194]},
      {stage2_8[96]}
   );
   gpc1_1 gpc2942 (
      {stage1_8[195]},
      {stage2_8[97]}
   );
   gpc1_1 gpc2943 (
      {stage1_8[196]},
      {stage2_8[98]}
   );
   gpc1_1 gpc2944 (
      {stage1_8[197]},
      {stage2_8[99]}
   );
   gpc1_1 gpc2945 (
      {stage1_8[198]},
      {stage2_8[100]}
   );
   gpc1_1 gpc2946 (
      {stage1_8[199]},
      {stage2_8[101]}
   );
   gpc1_1 gpc2947 (
      {stage1_8[200]},
      {stage2_8[102]}
   );
   gpc1_1 gpc2948 (
      {stage1_8[201]},
      {stage2_8[103]}
   );
   gpc1_1 gpc2949 (
      {stage1_8[202]},
      {stage2_8[104]}
   );
   gpc1_1 gpc2950 (
      {stage1_8[203]},
      {stage2_8[105]}
   );
   gpc1_1 gpc2951 (
      {stage1_8[204]},
      {stage2_8[106]}
   );
   gpc1_1 gpc2952 (
      {stage1_8[205]},
      {stage2_8[107]}
   );
   gpc1_1 gpc2953 (
      {stage1_9[211]},
      {stage2_9[72]}
   );
   gpc1_1 gpc2954 (
      {stage1_9[212]},
      {stage2_9[73]}
   );
   gpc1_1 gpc2955 (
      {stage1_9[213]},
      {stage2_9[74]}
   );
   gpc1_1 gpc2956 (
      {stage1_10[186]},
      {stage2_10[87]}
   );
   gpc1_1 gpc2957 (
      {stage1_10[187]},
      {stage2_10[88]}
   );
   gpc1_1 gpc2958 (
      {stage1_12[277]},
      {stage2_12[98]}
   );
   gpc1_1 gpc2959 (
      {stage1_12[278]},
      {stage2_12[99]}
   );
   gpc1_1 gpc2960 (
      {stage1_12[279]},
      {stage2_12[100]}
   );
   gpc1_1 gpc2961 (
      {stage1_12[280]},
      {stage2_12[101]}
   );
   gpc1_1 gpc2962 (
      {stage1_12[281]},
      {stage2_12[102]}
   );
   gpc1_1 gpc2963 (
      {stage1_14[238]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2964 (
      {stage1_14[239]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2965 (
      {stage1_14[240]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2966 (
      {stage1_14[241]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2967 (
      {stage1_14[242]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2968 (
      {stage1_14[243]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2969 (
      {stage1_14[244]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2970 (
      {stage1_14[245]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2971 (
      {stage1_14[246]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2972 (
      {stage1_14[247]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2973 (
      {stage1_14[248]},
      {stage2_14[90]}
   );
   gpc1_1 gpc2974 (
      {stage1_14[249]},
      {stage2_14[91]}
   );
   gpc1_1 gpc2975 (
      {stage1_14[250]},
      {stage2_14[92]}
   );
   gpc1_1 gpc2976 (
      {stage1_14[251]},
      {stage2_14[93]}
   );
   gpc1_1 gpc2977 (
      {stage1_14[252]},
      {stage2_14[94]}
   );
   gpc1_1 gpc2978 (
      {stage1_14[253]},
      {stage2_14[95]}
   );
   gpc1_1 gpc2979 (
      {stage1_14[254]},
      {stage2_14[96]}
   );
   gpc1_1 gpc2980 (
      {stage1_14[255]},
      {stage2_14[97]}
   );
   gpc1_1 gpc2981 (
      {stage1_14[256]},
      {stage2_14[98]}
   );
   gpc1_1 gpc2982 (
      {stage1_14[257]},
      {stage2_14[99]}
   );
   gpc1_1 gpc2983 (
      {stage1_14[258]},
      {stage2_14[100]}
   );
   gpc1_1 gpc2984 (
      {stage1_14[259]},
      {stage2_14[101]}
   );
   gpc1_1 gpc2985 (
      {stage1_14[260]},
      {stage2_14[102]}
   );
   gpc1_1 gpc2986 (
      {stage1_14[261]},
      {stage2_14[103]}
   );
   gpc1_1 gpc2987 (
      {stage1_14[262]},
      {stage2_14[104]}
   );
   gpc1_1 gpc2988 (
      {stage1_14[263]},
      {stage2_14[105]}
   );
   gpc1_1 gpc2989 (
      {stage1_14[264]},
      {stage2_14[106]}
   );
   gpc1_1 gpc2990 (
      {stage1_14[265]},
      {stage2_14[107]}
   );
   gpc1_1 gpc2991 (
      {stage1_14[266]},
      {stage2_14[108]}
   );
   gpc1_1 gpc2992 (
      {stage1_14[267]},
      {stage2_14[109]}
   );
   gpc1_1 gpc2993 (
      {stage1_14[268]},
      {stage2_14[110]}
   );
   gpc1_1 gpc2994 (
      {stage1_14[269]},
      {stage2_14[111]}
   );
   gpc1_1 gpc2995 (
      {stage1_14[270]},
      {stage2_14[112]}
   );
   gpc1_1 gpc2996 (
      {stage1_14[271]},
      {stage2_14[113]}
   );
   gpc1_1 gpc2997 (
      {stage1_14[272]},
      {stage2_14[114]}
   );
   gpc1_1 gpc2998 (
      {stage1_14[273]},
      {stage2_14[115]}
   );
   gpc1_1 gpc2999 (
      {stage1_14[274]},
      {stage2_14[116]}
   );
   gpc1_1 gpc3000 (
      {stage1_14[275]},
      {stage2_14[117]}
   );
   gpc1_1 gpc3001 (
      {stage1_14[276]},
      {stage2_14[118]}
   );
   gpc1_1 gpc3002 (
      {stage1_14[277]},
      {stage2_14[119]}
   );
   gpc1_1 gpc3003 (
      {stage1_14[278]},
      {stage2_14[120]}
   );
   gpc1_1 gpc3004 (
      {stage1_14[279]},
      {stage2_14[121]}
   );
   gpc1_1 gpc3005 (
      {stage1_14[280]},
      {stage2_14[122]}
   );
   gpc1_1 gpc3006 (
      {stage1_14[281]},
      {stage2_14[123]}
   );
   gpc1_1 gpc3007 (
      {stage1_14[282]},
      {stage2_14[124]}
   );
   gpc1_1 gpc3008 (
      {stage1_14[283]},
      {stage2_14[125]}
   );
   gpc1_1 gpc3009 (
      {stage1_14[284]},
      {stage2_14[126]}
   );
   gpc1_1 gpc3010 (
      {stage1_14[285]},
      {stage2_14[127]}
   );
   gpc1_1 gpc3011 (
      {stage1_14[286]},
      {stage2_14[128]}
   );
   gpc1_1 gpc3012 (
      {stage1_14[287]},
      {stage2_14[129]}
   );
   gpc1_1 gpc3013 (
      {stage1_14[288]},
      {stage2_14[130]}
   );
   gpc1_1 gpc3014 (
      {stage1_14[289]},
      {stage2_14[131]}
   );
   gpc1_1 gpc3015 (
      {stage1_14[290]},
      {stage2_14[132]}
   );
   gpc1_1 gpc3016 (
      {stage1_14[291]},
      {stage2_14[133]}
   );
   gpc1_1 gpc3017 (
      {stage1_14[292]},
      {stage2_14[134]}
   );
   gpc1_1 gpc3018 (
      {stage1_14[293]},
      {stage2_14[135]}
   );
   gpc1_1 gpc3019 (
      {stage1_14[294]},
      {stage2_14[136]}
   );
   gpc1_1 gpc3020 (
      {stage1_14[295]},
      {stage2_14[137]}
   );
   gpc1_1 gpc3021 (
      {stage1_14[296]},
      {stage2_14[138]}
   );
   gpc1_1 gpc3022 (
      {stage1_15[128]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3023 (
      {stage1_15[129]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3024 (
      {stage1_15[130]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3025 (
      {stage1_15[131]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3026 (
      {stage1_15[132]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3027 (
      {stage1_15[133]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3028 (
      {stage1_15[134]},
      {stage2_15[98]}
   );
   gpc1_1 gpc3029 (
      {stage1_15[135]},
      {stage2_15[99]}
   );
   gpc1_1 gpc3030 (
      {stage1_15[136]},
      {stage2_15[100]}
   );
   gpc1_1 gpc3031 (
      {stage1_15[137]},
      {stage2_15[101]}
   );
   gpc1_1 gpc3032 (
      {stage1_15[138]},
      {stage2_15[102]}
   );
   gpc1_1 gpc3033 (
      {stage1_15[139]},
      {stage2_15[103]}
   );
   gpc1_1 gpc3034 (
      {stage1_15[140]},
      {stage2_15[104]}
   );
   gpc1_1 gpc3035 (
      {stage1_15[141]},
      {stage2_15[105]}
   );
   gpc1_1 gpc3036 (
      {stage1_15[142]},
      {stage2_15[106]}
   );
   gpc1_1 gpc3037 (
      {stage1_15[143]},
      {stage2_15[107]}
   );
   gpc1_1 gpc3038 (
      {stage1_15[144]},
      {stage2_15[108]}
   );
   gpc1_1 gpc3039 (
      {stage1_15[145]},
      {stage2_15[109]}
   );
   gpc1_1 gpc3040 (
      {stage1_15[146]},
      {stage2_15[110]}
   );
   gpc1_1 gpc3041 (
      {stage1_15[147]},
      {stage2_15[111]}
   );
   gpc1_1 gpc3042 (
      {stage1_15[148]},
      {stage2_15[112]}
   );
   gpc1_1 gpc3043 (
      {stage1_15[149]},
      {stage2_15[113]}
   );
   gpc1_1 gpc3044 (
      {stage1_15[150]},
      {stage2_15[114]}
   );
   gpc1_1 gpc3045 (
      {stage1_15[151]},
      {stage2_15[115]}
   );
   gpc1_1 gpc3046 (
      {stage1_15[152]},
      {stage2_15[116]}
   );
   gpc1_1 gpc3047 (
      {stage1_15[153]},
      {stage2_15[117]}
   );
   gpc1_1 gpc3048 (
      {stage1_15[154]},
      {stage2_15[118]}
   );
   gpc1_1 gpc3049 (
      {stage1_15[155]},
      {stage2_15[119]}
   );
   gpc1_1 gpc3050 (
      {stage1_15[156]},
      {stage2_15[120]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[157]},
      {stage2_15[121]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[158]},
      {stage2_15[122]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[159]},
      {stage2_15[123]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[160]},
      {stage2_15[124]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[161]},
      {stage2_15[125]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[162]},
      {stage2_15[126]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[163]},
      {stage2_15[127]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[164]},
      {stage2_15[128]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[165]},
      {stage2_15[129]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[166]},
      {stage2_15[130]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[167]},
      {stage2_15[131]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[168]},
      {stage2_15[132]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[169]},
      {stage2_15[133]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[170]},
      {stage2_15[134]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[171]},
      {stage2_15[135]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[257]},
      {stage2_16[96]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[258]},
      {stage2_16[97]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[259]},
      {stage2_16[98]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[260]},
      {stage2_16[99]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[261]},
      {stage2_16[100]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[262]},
      {stage2_16[101]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[263]},
      {stage2_16[102]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[264]},
      {stage2_16[103]}
   );
   gpc1_1 gpc3074 (
      {stage1_17[234]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3075 (
      {stage1_17[235]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3076 (
      {stage1_17[236]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3077 (
      {stage1_17[237]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3078 (
      {stage1_17[238]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3079 (
      {stage1_17[239]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3080 (
      {stage1_17[240]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3081 (
      {stage1_17[241]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3082 (
      {stage1_17[242]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3083 (
      {stage1_17[243]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[244]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[245]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[246]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[247]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[248]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[249]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[250]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[251]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[252]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[253]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[254]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[255]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[256]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[257]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[258]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[259]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[260]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[261]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[262]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[263]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[264]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[265]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[266]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[267]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[268]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[269]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[270]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3111 (
      {stage1_18[198]},
      {stage2_18[79]}
   );
   gpc1_1 gpc3112 (
      {stage1_18[199]},
      {stage2_18[80]}
   );
   gpc1_1 gpc3113 (
      {stage1_18[200]},
      {stage2_18[81]}
   );
   gpc1_1 gpc3114 (
      {stage1_19[295]},
      {stage2_19[105]}
   );
   gpc1_1 gpc3115 (
      {stage1_19[296]},
      {stage2_19[106]}
   );
   gpc1_1 gpc3116 (
      {stage1_19[297]},
      {stage2_19[107]}
   );
   gpc1_1 gpc3117 (
      {stage1_19[298]},
      {stage2_19[108]}
   );
   gpc1_1 gpc3118 (
      {stage1_19[299]},
      {stage2_19[109]}
   );
   gpc1_1 gpc3119 (
      {stage1_20[172]},
      {stage2_20[111]}
   );
   gpc1_1 gpc3120 (
      {stage1_20[173]},
      {stage2_20[112]}
   );
   gpc1_1 gpc3121 (
      {stage1_20[174]},
      {stage2_20[113]}
   );
   gpc1_1 gpc3122 (
      {stage1_20[175]},
      {stage2_20[114]}
   );
   gpc1_1 gpc3123 (
      {stage1_20[176]},
      {stage2_20[115]}
   );
   gpc1_1 gpc3124 (
      {stage1_20[177]},
      {stage2_20[116]}
   );
   gpc1_1 gpc3125 (
      {stage1_20[178]},
      {stage2_20[117]}
   );
   gpc1_1 gpc3126 (
      {stage1_20[179]},
      {stage2_20[118]}
   );
   gpc1_1 gpc3127 (
      {stage1_20[180]},
      {stage2_20[119]}
   );
   gpc1_1 gpc3128 (
      {stage1_20[181]},
      {stage2_20[120]}
   );
   gpc1_1 gpc3129 (
      {stage1_20[182]},
      {stage2_20[121]}
   );
   gpc1_1 gpc3130 (
      {stage1_20[183]},
      {stage2_20[122]}
   );
   gpc1_1 gpc3131 (
      {stage1_20[184]},
      {stage2_20[123]}
   );
   gpc1_1 gpc3132 (
      {stage1_20[185]},
      {stage2_20[124]}
   );
   gpc1_1 gpc3133 (
      {stage1_20[186]},
      {stage2_20[125]}
   );
   gpc1_1 gpc3134 (
      {stage1_20[187]},
      {stage2_20[126]}
   );
   gpc1_1 gpc3135 (
      {stage1_20[188]},
      {stage2_20[127]}
   );
   gpc1_1 gpc3136 (
      {stage1_21[198]},
      {stage2_21[78]}
   );
   gpc1_1 gpc3137 (
      {stage1_24[194]},
      {stage2_24[82]}
   );
   gpc1_1 gpc3138 (
      {stage1_24[195]},
      {stage2_24[83]}
   );
   gpc1_1 gpc3139 (
      {stage1_24[196]},
      {stage2_24[84]}
   );
   gpc1_1 gpc3140 (
      {stage1_24[197]},
      {stage2_24[85]}
   );
   gpc1_1 gpc3141 (
      {stage1_24[198]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3142 (
      {stage1_24[199]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3143 (
      {stage1_24[200]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3144 (
      {stage1_24[201]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3145 (
      {stage1_24[202]},
      {stage2_24[90]}
   );
   gpc1_1 gpc3146 (
      {stage1_24[203]},
      {stage2_24[91]}
   );
   gpc1_1 gpc3147 (
      {stage1_24[204]},
      {stage2_24[92]}
   );
   gpc1_1 gpc3148 (
      {stage1_24[205]},
      {stage2_24[93]}
   );
   gpc1_1 gpc3149 (
      {stage1_24[206]},
      {stage2_24[94]}
   );
   gpc1_1 gpc3150 (
      {stage1_24[207]},
      {stage2_24[95]}
   );
   gpc1_1 gpc3151 (
      {stage1_24[208]},
      {stage2_24[96]}
   );
   gpc1_1 gpc3152 (
      {stage1_24[209]},
      {stage2_24[97]}
   );
   gpc1_1 gpc3153 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc3154 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc3155 (
      {stage1_25[209]},
      {stage2_25[62]}
   );
   gpc1_1 gpc3156 (
      {stage1_25[210]},
      {stage2_25[63]}
   );
   gpc1_1 gpc3157 (
      {stage1_25[211]},
      {stage2_25[64]}
   );
   gpc1_1 gpc3158 (
      {stage1_25[212]},
      {stage2_25[65]}
   );
   gpc1_1 gpc3159 (
      {stage1_25[213]},
      {stage2_25[66]}
   );
   gpc1_1 gpc3160 (
      {stage1_25[214]},
      {stage2_25[67]}
   );
   gpc1_1 gpc3161 (
      {stage1_25[215]},
      {stage2_25[68]}
   );
   gpc1_1 gpc3162 (
      {stage1_25[216]},
      {stage2_25[69]}
   );
   gpc1_1 gpc3163 (
      {stage1_25[217]},
      {stage2_25[70]}
   );
   gpc1_1 gpc3164 (
      {stage1_25[218]},
      {stage2_25[71]}
   );
   gpc1_1 gpc3165 (
      {stage1_25[219]},
      {stage2_25[72]}
   );
   gpc1_1 gpc3166 (
      {stage1_25[220]},
      {stage2_25[73]}
   );
   gpc1_1 gpc3167 (
      {stage1_25[221]},
      {stage2_25[74]}
   );
   gpc1_1 gpc3168 (
      {stage1_25[222]},
      {stage2_25[75]}
   );
   gpc1_1 gpc3169 (
      {stage1_25[223]},
      {stage2_25[76]}
   );
   gpc1_1 gpc3170 (
      {stage1_25[224]},
      {stage2_25[77]}
   );
   gpc1_1 gpc3171 (
      {stage1_25[225]},
      {stage2_25[78]}
   );
   gpc1_1 gpc3172 (
      {stage1_25[226]},
      {stage2_25[79]}
   );
   gpc1_1 gpc3173 (
      {stage1_25[227]},
      {stage2_25[80]}
   );
   gpc1_1 gpc3174 (
      {stage1_25[228]},
      {stage2_25[81]}
   );
   gpc1_1 gpc3175 (
      {stage1_25[229]},
      {stage2_25[82]}
   );
   gpc1_1 gpc3176 (
      {stage1_25[230]},
      {stage2_25[83]}
   );
   gpc1_1 gpc3177 (
      {stage1_25[231]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3178 (
      {stage1_25[232]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3179 (
      {stage1_25[233]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3180 (
      {stage1_25[234]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3181 (
      {stage1_28[243]},
      {stage2_28[66]}
   );
   gpc1_1 gpc3182 (
      {stage1_28[244]},
      {stage2_28[67]}
   );
   gpc1_1 gpc3183 (
      {stage1_28[245]},
      {stage2_28[68]}
   );
   gpc1_1 gpc3184 (
      {stage1_28[246]},
      {stage2_28[69]}
   );
   gpc1_1 gpc3185 (
      {stage1_28[247]},
      {stage2_28[70]}
   );
   gpc1_1 gpc3186 (
      {stage1_28[248]},
      {stage2_28[71]}
   );
   gpc1_1 gpc3187 (
      {stage1_28[249]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3188 (
      {stage1_28[250]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3189 (
      {stage1_28[251]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3190 (
      {stage1_29[186]},
      {stage2_29[71]}
   );
   gpc1_1 gpc3191 (
      {stage1_29[187]},
      {stage2_29[72]}
   );
   gpc1_1 gpc3192 (
      {stage1_29[188]},
      {stage2_29[73]}
   );
   gpc1_1 gpc3193 (
      {stage1_29[189]},
      {stage2_29[74]}
   );
   gpc1_1 gpc3194 (
      {stage1_29[190]},
      {stage2_29[75]}
   );
   gpc1_1 gpc3195 (
      {stage1_29[191]},
      {stage2_29[76]}
   );
   gpc1_1 gpc3196 (
      {stage1_29[192]},
      {stage2_29[77]}
   );
   gpc1_1 gpc3197 (
      {stage1_29[193]},
      {stage2_29[78]}
   );
   gpc1_1 gpc3198 (
      {stage1_29[194]},
      {stage2_29[79]}
   );
   gpc1_1 gpc3199 (
      {stage1_29[195]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3200 (
      {stage1_29[196]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3201 (
      {stage1_29[197]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3202 (
      {stage1_29[198]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3203 (
      {stage1_29[199]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3204 (
      {stage1_29[200]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3205 (
      {stage1_29[201]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3206 (
      {stage1_29[202]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3207 (
      {stage1_29[203]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3208 (
      {stage1_29[204]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3209 (
      {stage1_29[205]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3210 (
      {stage1_29[206]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3211 (
      {stage1_29[207]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3212 (
      {stage1_29[208]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3213 (
      {stage1_29[209]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3214 (
      {stage1_29[210]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3215 (
      {stage1_29[211]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3216 (
      {stage1_29[212]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3217 (
      {stage1_29[213]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3218 (
      {stage1_29[214]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3219 (
      {stage1_29[215]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3220 (
      {stage1_29[216]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3221 (
      {stage1_29[217]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3222 (
      {stage1_29[218]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3223 (
      {stage1_29[219]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3224 (
      {stage1_29[220]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3225 (
      {stage1_29[221]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3226 (
      {stage1_29[222]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3227 (
      {stage1_29[223]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3228 (
      {stage1_29[224]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3229 (
      {stage1_29[225]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3230 (
      {stage1_29[226]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3231 (
      {stage1_29[227]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3232 (
      {stage1_29[228]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3233 (
      {stage1_29[229]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3234 (
      {stage1_29[230]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3235 (
      {stage1_29[231]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3236 (
      {stage1_29[232]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3237 (
      {stage1_29[233]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3238 (
      {stage1_29[234]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3239 (
      {stage1_29[235]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3240 (
      {stage1_30[132]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3241 (
      {stage1_30[133]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3242 (
      {stage1_30[134]},
      {stage2_30[92]}
   );
   gpc1_1 gpc3243 (
      {stage1_30[135]},
      {stage2_30[93]}
   );
   gpc1_1 gpc3244 (
      {stage1_30[136]},
      {stage2_30[94]}
   );
   gpc1_1 gpc3245 (
      {stage1_30[137]},
      {stage2_30[95]}
   );
   gpc1_1 gpc3246 (
      {stage1_30[138]},
      {stage2_30[96]}
   );
   gpc1_1 gpc3247 (
      {stage1_30[139]},
      {stage2_30[97]}
   );
   gpc1_1 gpc3248 (
      {stage1_30[140]},
      {stage2_30[98]}
   );
   gpc1_1 gpc3249 (
      {stage1_30[141]},
      {stage2_30[99]}
   );
   gpc1_1 gpc3250 (
      {stage1_30[142]},
      {stage2_30[100]}
   );
   gpc1_1 gpc3251 (
      {stage1_30[143]},
      {stage2_30[101]}
   );
   gpc1_1 gpc3252 (
      {stage1_30[144]},
      {stage2_30[102]}
   );
   gpc1_1 gpc3253 (
      {stage1_30[145]},
      {stage2_30[103]}
   );
   gpc1_1 gpc3254 (
      {stage1_30[146]},
      {stage2_30[104]}
   );
   gpc1_1 gpc3255 (
      {stage1_30[147]},
      {stage2_30[105]}
   );
   gpc1_1 gpc3256 (
      {stage1_30[148]},
      {stage2_30[106]}
   );
   gpc1_1 gpc3257 (
      {stage1_30[149]},
      {stage2_30[107]}
   );
   gpc1_1 gpc3258 (
      {stage1_30[150]},
      {stage2_30[108]}
   );
   gpc1_1 gpc3259 (
      {stage1_30[151]},
      {stage2_30[109]}
   );
   gpc1_1 gpc3260 (
      {stage1_30[152]},
      {stage2_30[110]}
   );
   gpc1_1 gpc3261 (
      {stage1_30[153]},
      {stage2_30[111]}
   );
   gpc1_1 gpc3262 (
      {stage1_30[154]},
      {stage2_30[112]}
   );
   gpc1_1 gpc3263 (
      {stage1_30[155]},
      {stage2_30[113]}
   );
   gpc1_1 gpc3264 (
      {stage1_30[156]},
      {stage2_30[114]}
   );
   gpc1_1 gpc3265 (
      {stage1_30[157]},
      {stage2_30[115]}
   );
   gpc1_1 gpc3266 (
      {stage1_30[158]},
      {stage2_30[116]}
   );
   gpc1_1 gpc3267 (
      {stage1_30[159]},
      {stage2_30[117]}
   );
   gpc1_1 gpc3268 (
      {stage1_30[160]},
      {stage2_30[118]}
   );
   gpc1_1 gpc3269 (
      {stage1_30[161]},
      {stage2_30[119]}
   );
   gpc1_1 gpc3270 (
      {stage1_30[162]},
      {stage2_30[120]}
   );
   gpc1_1 gpc3271 (
      {stage1_30[163]},
      {stage2_30[121]}
   );
   gpc1_1 gpc3272 (
      {stage1_30[164]},
      {stage2_30[122]}
   );
   gpc1_1 gpc3273 (
      {stage1_30[165]},
      {stage2_30[123]}
   );
   gpc1_1 gpc3274 (
      {stage1_30[166]},
      {stage2_30[124]}
   );
   gpc1_1 gpc3275 (
      {stage1_30[167]},
      {stage2_30[125]}
   );
   gpc1_1 gpc3276 (
      {stage1_30[168]},
      {stage2_30[126]}
   );
   gpc1_1 gpc3277 (
      {stage1_30[169]},
      {stage2_30[127]}
   );
   gpc1_1 gpc3278 (
      {stage1_30[170]},
      {stage2_30[128]}
   );
   gpc1_1 gpc3279 (
      {stage1_30[171]},
      {stage2_30[129]}
   );
   gpc1_1 gpc3280 (
      {stage1_31[144]},
      {stage2_31[67]}
   );
   gpc1_1 gpc3281 (
      {stage1_31[145]},
      {stage2_31[68]}
   );
   gpc1_1 gpc3282 (
      {stage1_31[146]},
      {stage2_31[69]}
   );
   gpc1_1 gpc3283 (
      {stage1_31[147]},
      {stage2_31[70]}
   );
   gpc1_1 gpc3284 (
      {stage1_31[148]},
      {stage2_31[71]}
   );
   gpc1_1 gpc3285 (
      {stage1_31[149]},
      {stage2_31[72]}
   );
   gpc1_1 gpc3286 (
      {stage1_31[150]},
      {stage2_31[73]}
   );
   gpc1_1 gpc3287 (
      {stage1_31[151]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3288 (
      {stage1_31[152]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3289 (
      {stage1_31[153]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3290 (
      {stage1_31[154]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3291 (
      {stage1_31[155]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3292 (
      {stage1_31[156]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3293 (
      {stage1_31[157]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3294 (
      {stage1_31[158]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3295 (
      {stage1_31[159]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3296 (
      {stage1_31[160]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3297 (
      {stage1_32[132]},
      {stage2_32[46]}
   );
   gpc1_1 gpc3298 (
      {stage1_32[133]},
      {stage2_32[47]}
   );
   gpc1_1 gpc3299 (
      {stage1_32[134]},
      {stage2_32[48]}
   );
   gpc1_1 gpc3300 (
      {stage1_32[135]},
      {stage2_32[49]}
   );
   gpc1_1 gpc3301 (
      {stage1_32[136]},
      {stage2_32[50]}
   );
   gpc1_1 gpc3302 (
      {stage1_32[137]},
      {stage2_32[51]}
   );
   gpc1_1 gpc3303 (
      {stage1_32[138]},
      {stage2_32[52]}
   );
   gpc1_1 gpc3304 (
      {stage1_32[139]},
      {stage2_32[53]}
   );
   gpc1_1 gpc3305 (
      {stage1_32[140]},
      {stage2_32[54]}
   );
   gpc1_1 gpc3306 (
      {stage1_32[141]},
      {stage2_32[55]}
   );
   gpc1_1 gpc3307 (
      {stage1_32[142]},
      {stage2_32[56]}
   );
   gpc1_1 gpc3308 (
      {stage1_32[143]},
      {stage2_32[57]}
   );
   gpc1_1 gpc3309 (
      {stage1_32[144]},
      {stage2_32[58]}
   );
   gpc1_1 gpc3310 (
      {stage1_32[145]},
      {stage2_32[59]}
   );
   gpc1_1 gpc3311 (
      {stage1_32[146]},
      {stage2_32[60]}
   );
   gpc1_1 gpc3312 (
      {stage1_32[147]},
      {stage2_32[61]}
   );
   gpc1_1 gpc3313 (
      {stage1_32[148]},
      {stage2_32[62]}
   );
   gpc1_1 gpc3314 (
      {stage1_32[149]},
      {stage2_32[63]}
   );
   gpc1_1 gpc3315 (
      {stage1_32[150]},
      {stage2_32[64]}
   );
   gpc1163_5 gpc3316 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc3317 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc3318 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc3319 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc1163_5 gpc3320 (
      {stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_2[4]},
      {stage2_3[4]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc1163_5 gpc3321 (
      {stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_2[5]},
      {stage2_3[5]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1163_5 gpc3322 (
      {stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[6]},
      {stage2_3[6]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3323 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[0],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc3324 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[1],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc3325 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[2],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc3326 (
      {stage2_1[60], stage2_1[61], stage2_1[62], stage2_1[63], stage2_1[64], stage2_1[65]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[3],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc3327 (
      {stage2_1[66], stage2_1[67], stage2_1[68], stage2_1[69], stage2_1[70], stage2_1[71]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[4],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3328 (
      {stage2_1[72], stage2_1[73], stage2_1[74], stage2_1[75], stage2_1[76], stage2_1[77]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[5],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3329 (
      {stage2_1[78], stage2_1[79], stage2_1[80], stage2_1[81], stage2_1[82], stage2_1[83]},
      {stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage3_5[6],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3330 (
      {stage2_1[84], stage2_1[85], stage2_1[86], stage2_1[87], stage2_1[88], stage2_1[89]},
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage3_5[7],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3331 (
      {stage2_1[90], stage2_1[91], stage2_1[92], stage2_1[93], stage2_1[94], stage2_1[95]},
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60]},
      {stage3_5[8],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3332 (
      {stage2_1[96], stage2_1[97], stage2_1[98], stage2_1[99], stage2_1[100], stage2_1[101]},
      {stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage3_5[9],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3333 (
      {stage2_1[102], stage2_1[103], stage2_1[104], stage2_1[105], stage2_1[106], 1'b0},
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage3_5[10],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc606_5 gpc3334 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[11],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc606_5 gpc3335 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[12],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc606_5 gpc3336 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[13],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc606_5 gpc3337 (
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[14],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc606_5 gpc3338 (
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[15],stage3_4[22],stage3_3[22],stage3_2[22]}
   );
   gpc606_5 gpc3339 (
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[16],stage3_4[23],stage3_3[23],stage3_2[23]}
   );
   gpc615_5 gpc3340 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[17],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3341 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[18],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3342 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[19],stage3_4[26],stage3_3[26]}
   );
   gpc606_5 gpc3343 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[20],stage3_4[27]}
   );
   gpc606_5 gpc3344 (
      {stage2_4[45], stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[21],stage3_4[28]}
   );
   gpc606_5 gpc3345 (
      {stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[22],stage3_4[29]}
   );
   gpc615_5 gpc3346 (
      {stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[12],stage3_5[23],stage3_4[30]}
   );
   gpc615_5 gpc3347 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[13],stage3_5[24],stage3_4[31]}
   );
   gpc615_5 gpc3348 (
      {stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[14],stage3_5[25],stage3_4[32]}
   );
   gpc615_5 gpc3349 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[15],stage3_5[26],stage3_4[33]}
   );
   gpc615_5 gpc3350 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[16],stage3_5[27],stage3_4[34]}
   );
   gpc606_5 gpc3351 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[17],stage3_5[28]}
   );
   gpc606_5 gpc3352 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[18],stage3_5[29]}
   );
   gpc606_5 gpc3353 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[19],stage3_5[30]}
   );
   gpc606_5 gpc3354 (
      {stage2_5[41], stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[11],stage3_7[14],stage3_6[20],stage3_5[31]}
   );
   gpc606_5 gpc3355 (
      {stage2_5[47], stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[12],stage3_7[15],stage3_6[21],stage3_5[32]}
   );
   gpc606_5 gpc3356 (
      {stage2_5[53], stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[13],stage3_7[16],stage3_6[22],stage3_5[33]}
   );
   gpc606_5 gpc3357 (
      {stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[14],stage3_7[17],stage3_6[23],stage3_5[34]}
   );
   gpc606_5 gpc3358 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[15],stage3_7[18],stage3_6[24],stage3_5[35]}
   );
   gpc615_5 gpc3359 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[48]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[8],stage3_8[16],stage3_7[19],stage3_6[25]}
   );
   gpc615_5 gpc3360 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[49]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[9],stage3_8[17],stage3_7[20],stage3_6[26]}
   );
   gpc615_5 gpc3361 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[50]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[10],stage3_8[18],stage3_7[21],stage3_6[27]}
   );
   gpc615_5 gpc3362 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[51]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[11],stage3_8[19],stage3_7[22],stage3_6[28]}
   );
   gpc615_5 gpc3363 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[52]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[12],stage3_8[20],stage3_7[23],stage3_6[29]}
   );
   gpc615_5 gpc3364 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[53]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[13],stage3_8[21],stage3_7[24],stage3_6[30]}
   );
   gpc615_5 gpc3365 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[54]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[14],stage3_8[22],stage3_7[25],stage3_6[31]}
   );
   gpc615_5 gpc3366 (
      {stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage2_8[42]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[7],stage3_9[15],stage3_8[23],stage3_7[26]}
   );
   gpc615_5 gpc3367 (
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64]},
      {stage2_8[43]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[8],stage3_9[16],stage3_8[24],stage3_7[27]}
   );
   gpc615_5 gpc3368 (
      {stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69]},
      {stage2_8[44]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[9],stage3_9[17],stage3_8[25],stage3_7[28]}
   );
   gpc1343_5 gpc3369 (
      {stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[3],stage3_10[10],stage3_9[18],stage3_8[26]}
   );
   gpc1343_5 gpc3370 (
      {stage2_8[48], stage2_8[49], stage2_8[50]},
      {stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25]},
      {stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_11[1]},
      {stage3_12[1],stage3_11[4],stage3_10[11],stage3_9[19],stage3_8[27]}
   );
   gpc1343_5 gpc3371 (
      {stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_10[6], stage2_10[7], stage2_10[8]},
      {stage2_11[2]},
      {stage3_12[2],stage3_11[5],stage3_10[12],stage3_9[20],stage3_8[28]}
   );
   gpc606_5 gpc3372 (
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13], stage2_10[14]},
      {stage3_12[3],stage3_11[6],stage3_10[13],stage3_9[21],stage3_8[29]}
   );
   gpc606_5 gpc3373 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage3_12[4],stage3_11[7],stage3_10[14],stage3_9[22],stage3_8[30]}
   );
   gpc606_5 gpc3374 (
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25], stage2_10[26]},
      {stage3_12[5],stage3_11[8],stage3_10[15],stage3_9[23],stage3_8[31]}
   );
   gpc606_5 gpc3375 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31], stage2_10[32]},
      {stage3_12[6],stage3_11[9],stage3_10[16],stage3_9[24],stage3_8[32]}
   );
   gpc606_5 gpc3376 (
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage3_12[7],stage3_11[10],stage3_10[17],stage3_9[25],stage3_8[33]}
   );
   gpc606_5 gpc3377 (
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage3_12[8],stage3_11[11],stage3_10[18],stage3_9[26],stage3_8[34]}
   );
   gpc606_5 gpc3378 (
      {stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94], stage2_8[95]},
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage3_12[9],stage3_11[12],stage3_10[19],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc3379 (
      {stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100], stage2_8[101]},
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage3_12[10],stage3_11[13],stage3_10[20],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc3380 (
      {stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106], stage2_8[107]},
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage3_12[11],stage3_11[14],stage3_10[21],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc3381 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage3_13[0],stage3_12[12],stage3_11[15],stage3_10[22],stage3_9[30]}
   );
   gpc615_5 gpc3382 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67]},
      {stage2_11[9]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[13],stage3_11[16],stage3_10[23]}
   );
   gpc615_5 gpc3383 (
      {stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72]},
      {stage2_11[10]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[14],stage3_11[17],stage3_10[24]}
   );
   gpc615_5 gpc3384 (
      {stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage2_11[11]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[15],stage3_11[18],stage3_10[25]}
   );
   gpc615_5 gpc3385 (
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82]},
      {stage2_11[12]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[16],stage3_11[19],stage3_10[26]}
   );
   gpc615_5 gpc3386 (
      {stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87]},
      {stage2_11[13]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[17],stage3_11[20],stage3_10[27]}
   );
   gpc606_5 gpc3387 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[5],stage3_13[6],stage3_12[18],stage3_11[21]}
   );
   gpc606_5 gpc3388 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[6],stage3_13[7],stage3_12[19],stage3_11[22]}
   );
   gpc606_5 gpc3389 (
      {stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[7],stage3_13[8],stage3_12[20],stage3_11[23]}
   );
   gpc606_5 gpc3390 (
      {stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[8],stage3_13[9],stage3_12[21],stage3_11[24]}
   );
   gpc606_5 gpc3391 (
      {stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[9],stage3_13[10],stage3_12[22],stage3_11[25]}
   );
   gpc606_5 gpc3392 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[10],stage3_13[11],stage3_12[23],stage3_11[26]}
   );
   gpc606_5 gpc3393 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[11],stage3_13[12],stage3_12[24],stage3_11[27]}
   );
   gpc606_5 gpc3394 (
      {stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[12],stage3_13[13],stage3_12[25],stage3_11[28]}
   );
   gpc606_5 gpc3395 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[13],stage3_13[14],stage3_12[26],stage3_11[29]}
   );
   gpc606_5 gpc3396 (
      {stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[14],stage3_13[15],stage3_12[27],stage3_11[30]}
   );
   gpc606_5 gpc3397 (
      {stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[15],stage3_13[16],stage3_12[28],stage3_11[31]}
   );
   gpc606_5 gpc3398 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[11],stage3_14[16],stage3_13[17],stage3_12[29]}
   );
   gpc606_5 gpc3399 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[12],stage3_14[17],stage3_13[18],stage3_12[30]}
   );
   gpc606_5 gpc3400 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[13],stage3_14[18],stage3_13[19],stage3_12[31]}
   );
   gpc606_5 gpc3401 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[14],stage3_14[19],stage3_13[20],stage3_12[32]}
   );
   gpc606_5 gpc3402 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[15],stage3_14[20],stage3_13[21],stage3_12[33]}
   );
   gpc606_5 gpc3403 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[16],stage3_14[21],stage3_13[22],stage3_12[34]}
   );
   gpc606_5 gpc3404 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[17],stage3_14[22],stage3_13[23],stage3_12[35]}
   );
   gpc606_5 gpc3405 (
      {stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[18],stage3_14[23],stage3_13[24],stage3_12[36]}
   );
   gpc606_5 gpc3406 (
      {stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[19],stage3_14[24],stage3_13[25],stage3_12[37]}
   );
   gpc606_5 gpc3407 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[20],stage3_14[25],stage3_13[26],stage3_12[38]}
   );
   gpc606_5 gpc3408 (
      {stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94], stage2_12[95]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[21],stage3_14[26],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc3409 (
      {stage2_12[96], stage2_12[97], stage2_12[98], stage2_12[99], stage2_12[100], stage2_12[101]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[22],stage3_14[27],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc3410 (
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[23],stage3_14[28],stage3_13[29]}
   );
   gpc606_5 gpc3411 (
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[24],stage3_14[29],stage3_13[30]}
   );
   gpc606_5 gpc3412 (
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[25],stage3_14[30],stage3_13[31]}
   );
   gpc606_5 gpc3413 (
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[26],stage3_14[31],stage3_13[32]}
   );
   gpc615_5 gpc3414 (
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94]},
      {stage2_14[72]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[27],stage3_14[32],stage3_13[33]}
   );
   gpc615_5 gpc3415 (
      {stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_15[30]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[5],stage3_16[17],stage3_15[28],stage3_14[33]}
   );
   gpc615_5 gpc3416 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[31]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[6],stage3_16[18],stage3_15[29],stage3_14[34]}
   );
   gpc615_5 gpc3417 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[32]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[7],stage3_16[19],stage3_15[30],stage3_14[35]}
   );
   gpc615_5 gpc3418 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[33]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[8],stage3_16[20],stage3_15[31],stage3_14[36]}
   );
   gpc615_5 gpc3419 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[34]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[9],stage3_16[21],stage3_15[32],stage3_14[37]}
   );
   gpc615_5 gpc3420 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], stage2_14[102]},
      {stage2_15[35]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[10],stage3_16[22],stage3_15[33],stage3_14[38]}
   );
   gpc615_5 gpc3421 (
      {stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_15[36]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[11],stage3_16[23],stage3_15[34],stage3_14[39]}
   );
   gpc615_5 gpc3422 (
      {stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111], stage2_14[112]},
      {stage2_15[37]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[12],stage3_16[24],stage3_15[35],stage3_14[40]}
   );
   gpc615_5 gpc3423 (
      {stage2_14[113], stage2_14[114], stage2_14[115], stage2_14[116], stage2_14[117]},
      {stage2_15[38]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[13],stage3_16[25],stage3_15[36],stage3_14[41]}
   );
   gpc615_5 gpc3424 (
      {stage2_14[118], stage2_14[119], stage2_14[120], stage2_14[121], stage2_14[122]},
      {stage2_15[39]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[14],stage3_16[26],stage3_15[37],stage3_14[42]}
   );
   gpc615_5 gpc3425 (
      {stage2_14[123], stage2_14[124], stage2_14[125], stage2_14[126], stage2_14[127]},
      {stage2_15[40]},
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage3_18[10],stage3_17[15],stage3_16[27],stage3_15[38],stage3_14[43]}
   );
   gpc615_5 gpc3426 (
      {stage2_14[128], stage2_14[129], stage2_14[130], stage2_14[131], stage2_14[132]},
      {stage2_15[41]},
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage3_18[11],stage3_17[16],stage3_16[28],stage3_15[39],stage3_14[44]}
   );
   gpc2135_5 gpc3427 (
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46]},
      {stage2_16[72], stage2_16[73], stage2_16[74]},
      {stage2_17[0]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[12],stage3_17[17],stage3_16[29],stage3_15[40]}
   );
   gpc606_5 gpc3428 (
      {stage2_15[47], stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[1],stage3_18[13],stage3_17[18],stage3_16[30],stage3_15[41]}
   );
   gpc606_5 gpc3429 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[2],stage3_18[14],stage3_17[19],stage3_16[31],stage3_15[42]}
   );
   gpc606_5 gpc3430 (
      {stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[3],stage3_18[15],stage3_17[20],stage3_16[32],stage3_15[43]}
   );
   gpc606_5 gpc3431 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69], stage2_15[70]},
      {stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24]},
      {stage3_19[4],stage3_18[16],stage3_17[21],stage3_16[33],stage3_15[44]}
   );
   gpc606_5 gpc3432 (
      {stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76]},
      {stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30]},
      {stage3_19[5],stage3_18[17],stage3_17[22],stage3_16[34],stage3_15[45]}
   );
   gpc606_5 gpc3433 (
      {stage2_15[77], stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36]},
      {stage3_19[6],stage3_18[18],stage3_17[23],stage3_16[35],stage3_15[46]}
   );
   gpc606_5 gpc3434 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87], stage2_15[88]},
      {stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42]},
      {stage3_19[7],stage3_18[19],stage3_17[24],stage3_16[36],stage3_15[47]}
   );
   gpc606_5 gpc3435 (
      {stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92], stage2_15[93], stage2_15[94]},
      {stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48]},
      {stage3_19[8],stage3_18[20],stage3_17[25],stage3_16[37],stage3_15[48]}
   );
   gpc606_5 gpc3436 (
      {stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80]},
      {stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6], stage2_18[7]},
      {stage3_20[0],stage3_19[9],stage3_18[21],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc3437 (
      {stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[10],stage3_18[22],stage3_17[27]}
   );
   gpc606_5 gpc3438 (
      {stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[11],stage3_18[23],stage3_17[28]}
   );
   gpc606_5 gpc3439 (
      {stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[12],stage3_18[24],stage3_17[29]}
   );
   gpc606_5 gpc3440 (
      {stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[13],stage3_18[25],stage3_17[30]}
   );
   gpc606_5 gpc3441 (
      {stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[5],stage3_19[14],stage3_18[26],stage3_17[31]}
   );
   gpc606_5 gpc3442 (
      {stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83], stage2_17[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage3_21[5],stage3_20[6],stage3_19[15],stage3_18[27],stage3_17[32]}
   );
   gpc606_5 gpc3443 (
      {stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89], stage2_17[90]},
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage3_21[6],stage3_20[7],stage3_19[16],stage3_18[28],stage3_17[33]}
   );
   gpc606_5 gpc3444 (
      {stage2_17[91], stage2_17[92], stage2_17[93], stage2_17[94], stage2_17[95], stage2_17[96]},
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage3_21[7],stage3_20[8],stage3_19[17],stage3_18[29],stage3_17[34]}
   );
   gpc606_5 gpc3445 (
      {stage2_17[97], stage2_17[98], stage2_17[99], stage2_17[100], stage2_17[101], stage2_17[102]},
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage3_21[8],stage3_20[9],stage3_19[18],stage3_18[30],stage3_17[35]}
   );
   gpc606_5 gpc3446 (
      {stage2_17[103], stage2_17[104], stage2_17[105], stage2_17[106], stage2_17[107], stage2_17[108]},
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage3_21[9],stage3_20[10],stage3_19[19],stage3_18[31],stage3_17[36]}
   );
   gpc1343_5 gpc3447 (
      {stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[10],stage3_20[11],stage3_19[20],stage3_18[32]}
   );
   gpc1343_5 gpc3448 (
      {stage2_18[11], stage2_18[12], stage2_18[13]},
      {stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[11],stage3_20[12],stage3_19[21],stage3_18[33]}
   );
   gpc1343_5 gpc3449 (
      {stage2_18[14], stage2_18[15], stage2_18[16]},
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71]},
      {stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_21[2]},
      {stage3_22[2],stage3_21[12],stage3_20[13],stage3_19[22],stage3_18[34]}
   );
   gpc1343_5 gpc3450 (
      {stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[72], stage2_19[73], stage2_19[74], stage2_19[75]},
      {stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage2_21[3]},
      {stage3_22[3],stage3_21[13],stage3_20[14],stage3_19[23],stage3_18[35]}
   );
   gpc615_5 gpc3451 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[76]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[4],stage3_21[14],stage3_20[15],stage3_19[24],stage3_18[36]}
   );
   gpc615_5 gpc3452 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[77]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[5],stage3_21[15],stage3_20[16],stage3_19[25],stage3_18[37]}
   );
   gpc615_5 gpc3453 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[78]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[6],stage3_21[16],stage3_20[17],stage3_19[26],stage3_18[38]}
   );
   gpc615_5 gpc3454 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[79]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[7],stage3_21[17],stage3_20[18],stage3_19[27],stage3_18[39]}
   );
   gpc615_5 gpc3455 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[80]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[8],stage3_21[18],stage3_20[19],stage3_19[28],stage3_18[40]}
   );
   gpc615_5 gpc3456 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[81]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[9],stage3_21[19],stage3_20[20],stage3_19[29],stage3_18[41]}
   );
   gpc615_5 gpc3457 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[82]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[10],stage3_21[20],stage3_20[21],stage3_19[30],stage3_18[42]}
   );
   gpc615_5 gpc3458 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[83]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[11],stage3_21[21],stage3_20[22],stage3_19[31],stage3_18[43]}
   );
   gpc615_5 gpc3459 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[84]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[12],stage3_21[22],stage3_20[23],stage3_19[32],stage3_18[44]}
   );
   gpc615_5 gpc3460 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[85]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[13],stage3_21[23],stage3_20[24],stage3_19[33],stage3_18[45]}
   );
   gpc615_5 gpc3461 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[86]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[14],stage3_21[24],stage3_20[25],stage3_19[34],stage3_18[46]}
   );
   gpc615_5 gpc3462 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[87]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[15],stage3_21[25],stage3_20[26],stage3_19[35],stage3_18[47]}
   );
   gpc615_5 gpc3463 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[84]},
      {stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage3_23[0],stage3_22[16],stage3_21[26],stage3_20[27],stage3_19[36]}
   );
   gpc615_5 gpc3464 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[85]},
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage3_23[1],stage3_22[17],stage3_21[27],stage3_20[28],stage3_19[37]}
   );
   gpc606_5 gpc3465 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[18],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3466 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[3],stage3_22[19],stage3_21[29],stage3_20[30]}
   );
   gpc606_5 gpc3467 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[4],stage3_22[20],stage3_21[30],stage3_20[31]}
   );
   gpc606_5 gpc3468 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[5],stage3_22[21],stage3_21[31],stage3_20[32]}
   );
   gpc606_5 gpc3469 (
      {stage2_20[110], stage2_20[111], stage2_20[112], stage2_20[113], stage2_20[114], stage2_20[115]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[6],stage3_22[22],stage3_21[32],stage3_20[33]}
   );
   gpc1163_5 gpc3470 (
      {stage2_21[16], stage2_21[17], stage2_21[18]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage2_23[0]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[5],stage3_23[7],stage3_22[23],stage3_21[33]}
   );
   gpc1163_5 gpc3471 (
      {stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[1]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[6],stage3_23[8],stage3_22[24],stage3_21[34]}
   );
   gpc1163_5 gpc3472 (
      {stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage2_23[2]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[7],stage3_23[9],stage3_22[25],stage3_21[35]}
   );
   gpc1163_5 gpc3473 (
      {stage2_21[25], stage2_21[26], stage2_21[27]},
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53]},
      {stage2_23[3]},
      {stage2_24[3]},
      {stage3_25[3],stage3_24[8],stage3_23[10],stage3_22[26],stage3_21[36]}
   );
   gpc1163_5 gpc3474 (
      {stage2_21[28], stage2_21[29], stage2_21[30]},
      {stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[4]},
      {stage2_24[4]},
      {stage3_25[4],stage3_24[9],stage3_23[11],stage3_22[27],stage3_21[37]}
   );
   gpc1163_5 gpc3475 (
      {stage2_21[31], stage2_21[32], stage2_21[33]},
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65]},
      {stage2_23[5]},
      {stage2_24[5]},
      {stage3_25[5],stage3_24[10],stage3_23[12],stage3_22[28],stage3_21[38]}
   );
   gpc606_5 gpc3476 (
      {stage2_21[34], stage2_21[35], stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[6],stage3_24[11],stage3_23[13],stage3_22[29],stage3_21[39]}
   );
   gpc606_5 gpc3477 (
      {stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[7],stage3_24[12],stage3_23[14],stage3_22[30],stage3_21[40]}
   );
   gpc606_5 gpc3478 (
      {stage2_21[46], stage2_21[47], stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[8],stage3_24[13],stage3_23[15],stage3_22[31],stage3_21[41]}
   );
   gpc606_5 gpc3479 (
      {stage2_21[52], stage2_21[53], stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[9],stage3_24[14],stage3_23[16],stage3_22[32],stage3_21[42]}
   );
   gpc606_5 gpc3480 (
      {stage2_21[58], stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[10],stage3_24[15],stage3_23[17],stage3_22[33],stage3_21[43]}
   );
   gpc615_5 gpc3481 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40]},
      {stage2_24[6]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[11],stage3_24[16],stage3_23[18]}
   );
   gpc615_5 gpc3482 (
      {stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45]},
      {stage2_24[7]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[1],stage3_25[12],stage3_24[17],stage3_23[19]}
   );
   gpc615_5 gpc3483 (
      {stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_24[8]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[2],stage3_25[13],stage3_24[18],stage3_23[20]}
   );
   gpc615_5 gpc3484 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55]},
      {stage2_24[9]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[3],stage3_25[14],stage3_24[19],stage3_23[21]}
   );
   gpc615_5 gpc3485 (
      {stage2_23[56], stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60]},
      {stage2_24[10]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[4],stage3_25[15],stage3_24[20],stage3_23[22]}
   );
   gpc615_5 gpc3486 (
      {stage2_23[61], stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65]},
      {stage2_24[11]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[5],stage3_25[16],stage3_24[21],stage3_23[23]}
   );
   gpc615_5 gpc3487 (
      {stage2_23[66], stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70]},
      {stage2_24[12]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[6],stage3_25[17],stage3_24[22],stage3_23[24]}
   );
   gpc615_5 gpc3488 (
      {stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75]},
      {stage2_24[13]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[7],stage3_25[18],stage3_24[23],stage3_23[25]}
   );
   gpc615_5 gpc3489 (
      {stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_24[14]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[8],stage3_25[19],stage3_24[24],stage3_23[26]}
   );
   gpc615_5 gpc3490 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85]},
      {stage2_24[15]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[9],stage3_25[20],stage3_24[25],stage3_23[27]}
   );
   gpc615_5 gpc3491 (
      {stage2_23[86], stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90]},
      {stage2_24[16]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[10],stage3_25[21],stage3_24[26],stage3_23[28]}
   );
   gpc606_5 gpc3492 (
      {stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[11],stage3_26[11],stage3_25[22],stage3_24[27]}
   );
   gpc606_5 gpc3493 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[12],stage3_26[12],stage3_25[23],stage3_24[28]}
   );
   gpc606_5 gpc3494 (
      {stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[13],stage3_26[13],stage3_25[24],stage3_24[29]}
   );
   gpc606_5 gpc3495 (
      {stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[14],stage3_26[14],stage3_25[25],stage3_24[30]}
   );
   gpc606_5 gpc3496 (
      {stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[15],stage3_26[15],stage3_25[26],stage3_24[31]}
   );
   gpc606_5 gpc3497 (
      {stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[16],stage3_26[16],stage3_25[27],stage3_24[32]}
   );
   gpc606_5 gpc3498 (
      {stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[17],stage3_26[17],stage3_25[28],stage3_24[33]}
   );
   gpc606_5 gpc3499 (
      {stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[18],stage3_26[18],stage3_25[29],stage3_24[34]}
   );
   gpc606_5 gpc3500 (
      {stage2_24[65], stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70]},
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53]},
      {stage3_28[8],stage3_27[19],stage3_26[19],stage3_25[30],stage3_24[35]}
   );
   gpc606_5 gpc3501 (
      {stage2_24[71], stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76]},
      {stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59]},
      {stage3_28[9],stage3_27[20],stage3_26[20],stage3_25[31],stage3_24[36]}
   );
   gpc606_5 gpc3502 (
      {stage2_24[77], stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82]},
      {stage2_26[60], stage2_26[61], stage2_26[62], stage2_26[63], stage2_26[64], stage2_26[65]},
      {stage3_28[10],stage3_27[21],stage3_26[21],stage3_25[32],stage3_24[37]}
   );
   gpc606_5 gpc3503 (
      {stage2_24[83], stage2_24[84], stage2_24[85], stage2_24[86], stage2_24[87], stage2_24[88]},
      {stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71]},
      {stage3_28[11],stage3_27[22],stage3_26[22],stage3_25[33],stage3_24[38]}
   );
   gpc606_5 gpc3504 (
      {stage2_24[89], stage2_24[90], stage2_24[91], stage2_24[92], stage2_24[93], stage2_24[94]},
      {stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76], stage2_26[77]},
      {stage3_28[12],stage3_27[23],stage3_26[23],stage3_25[34],stage3_24[39]}
   );
   gpc606_5 gpc3505 (
      {stage2_24[95], stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], 1'b0},
      {stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage3_28[13],stage3_27[24],stage3_26[24],stage3_25[35],stage3_24[40]}
   );
   gpc606_5 gpc3506 (
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[14],stage3_27[25],stage3_26[25],stage3_25[36]}
   );
   gpc606_5 gpc3507 (
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[15],stage3_27[26],stage3_26[26],stage3_25[37]}
   );
   gpc606_5 gpc3508 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[16],stage3_27[27],stage3_26[27],stage3_25[38]}
   );
   gpc606_5 gpc3509 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], 1'b0, 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[17],stage3_27[28],stage3_26[28],stage3_25[39]}
   );
   gpc615_5 gpc3510 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88]},
      {stage2_27[24]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[4],stage3_28[18],stage3_27[29],stage3_26[29]}
   );
   gpc615_5 gpc3511 (
      {stage2_26[89], stage2_26[90], stage2_26[91], stage2_26[92], stage2_26[93]},
      {stage2_27[25]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[5],stage3_28[19],stage3_27[30],stage3_26[30]}
   );
   gpc615_5 gpc3512 (
      {stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97], stage2_26[98]},
      {stage2_27[26]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[6],stage3_28[20],stage3_27[31],stage3_26[31]}
   );
   gpc606_5 gpc3513 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[3],stage3_29[7],stage3_28[21],stage3_27[32]}
   );
   gpc606_5 gpc3514 (
      {stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[4],stage3_29[8],stage3_28[22],stage3_27[33]}
   );
   gpc606_5 gpc3515 (
      {stage2_27[39], stage2_27[40], stage2_27[41], stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[5],stage3_29[9],stage3_28[23],stage3_27[34]}
   );
   gpc615_5 gpc3516 (
      {stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48], stage2_27[49]},
      {stage2_28[18]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[6],stage3_29[10],stage3_28[24],stage3_27[35]}
   );
   gpc615_5 gpc3517 (
      {stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54]},
      {stage2_28[19]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[7],stage3_29[11],stage3_28[25],stage3_27[36]}
   );
   gpc615_5 gpc3518 (
      {stage2_27[55], stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[20]},
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage3_31[5],stage3_30[8],stage3_29[12],stage3_28[26],stage3_27[37]}
   );
   gpc615_5 gpc3519 (
      {stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63], stage2_27[64]},
      {stage2_28[21]},
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage3_31[6],stage3_30[9],stage3_29[13],stage3_28[27],stage3_27[38]}
   );
   gpc615_5 gpc3520 (
      {stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_28[22]},
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage3_31[7],stage3_30[10],stage3_29[14],stage3_28[28],stage3_27[39]}
   );
   gpc606_5 gpc3521 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[8],stage3_30[11],stage3_29[15],stage3_28[29]}
   );
   gpc606_5 gpc3522 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[9],stage3_30[12],stage3_29[16],stage3_28[30]}
   );
   gpc606_5 gpc3523 (
      {stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[10],stage3_30[13],stage3_29[17],stage3_28[31]}
   );
   gpc606_5 gpc3524 (
      {stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[11],stage3_30[14],stage3_29[18],stage3_28[32]}
   );
   gpc606_5 gpc3525 (
      {stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[12],stage3_30[15],stage3_29[19],stage3_28[33]}
   );
   gpc606_5 gpc3526 (
      {stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[13],stage3_30[16],stage3_29[20],stage3_28[34]}
   );
   gpc615_5 gpc3527 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[48]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[14],stage3_30[17],stage3_29[21],stage3_28[35]}
   );
   gpc615_5 gpc3528 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[49]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[15],stage3_30[18],stage3_29[22],stage3_28[36]}
   );
   gpc1163_5 gpc3529 (
      {stage2_29[50], stage2_29[51], stage2_29[52]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[8],stage3_31[16],stage3_30[19],stage3_29[23]}
   );
   gpc1163_5 gpc3530 (
      {stage2_29[53], stage2_29[54], stage2_29[55]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[9],stage3_31[17],stage3_30[20],stage3_29[24]}
   );
   gpc1163_5 gpc3531 (
      {stage2_29[56], stage2_29[57], stage2_29[58]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[10],stage3_31[18],stage3_30[21],stage3_29[25]}
   );
   gpc1163_5 gpc3532 (
      {stage2_29[59], stage2_29[60], stage2_29[61]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[11],stage3_31[19],stage3_30[22],stage3_29[26]}
   );
   gpc1163_5 gpc3533 (
      {stage2_29[62], stage2_29[63], stage2_29[64]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[12],stage3_31[20],stage3_30[23],stage3_29[27]}
   );
   gpc606_5 gpc3534 (
      {stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[13],stage3_31[21],stage3_30[24],stage3_29[28]}
   );
   gpc606_5 gpc3535 (
      {stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[14],stage3_31[22],stage3_30[25],stage3_29[29]}
   );
   gpc606_5 gpc3536 (
      {stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[15],stage3_31[23],stage3_30[26],stage3_29[30]}
   );
   gpc606_5 gpc3537 (
      {stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[16],stage3_31[24],stage3_30[27],stage3_29[31]}
   );
   gpc606_5 gpc3538 (
      {stage2_29[89], stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[17],stage3_31[25],stage3_30[28],stage3_29[32]}
   );
   gpc606_5 gpc3539 (
      {stage2_29[95], stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[18],stage3_31[26],stage3_30[29],stage3_29[33]}
   );
   gpc606_5 gpc3540 (
      {stage2_29[101], stage2_29[102], stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[19],stage3_31[27],stage3_30[30],stage3_29[34]}
   );
   gpc606_5 gpc3541 (
      {stage2_29[107], stage2_29[108], stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[20],stage3_31[28],stage3_30[31],stage3_29[35]}
   );
   gpc606_5 gpc3542 (
      {stage2_29[113], stage2_29[114], stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[21],stage3_31[29],stage3_30[32],stage3_29[36]}
   );
   gpc606_5 gpc3543 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_32[5], stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10]},
      {stage3_34[0],stage3_33[14],stage3_32[22],stage3_31[30],stage3_30[33]}
   );
   gpc606_5 gpc3544 (
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_32[11], stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16]},
      {stage3_34[1],stage3_33[15],stage3_32[23],stage3_31[31],stage3_30[34]}
   );
   gpc606_5 gpc3545 (
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22]},
      {stage3_34[2],stage3_33[16],stage3_32[24],stage3_31[32],stage3_30[35]}
   );
   gpc606_5 gpc3546 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101]},
      {stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28]},
      {stage3_34[3],stage3_33[17],stage3_32[25],stage3_31[33],stage3_30[36]}
   );
   gpc606_5 gpc3547 (
      {stage2_30[102], stage2_30[103], stage2_30[104], stage2_30[105], stage2_30[106], stage2_30[107]},
      {stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34]},
      {stage3_34[4],stage3_33[18],stage3_32[26],stage3_31[34],stage3_30[37]}
   );
   gpc606_5 gpc3548 (
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[5],stage3_33[19],stage3_32[27],stage3_31[35]}
   );
   gpc606_5 gpc3549 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[6],stage3_33[20],stage3_32[28],stage3_31[36]}
   );
   gpc606_5 gpc3550 (
      {stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[7],stage3_33[21],stage3_32[29],stage3_31[37]}
   );
   gpc606_5 gpc3551 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[8],stage3_33[22],stage3_32[30],stage3_31[38]}
   );
   gpc606_5 gpc3552 (
      {stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[9],stage3_33[23],stage3_32[31]}
   );
   gpc606_5 gpc3553 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45], stage2_32[46]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[10],stage3_33[24],stage3_32[32]}
   );
   gpc606_5 gpc3554 (
      {stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50], stage2_32[51], stage2_32[52]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[6],stage3_34[11],stage3_33[25],stage3_32[33]}
   );
   gpc606_5 gpc3555 (
      {stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56], stage2_32[57], stage2_32[58]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[7],stage3_34[12],stage3_33[26],stage3_32[34]}
   );
   gpc606_5 gpc3556 (
      {stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62], stage2_32[63], stage2_32[64]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[8],stage3_34[13],stage3_33[27],stage3_32[35]}
   );
   gpc606_5 gpc3557 (
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[5],stage3_35[9],stage3_34[14],stage3_33[28]}
   );
   gpc606_5 gpc3558 (
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[6],stage3_35[10],stage3_34[15],stage3_33[29]}
   );
   gpc1_1 gpc3559 (
      {stage2_0[21]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3560 (
      {stage2_2[43]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3561 (
      {stage2_2[44]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3562 (
      {stage2_2[45]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3563 (
      {stage2_2[46]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3564 (
      {stage2_2[47]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3565 (
      {stage2_2[48]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3566 (
      {stage2_2[49]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3567 (
      {stage2_2[50]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3568 (
      {stage2_4[82]},
      {stage3_4[35]}
   );
   gpc1_1 gpc3569 (
      {stage2_4[83]},
      {stage3_4[36]}
   );
   gpc1_1 gpc3570 (
      {stage2_4[84]},
      {stage3_4[37]}
   );
   gpc1_1 gpc3571 (
      {stage2_4[85]},
      {stage3_4[38]}
   );
   gpc1_1 gpc3572 (
      {stage2_4[86]},
      {stage3_4[39]}
   );
   gpc1_1 gpc3573 (
      {stage2_4[87]},
      {stage3_4[40]}
   );
   gpc1_1 gpc3574 (
      {stage2_4[88]},
      {stage3_4[41]}
   );
   gpc1_1 gpc3575 (
      {stage2_4[89]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3576 (
      {stage2_4[90]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3577 (
      {stage2_5[71]},
      {stage3_5[36]}
   );
   gpc1_1 gpc3578 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3579 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3580 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3581 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3582 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3583 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3584 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3585 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3586 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3587 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3588 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3589 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3590 (
      {stage2_6[83]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3591 (
      {stage2_6[84]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3592 (
      {stage2_6[85]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3593 (
      {stage2_6[86]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3594 (
      {stage2_6[87]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3595 (
      {stage2_6[88]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3596 (
      {stage2_6[89]},
      {stage3_6[38]}
   );
   gpc1_1 gpc3597 (
      {stage2_6[90]},
      {stage3_6[39]}
   );
   gpc1_1 gpc3598 (
      {stage2_6[91]},
      {stage3_6[40]}
   );
   gpc1_1 gpc3599 (
      {stage2_6[92]},
      {stage3_6[41]}
   );
   gpc1_1 gpc3600 (
      {stage2_6[93]},
      {stage3_6[42]}
   );
   gpc1_1 gpc3601 (
      {stage2_7[70]},
      {stage3_7[29]}
   );
   gpc1_1 gpc3602 (
      {stage2_7[71]},
      {stage3_7[30]}
   );
   gpc1_1 gpc3603 (
      {stage2_7[72]},
      {stage3_7[31]}
   );
   gpc1_1 gpc3604 (
      {stage2_7[73]},
      {stage3_7[32]}
   );
   gpc1_1 gpc3605 (
      {stage2_7[74]},
      {stage3_7[33]}
   );
   gpc1_1 gpc3606 (
      {stage2_7[75]},
      {stage3_7[34]}
   );
   gpc1_1 gpc3607 (
      {stage2_7[76]},
      {stage3_7[35]}
   );
   gpc1_1 gpc3608 (
      {stage2_7[77]},
      {stage3_7[36]}
   );
   gpc1_1 gpc3609 (
      {stage2_7[78]},
      {stage3_7[37]}
   );
   gpc1_1 gpc3610 (
      {stage2_7[79]},
      {stage3_7[38]}
   );
   gpc1_1 gpc3611 (
      {stage2_7[80]},
      {stage3_7[39]}
   );
   gpc1_1 gpc3612 (
      {stage2_7[81]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3613 (
      {stage2_7[82]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3614 (
      {stage2_7[83]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3615 (
      {stage2_7[84]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3616 (
      {stage2_7[85]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3617 (
      {stage2_7[86]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3618 (
      {stage2_7[87]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3619 (
      {stage2_7[88]},
      {stage3_7[47]}
   );
   gpc1_1 gpc3620 (
      {stage2_7[89]},
      {stage3_7[48]}
   );
   gpc1_1 gpc3621 (
      {stage2_7[90]},
      {stage3_7[49]}
   );
   gpc1_1 gpc3622 (
      {stage2_7[91]},
      {stage3_7[50]}
   );
   gpc1_1 gpc3623 (
      {stage2_7[92]},
      {stage3_7[51]}
   );
   gpc1_1 gpc3624 (
      {stage2_7[93]},
      {stage3_7[52]}
   );
   gpc1_1 gpc3625 (
      {stage2_7[94]},
      {stage3_7[53]}
   );
   gpc1_1 gpc3626 (
      {stage2_7[95]},
      {stage3_7[54]}
   );
   gpc1_1 gpc3627 (
      {stage2_7[96]},
      {stage3_7[55]}
   );
   gpc1_1 gpc3628 (
      {stage2_7[97]},
      {stage3_7[56]}
   );
   gpc1_1 gpc3629 (
      {stage2_7[98]},
      {stage3_7[57]}
   );
   gpc1_1 gpc3630 (
      {stage2_7[99]},
      {stage3_7[58]}
   );
   gpc1_1 gpc3631 (
      {stage2_7[100]},
      {stage3_7[59]}
   );
   gpc1_1 gpc3632 (
      {stage2_7[101]},
      {stage3_7[60]}
   );
   gpc1_1 gpc3633 (
      {stage2_7[102]},
      {stage3_7[61]}
   );
   gpc1_1 gpc3634 (
      {stage2_7[103]},
      {stage3_7[62]}
   );
   gpc1_1 gpc3635 (
      {stage2_7[104]},
      {stage3_7[63]}
   );
   gpc1_1 gpc3636 (
      {stage2_7[105]},
      {stage3_7[64]}
   );
   gpc1_1 gpc3637 (
      {stage2_7[106]},
      {stage3_7[65]}
   );
   gpc1_1 gpc3638 (
      {stage2_7[107]},
      {stage3_7[66]}
   );
   gpc1_1 gpc3639 (
      {stage2_7[108]},
      {stage3_7[67]}
   );
   gpc1_1 gpc3640 (
      {stage2_7[109]},
      {stage3_7[68]}
   );
   gpc1_1 gpc3641 (
      {stage2_9[36]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3642 (
      {stage2_9[37]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3643 (
      {stage2_9[38]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3644 (
      {stage2_9[39]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3645 (
      {stage2_9[40]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3646 (
      {stage2_9[41]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3647 (
      {stage2_9[42]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3648 (
      {stage2_9[43]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3649 (
      {stage2_9[44]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3650 (
      {stage2_9[45]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3651 (
      {stage2_9[46]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3652 (
      {stage2_9[47]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3653 (
      {stage2_9[48]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[49]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[50]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[51]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[52]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3658 (
      {stage2_9[53]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3659 (
      {stage2_9[54]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3660 (
      {stage2_9[55]},
      {stage3_9[50]}
   );
   gpc1_1 gpc3661 (
      {stage2_9[56]},
      {stage3_9[51]}
   );
   gpc1_1 gpc3662 (
      {stage2_9[57]},
      {stage3_9[52]}
   );
   gpc1_1 gpc3663 (
      {stage2_9[58]},
      {stage3_9[53]}
   );
   gpc1_1 gpc3664 (
      {stage2_9[59]},
      {stage3_9[54]}
   );
   gpc1_1 gpc3665 (
      {stage2_9[60]},
      {stage3_9[55]}
   );
   gpc1_1 gpc3666 (
      {stage2_9[61]},
      {stage3_9[56]}
   );
   gpc1_1 gpc3667 (
      {stage2_9[62]},
      {stage3_9[57]}
   );
   gpc1_1 gpc3668 (
      {stage2_9[63]},
      {stage3_9[58]}
   );
   gpc1_1 gpc3669 (
      {stage2_9[64]},
      {stage3_9[59]}
   );
   gpc1_1 gpc3670 (
      {stage2_9[65]},
      {stage3_9[60]}
   );
   gpc1_1 gpc3671 (
      {stage2_9[66]},
      {stage3_9[61]}
   );
   gpc1_1 gpc3672 (
      {stage2_9[67]},
      {stage3_9[62]}
   );
   gpc1_1 gpc3673 (
      {stage2_9[68]},
      {stage3_9[63]}
   );
   gpc1_1 gpc3674 (
      {stage2_9[69]},
      {stage3_9[64]}
   );
   gpc1_1 gpc3675 (
      {stage2_9[70]},
      {stage3_9[65]}
   );
   gpc1_1 gpc3676 (
      {stage2_9[71]},
      {stage3_9[66]}
   );
   gpc1_1 gpc3677 (
      {stage2_9[72]},
      {stage3_9[67]}
   );
   gpc1_1 gpc3678 (
      {stage2_9[73]},
      {stage3_9[68]}
   );
   gpc1_1 gpc3679 (
      {stage2_9[74]},
      {stage3_9[69]}
   );
   gpc1_1 gpc3680 (
      {stage2_10[88]},
      {stage3_10[28]}
   );
   gpc1_1 gpc3681 (
      {stage2_11[80]},
      {stage3_11[32]}
   );
   gpc1_1 gpc3682 (
      {stage2_11[81]},
      {stage3_11[33]}
   );
   gpc1_1 gpc3683 (
      {stage2_11[82]},
      {stage3_11[34]}
   );
   gpc1_1 gpc3684 (
      {stage2_11[83]},
      {stage3_11[35]}
   );
   gpc1_1 gpc3685 (
      {stage2_11[84]},
      {stage3_11[36]}
   );
   gpc1_1 gpc3686 (
      {stage2_11[85]},
      {stage3_11[37]}
   );
   gpc1_1 gpc3687 (
      {stage2_11[86]},
      {stage3_11[38]}
   );
   gpc1_1 gpc3688 (
      {stage2_11[87]},
      {stage3_11[39]}
   );
   gpc1_1 gpc3689 (
      {stage2_11[88]},
      {stage3_11[40]}
   );
   gpc1_1 gpc3690 (
      {stage2_11[89]},
      {stage3_11[41]}
   );
   gpc1_1 gpc3691 (
      {stage2_11[90]},
      {stage3_11[42]}
   );
   gpc1_1 gpc3692 (
      {stage2_11[91]},
      {stage3_11[43]}
   );
   gpc1_1 gpc3693 (
      {stage2_12[102]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3694 (
      {stage2_13[95]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3695 (
      {stage2_13[96]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3696 (
      {stage2_13[97]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3697 (
      {stage2_13[98]},
      {stage3_13[37]}
   );
   gpc1_1 gpc3698 (
      {stage2_13[99]},
      {stage3_13[38]}
   );
   gpc1_1 gpc3699 (
      {stage2_13[100]},
      {stage3_13[39]}
   );
   gpc1_1 gpc3700 (
      {stage2_13[101]},
      {stage3_13[40]}
   );
   gpc1_1 gpc3701 (
      {stage2_14[133]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3702 (
      {stage2_14[134]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3703 (
      {stage2_14[135]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3704 (
      {stage2_14[136]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3705 (
      {stage2_14[137]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3706 (
      {stage2_14[138]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[95]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[96]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[97]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[98]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[99]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[100]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[101]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[102]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[103]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[104]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3717 (
      {stage2_15[105]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3718 (
      {stage2_15[106]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3719 (
      {stage2_15[107]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3720 (
      {stage2_15[108]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3721 (
      {stage2_15[109]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3722 (
      {stage2_15[110]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3723 (
      {stage2_15[111]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3724 (
      {stage2_15[112]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3725 (
      {stage2_15[113]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3726 (
      {stage2_15[114]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3727 (
      {stage2_15[115]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3728 (
      {stage2_15[116]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3729 (
      {stage2_15[117]},
      {stage3_15[71]}
   );
   gpc1_1 gpc3730 (
      {stage2_15[118]},
      {stage3_15[72]}
   );
   gpc1_1 gpc3731 (
      {stage2_15[119]},
      {stage3_15[73]}
   );
   gpc1_1 gpc3732 (
      {stage2_15[120]},
      {stage3_15[74]}
   );
   gpc1_1 gpc3733 (
      {stage2_15[121]},
      {stage3_15[75]}
   );
   gpc1_1 gpc3734 (
      {stage2_15[122]},
      {stage3_15[76]}
   );
   gpc1_1 gpc3735 (
      {stage2_15[123]},
      {stage3_15[77]}
   );
   gpc1_1 gpc3736 (
      {stage2_15[124]},
      {stage3_15[78]}
   );
   gpc1_1 gpc3737 (
      {stage2_15[125]},
      {stage3_15[79]}
   );
   gpc1_1 gpc3738 (
      {stage2_15[126]},
      {stage3_15[80]}
   );
   gpc1_1 gpc3739 (
      {stage2_15[127]},
      {stage3_15[81]}
   );
   gpc1_1 gpc3740 (
      {stage2_15[128]},
      {stage3_15[82]}
   );
   gpc1_1 gpc3741 (
      {stage2_15[129]},
      {stage3_15[83]}
   );
   gpc1_1 gpc3742 (
      {stage2_15[130]},
      {stage3_15[84]}
   );
   gpc1_1 gpc3743 (
      {stage2_15[131]},
      {stage3_15[85]}
   );
   gpc1_1 gpc3744 (
      {stage2_15[132]},
      {stage3_15[86]}
   );
   gpc1_1 gpc3745 (
      {stage2_15[133]},
      {stage3_15[87]}
   );
   gpc1_1 gpc3746 (
      {stage2_15[134]},
      {stage3_15[88]}
   );
   gpc1_1 gpc3747 (
      {stage2_15[135]},
      {stage3_15[89]}
   );
   gpc1_1 gpc3748 (
      {stage2_16[81]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3749 (
      {stage2_16[82]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3750 (
      {stage2_16[83]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3751 (
      {stage2_16[84]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3752 (
      {stage2_16[85]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3753 (
      {stage2_16[86]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3754 (
      {stage2_16[87]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3755 (
      {stage2_16[88]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3756 (
      {stage2_16[89]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3757 (
      {stage2_16[90]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3758 (
      {stage2_16[91]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3759 (
      {stage2_16[92]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3760 (
      {stage2_16[93]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3761 (
      {stage2_16[94]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3762 (
      {stage2_16[95]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3763 (
      {stage2_16[96]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3764 (
      {stage2_16[97]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3765 (
      {stage2_16[98]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3766 (
      {stage2_16[99]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3767 (
      {stage2_16[100]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3768 (
      {stage2_16[101]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3769 (
      {stage2_16[102]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3770 (
      {stage2_16[103]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3771 (
      {stage2_17[109]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3772 (
      {stage2_17[110]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3773 (
      {stage2_17[111]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3774 (
      {stage2_17[112]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3775 (
      {stage2_17[113]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3776 (
      {stage2_17[114]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3777 (
      {stage2_17[115]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3778 (
      {stage2_17[116]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3779 (
      {stage2_17[117]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3780 (
      {stage2_17[118]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3781 (
      {stage2_17[119]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3782 (
      {stage2_17[120]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3783 (
      {stage2_17[121]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3784 (
      {stage2_18[80]},
      {stage3_18[48]}
   );
   gpc1_1 gpc3785 (
      {stage2_18[81]},
      {stage3_18[49]}
   );
   gpc1_1 gpc3786 (
      {stage2_19[98]},
      {stage3_19[38]}
   );
   gpc1_1 gpc3787 (
      {stage2_19[99]},
      {stage3_19[39]}
   );
   gpc1_1 gpc3788 (
      {stage2_19[100]},
      {stage3_19[40]}
   );
   gpc1_1 gpc3789 (
      {stage2_19[101]},
      {stage3_19[41]}
   );
   gpc1_1 gpc3790 (
      {stage2_19[102]},
      {stage3_19[42]}
   );
   gpc1_1 gpc3791 (
      {stage2_19[103]},
      {stage3_19[43]}
   );
   gpc1_1 gpc3792 (
      {stage2_19[104]},
      {stage3_19[44]}
   );
   gpc1_1 gpc3793 (
      {stage2_19[105]},
      {stage3_19[45]}
   );
   gpc1_1 gpc3794 (
      {stage2_19[106]},
      {stage3_19[46]}
   );
   gpc1_1 gpc3795 (
      {stage2_19[107]},
      {stage3_19[47]}
   );
   gpc1_1 gpc3796 (
      {stage2_19[108]},
      {stage3_19[48]}
   );
   gpc1_1 gpc3797 (
      {stage2_19[109]},
      {stage3_19[49]}
   );
   gpc1_1 gpc3798 (
      {stage2_20[116]},
      {stage3_20[34]}
   );
   gpc1_1 gpc3799 (
      {stage2_20[117]},
      {stage3_20[35]}
   );
   gpc1_1 gpc3800 (
      {stage2_20[118]},
      {stage3_20[36]}
   );
   gpc1_1 gpc3801 (
      {stage2_20[119]},
      {stage3_20[37]}
   );
   gpc1_1 gpc3802 (
      {stage2_20[120]},
      {stage3_20[38]}
   );
   gpc1_1 gpc3803 (
      {stage2_20[121]},
      {stage3_20[39]}
   );
   gpc1_1 gpc3804 (
      {stage2_20[122]},
      {stage3_20[40]}
   );
   gpc1_1 gpc3805 (
      {stage2_20[123]},
      {stage3_20[41]}
   );
   gpc1_1 gpc3806 (
      {stage2_20[124]},
      {stage3_20[42]}
   );
   gpc1_1 gpc3807 (
      {stage2_20[125]},
      {stage3_20[43]}
   );
   gpc1_1 gpc3808 (
      {stage2_20[126]},
      {stage3_20[44]}
   );
   gpc1_1 gpc3809 (
      {stage2_20[127]},
      {stage3_20[45]}
   );
   gpc1_1 gpc3810 (
      {stage2_21[64]},
      {stage3_21[44]}
   );
   gpc1_1 gpc3811 (
      {stage2_21[65]},
      {stage3_21[45]}
   );
   gpc1_1 gpc3812 (
      {stage2_21[66]},
      {stage3_21[46]}
   );
   gpc1_1 gpc3813 (
      {stage2_21[67]},
      {stage3_21[47]}
   );
   gpc1_1 gpc3814 (
      {stage2_21[68]},
      {stage3_21[48]}
   );
   gpc1_1 gpc3815 (
      {stage2_21[69]},
      {stage3_21[49]}
   );
   gpc1_1 gpc3816 (
      {stage2_21[70]},
      {stage3_21[50]}
   );
   gpc1_1 gpc3817 (
      {stage2_21[71]},
      {stage3_21[51]}
   );
   gpc1_1 gpc3818 (
      {stage2_21[72]},
      {stage3_21[52]}
   );
   gpc1_1 gpc3819 (
      {stage2_21[73]},
      {stage3_21[53]}
   );
   gpc1_1 gpc3820 (
      {stage2_21[74]},
      {stage3_21[54]}
   );
   gpc1_1 gpc3821 (
      {stage2_21[75]},
      {stage3_21[55]}
   );
   gpc1_1 gpc3822 (
      {stage2_21[76]},
      {stage3_21[56]}
   );
   gpc1_1 gpc3823 (
      {stage2_21[77]},
      {stage3_21[57]}
   );
   gpc1_1 gpc3824 (
      {stage2_21[78]},
      {stage3_21[58]}
   );
   gpc1_1 gpc3825 (
      {stage2_22[66]},
      {stage3_22[34]}
   );
   gpc1_1 gpc3826 (
      {stage2_22[67]},
      {stage3_22[35]}
   );
   gpc1_1 gpc3827 (
      {stage2_22[68]},
      {stage3_22[36]}
   );
   gpc1_1 gpc3828 (
      {stage2_22[69]},
      {stage3_22[37]}
   );
   gpc1_1 gpc3829 (
      {stage2_22[70]},
      {stage3_22[38]}
   );
   gpc1_1 gpc3830 (
      {stage2_22[71]},
      {stage3_22[39]}
   );
   gpc1_1 gpc3831 (
      {stage2_22[72]},
      {stage3_22[40]}
   );
   gpc1_1 gpc3832 (
      {stage2_22[73]},
      {stage3_22[41]}
   );
   gpc1_1 gpc3833 (
      {stage2_22[74]},
      {stage3_22[42]}
   );
   gpc1_1 gpc3834 (
      {stage2_22[75]},
      {stage3_22[43]}
   );
   gpc1_1 gpc3835 (
      {stage2_22[76]},
      {stage3_22[44]}
   );
   gpc1_1 gpc3836 (
      {stage2_22[77]},
      {stage3_22[45]}
   );
   gpc1_1 gpc3837 (
      {stage2_22[78]},
      {stage3_22[46]}
   );
   gpc1_1 gpc3838 (
      {stage2_23[91]},
      {stage3_23[29]}
   );
   gpc1_1 gpc3839 (
      {stage2_23[92]},
      {stage3_23[30]}
   );
   gpc1_1 gpc3840 (
      {stage2_23[93]},
      {stage3_23[31]}
   );
   gpc1_1 gpc3841 (
      {stage2_23[94]},
      {stage3_23[32]}
   );
   gpc1_1 gpc3842 (
      {stage2_23[95]},
      {stage3_23[33]}
   );
   gpc1_1 gpc3843 (
      {stage2_23[96]},
      {stage3_23[34]}
   );
   gpc1_1 gpc3844 (
      {stage2_23[97]},
      {stage3_23[35]}
   );
   gpc1_1 gpc3845 (
      {stage2_23[98]},
      {stage3_23[36]}
   );
   gpc1_1 gpc3846 (
      {stage2_23[99]},
      {stage3_23[37]}
   );
   gpc1_1 gpc3847 (
      {stage2_23[100]},
      {stage3_23[38]}
   );
   gpc1_1 gpc3848 (
      {stage2_23[101]},
      {stage3_23[39]}
   );
   gpc1_1 gpc3849 (
      {stage2_23[102]},
      {stage3_23[40]}
   );
   gpc1_1 gpc3850 (
      {stage2_23[103]},
      {stage3_23[41]}
   );
   gpc1_1 gpc3851 (
      {stage2_23[104]},
      {stage3_23[42]}
   );
   gpc1_1 gpc3852 (
      {stage2_23[105]},
      {stage3_23[43]}
   );
   gpc1_1 gpc3853 (
      {stage2_23[106]},
      {stage3_23[44]}
   );
   gpc1_1 gpc3854 (
      {stage2_23[107]},
      {stage3_23[45]}
   );
   gpc1_1 gpc3855 (
      {stage2_23[108]},
      {stage3_23[46]}
   );
   gpc1_1 gpc3856 (
      {stage2_23[109]},
      {stage3_23[47]}
   );
   gpc1_1 gpc3857 (
      {stage2_27[70]},
      {stage3_27[40]}
   );
   gpc1_1 gpc3858 (
      {stage2_27[71]},
      {stage3_27[41]}
   );
   gpc1_1 gpc3859 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc3860 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc3861 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc3862 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc3863 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc3864 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc3865 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc3866 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc3867 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc3868 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc3869 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc3870 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc3871 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc3872 (
      {stage2_27[85]},
      {stage3_27[55]}
   );
   gpc1_1 gpc3873 (
      {stage2_27[86]},
      {stage3_27[56]}
   );
   gpc1_1 gpc3874 (
      {stage2_27[87]},
      {stage3_27[57]}
   );
   gpc1_1 gpc3875 (
      {stage2_27[88]},
      {stage3_27[58]}
   );
   gpc1_1 gpc3876 (
      {stage2_27[89]},
      {stage3_27[59]}
   );
   gpc1_1 gpc3877 (
      {stage2_27[90]},
      {stage3_27[60]}
   );
   gpc1_1 gpc3878 (
      {stage2_27[91]},
      {stage3_27[61]}
   );
   gpc1_1 gpc3879 (
      {stage2_27[92]},
      {stage3_27[62]}
   );
   gpc1_1 gpc3880 (
      {stage2_27[93]},
      {stage3_27[63]}
   );
   gpc1_1 gpc3881 (
      {stage2_27[94]},
      {stage3_27[64]}
   );
   gpc1_1 gpc3882 (
      {stage2_27[95]},
      {stage3_27[65]}
   );
   gpc1_1 gpc3883 (
      {stage2_27[96]},
      {stage3_27[66]}
   );
   gpc1_1 gpc3884 (
      {stage2_28[69]},
      {stage3_28[37]}
   );
   gpc1_1 gpc3885 (
      {stage2_28[70]},
      {stage3_28[38]}
   );
   gpc1_1 gpc3886 (
      {stage2_28[71]},
      {stage3_28[39]}
   );
   gpc1_1 gpc3887 (
      {stage2_28[72]},
      {stage3_28[40]}
   );
   gpc1_1 gpc3888 (
      {stage2_28[73]},
      {stage3_28[41]}
   );
   gpc1_1 gpc3889 (
      {stage2_28[74]},
      {stage3_28[42]}
   );
   gpc1_1 gpc3890 (
      {stage2_29[119]},
      {stage3_29[37]}
   );
   gpc1_1 gpc3891 (
      {stage2_29[120]},
      {stage3_29[38]}
   );
   gpc1_1 gpc3892 (
      {stage2_30[108]},
      {stage3_30[38]}
   );
   gpc1_1 gpc3893 (
      {stage2_30[109]},
      {stage3_30[39]}
   );
   gpc1_1 gpc3894 (
      {stage2_30[110]},
      {stage3_30[40]}
   );
   gpc1_1 gpc3895 (
      {stage2_30[111]},
      {stage3_30[41]}
   );
   gpc1_1 gpc3896 (
      {stage2_30[112]},
      {stage3_30[42]}
   );
   gpc1_1 gpc3897 (
      {stage2_30[113]},
      {stage3_30[43]}
   );
   gpc1_1 gpc3898 (
      {stage2_30[114]},
      {stage3_30[44]}
   );
   gpc1_1 gpc3899 (
      {stage2_30[115]},
      {stage3_30[45]}
   );
   gpc1_1 gpc3900 (
      {stage2_30[116]},
      {stage3_30[46]}
   );
   gpc1_1 gpc3901 (
      {stage2_30[117]},
      {stage3_30[47]}
   );
   gpc1_1 gpc3902 (
      {stage2_30[118]},
      {stage3_30[48]}
   );
   gpc1_1 gpc3903 (
      {stage2_30[119]},
      {stage3_30[49]}
   );
   gpc1_1 gpc3904 (
      {stage2_30[120]},
      {stage3_30[50]}
   );
   gpc1_1 gpc3905 (
      {stage2_30[121]},
      {stage3_30[51]}
   );
   gpc1_1 gpc3906 (
      {stage2_30[122]},
      {stage3_30[52]}
   );
   gpc1_1 gpc3907 (
      {stage2_30[123]},
      {stage3_30[53]}
   );
   gpc1_1 gpc3908 (
      {stage2_30[124]},
      {stage3_30[54]}
   );
   gpc1_1 gpc3909 (
      {stage2_30[125]},
      {stage3_30[55]}
   );
   gpc1_1 gpc3910 (
      {stage2_30[126]},
      {stage3_30[56]}
   );
   gpc1_1 gpc3911 (
      {stage2_30[127]},
      {stage3_30[57]}
   );
   gpc1_1 gpc3912 (
      {stage2_30[128]},
      {stage3_30[58]}
   );
   gpc1_1 gpc3913 (
      {stage2_30[129]},
      {stage3_30[59]}
   );
   gpc1_1 gpc3914 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc3915 (
      {stage2_33[36]},
      {stage3_33[30]}
   );
   gpc1_1 gpc3916 (
      {stage2_33[37]},
      {stage3_33[31]}
   );
   gpc1_1 gpc3917 (
      {stage2_33[38]},
      {stage3_33[32]}
   );
   gpc1_1 gpc3918 (
      {stage2_33[39]},
      {stage3_33[33]}
   );
   gpc1_1 gpc3919 (
      {stage2_33[40]},
      {stage3_33[34]}
   );
   gpc1_1 gpc3920 (
      {stage2_33[41]},
      {stage3_33[35]}
   );
   gpc1_1 gpc3921 (
      {stage2_33[42]},
      {stage3_33[36]}
   );
   gpc1_1 gpc3922 (
      {stage2_33[43]},
      {stage3_33[37]}
   );
   gpc1_1 gpc3923 (
      {stage2_33[44]},
      {stage3_33[38]}
   );
   gpc1_1 gpc3924 (
      {stage2_33[45]},
      {stage3_33[39]}
   );
   gpc1_1 gpc3925 (
      {stage2_34[30]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3926 (
      {stage2_34[31]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3927 (
      {stage2_34[32]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3928 (
      {stage2_34[33]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3929 (
      {stage2_34[34]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3930 (
      {stage2_34[35]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3931 (
      {stage2_35[12]},
      {stage3_35[11]}
   );
   gpc1_1 gpc3932 (
      {stage2_35[13]},
      {stage3_35[12]}
   );
   gpc606_5 gpc3933 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc3934 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc3935 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc3936 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc3937 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc3938 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc3939 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc615_5 gpc3940 (
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc3941 (
      {stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21]},
      {stage3_4[25]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[5],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc3942 (
      {stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25], stage3_3[26]},
      {stage3_4[26]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[6],stage4_5[8],stage4_4[9],stage4_3[9]}
   );
   gpc606_5 gpc3943 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[7],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc3944 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[8],stage4_5[10],stage4_4[11]}
   );
   gpc1163_5 gpc3945 (
      {stage3_5[18], stage3_5[19], stage3_5[20]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[0]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[2],stage4_7[5],stage4_6[9],stage4_5[11]}
   );
   gpc1163_5 gpc3946 (
      {stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[1]},
      {stage3_8[1]},
      {stage4_9[1],stage4_8[3],stage4_7[6],stage4_6[10],stage4_5[12]}
   );
   gpc606_5 gpc3947 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage4_9[2],stage4_8[4],stage4_7[7],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc3948 (
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage4_9[3],stage4_8[5],stage4_7[8],stage4_6[12],stage4_5[14]}
   );
   gpc606_5 gpc3949 (
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage4_9[4],stage4_8[6],stage4_7[9],stage4_6[13],stage4_5[15]}
   );
   gpc615_5 gpc3950 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[20]},
      {stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6], stage3_8[7]},
      {stage4_10[0],stage4_9[5],stage4_8[7],stage4_7[10],stage4_6[14]}
   );
   gpc615_5 gpc3951 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[21]},
      {stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13]},
      {stage4_10[1],stage4_9[6],stage4_8[8],stage4_7[11],stage4_6[15]}
   );
   gpc615_5 gpc3952 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[22]},
      {stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19]},
      {stage4_10[2],stage4_9[7],stage4_8[9],stage4_7[12],stage4_6[16]}
   );
   gpc615_5 gpc3953 (
      {stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27]},
      {stage3_8[20]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[8],stage4_8[10],stage4_7[13]}
   );
   gpc615_5 gpc3954 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[21]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[9],stage4_8[11],stage4_7[14]}
   );
   gpc615_5 gpc3955 (
      {stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36], stage3_7[37]},
      {stage3_8[22]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[10],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc3956 (
      {stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41], stage3_7[42]},
      {stage3_8[23]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[11],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc3957 (
      {stage3_7[43], stage3_7[44], stage3_7[45], stage3_7[46], stage3_7[47]},
      {stage3_8[24]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[12],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc3958 (
      {stage3_7[48], stage3_7[49], stage3_7[50], stage3_7[51], stage3_7[52]},
      {stage3_8[25]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[8],stage4_9[13],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc3959 (
      {stage3_7[53], stage3_7[54], stage3_7[55], stage3_7[56], stage3_7[57]},
      {stage3_8[26]},
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage4_11[6],stage4_10[9],stage4_9[14],stage4_8[16],stage4_7[19]}
   );
   gpc615_5 gpc3960 (
      {stage3_7[58], stage3_7[59], stage3_7[60], stage3_7[61], stage3_7[62]},
      {stage3_8[27]},
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage4_11[7],stage4_10[10],stage4_9[15],stage4_8[17],stage4_7[20]}
   );
   gpc606_5 gpc3961 (
      {stage3_8[28], stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[8],stage4_10[11],stage4_9[16],stage4_8[18]}
   );
   gpc623_5 gpc3962 (
      {stage3_9[48], stage3_9[49], stage3_9[50]},
      {stage3_10[6], stage3_10[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[9],stage4_10[12],stage4_9[17]}
   );
   gpc623_5 gpc3963 (
      {stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_10[8], stage3_10[9]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[2],stage4_11[10],stage4_10[13],stage4_9[18]}
   );
   gpc623_5 gpc3964 (
      {stage3_9[54], stage3_9[55], stage3_9[56]},
      {stage3_10[10], stage3_10[11]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[3],stage4_11[11],stage4_10[14],stage4_9[19]}
   );
   gpc623_5 gpc3965 (
      {stage3_9[57], stage3_9[58], stage3_9[59]},
      {stage3_10[12], stage3_10[13]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[4],stage4_11[12],stage4_10[15],stage4_9[20]}
   );
   gpc623_5 gpc3966 (
      {stage3_9[60], stage3_9[61], stage3_9[62]},
      {stage3_10[14], stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[5],stage4_11[13],stage4_10[16],stage4_9[21]}
   );
   gpc623_5 gpc3967 (
      {stage3_9[63], stage3_9[64], stage3_9[65]},
      {stage3_10[16], stage3_10[17]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[6],stage4_11[14],stage4_10[17],stage4_9[22]}
   );
   gpc1163_5 gpc3968 (
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[6],stage4_12[7],stage4_11[15]}
   );
   gpc606_5 gpc3969 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[7],stage4_12[8]}
   );
   gpc606_5 gpc3970 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage4_16[1],stage4_15[2],stage4_14[2],stage4_13[8],stage4_12[9]}
   );
   gpc606_5 gpc3971 (
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18]},
      {stage4_16[2],stage4_15[3],stage4_14[3],stage4_13[9],stage4_12[10]}
   );
   gpc606_5 gpc3972 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage4_16[3],stage4_15[4],stage4_14[4],stage4_13[10],stage4_12[11]}
   );
   gpc606_5 gpc3973 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage4_16[4],stage4_15[5],stage4_14[5],stage4_13[11],stage4_12[12]}
   );
   gpc606_5 gpc3974 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], stage3_14[36]},
      {stage4_16[5],stage4_15[6],stage4_14[6],stage4_13[12],stage4_12[13]}
   );
   gpc2135_5 gpc3975 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[37], stage3_14[38], stage3_14[39]},
      {stage3_15[0]},
      {stage3_16[0], stage3_16[1]},
      {stage4_17[0],stage4_16[6],stage4_15[7],stage4_14[7],stage4_13[13]}
   );
   gpc2135_5 gpc3976 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[40], stage3_14[41], stage3_14[42]},
      {stage3_15[1]},
      {stage3_16[2], stage3_16[3]},
      {stage4_17[1],stage4_16[7],stage4_15[8],stage4_14[8],stage4_13[14]}
   );
   gpc2135_5 gpc3977 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[43], stage3_14[44], stage3_14[45]},
      {stage3_15[2]},
      {stage3_16[4], stage3_16[5]},
      {stage4_17[2],stage4_16[8],stage4_15[9],stage4_14[9],stage4_13[15]}
   );
   gpc2135_5 gpc3978 (
      {stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_14[46], stage3_14[47], stage3_14[48]},
      {stage3_15[3]},
      {stage3_16[6], stage3_16[7]},
      {stage4_17[3],stage4_16[9],stage4_15[10],stage4_14[10],stage4_13[16]}
   );
   gpc2135_5 gpc3979 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_14[49], stage3_14[50], 1'b0},
      {stage3_15[4]},
      {stage3_16[8], stage3_16[9]},
      {stage4_17[4],stage4_16[10],stage4_15[11],stage4_14[11],stage4_13[17]}
   );
   gpc606_5 gpc3980 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10]},
      {stage4_17[5],stage4_16[11],stage4_15[12],stage4_14[12],stage4_13[18]}
   );
   gpc2135_5 gpc3981 (
      {stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage3_16[10], stage3_16[11], stage3_16[12]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[6],stage4_16[12],stage4_15[13]}
   );
   gpc2135_5 gpc3982 (
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage3_17[1]},
      {stage3_18[2], stage3_18[3]},
      {stage4_19[1],stage4_18[1],stage4_17[7],stage4_16[13],stage4_15[14]}
   );
   gpc2135_5 gpc3983 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[2]},
      {stage3_18[4], stage3_18[5]},
      {stage4_19[2],stage4_18[2],stage4_17[8],stage4_16[14],stage4_15[15]}
   );
   gpc2135_5 gpc3984 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[19], stage3_16[20], stage3_16[21]},
      {stage3_17[3]},
      {stage3_18[6], stage3_18[7]},
      {stage4_19[3],stage4_18[3],stage4_17[9],stage4_16[15],stage4_15[16]}
   );
   gpc2135_5 gpc3985 (
      {stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage3_16[22], stage3_16[23], stage3_16[24]},
      {stage3_17[4]},
      {stage3_18[8], stage3_18[9]},
      {stage4_19[4],stage4_18[4],stage4_17[10],stage4_16[16],stage4_15[17]}
   );
   gpc2135_5 gpc3986 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40]},
      {stage3_16[25], stage3_16[26], stage3_16[27]},
      {stage3_17[5]},
      {stage3_18[10], stage3_18[11]},
      {stage4_19[5],stage4_18[5],stage4_17[11],stage4_16[17],stage4_15[18]}
   );
   gpc2135_5 gpc3987 (
      {stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45]},
      {stage3_16[28], stage3_16[29], stage3_16[30]},
      {stage3_17[6]},
      {stage3_18[12], stage3_18[13]},
      {stage4_19[6],stage4_18[6],stage4_17[12],stage4_16[18],stage4_15[19]}
   );
   gpc2135_5 gpc3988 (
      {stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49], stage3_15[50]},
      {stage3_16[31], stage3_16[32], stage3_16[33]},
      {stage3_17[7]},
      {stage3_18[14], stage3_18[15]},
      {stage4_19[7],stage4_18[7],stage4_17[13],stage4_16[19],stage4_15[20]}
   );
   gpc2135_5 gpc3989 (
      {stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54], stage3_15[55]},
      {stage3_16[34], stage3_16[35], stage3_16[36]},
      {stage3_17[8]},
      {stage3_18[16], stage3_18[17]},
      {stage4_19[8],stage4_18[8],stage4_17[14],stage4_16[20],stage4_15[21]}
   );
   gpc2135_5 gpc3990 (
      {stage3_15[56], stage3_15[57], stage3_15[58], stage3_15[59], stage3_15[60]},
      {stage3_16[37], stage3_16[38], stage3_16[39]},
      {stage3_17[9]},
      {stage3_18[18], stage3_18[19]},
      {stage4_19[9],stage4_18[9],stage4_17[15],stage4_16[21],stage4_15[22]}
   );
   gpc615_5 gpc3991 (
      {stage3_15[61], stage3_15[62], stage3_15[63], stage3_15[64], stage3_15[65]},
      {stage3_16[40]},
      {stage3_17[10], stage3_17[11], stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15]},
      {stage4_19[10],stage4_18[10],stage4_17[16],stage4_16[22],stage4_15[23]}
   );
   gpc606_5 gpc3992 (
      {stage3_16[41], stage3_16[42], stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46]},
      {stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage4_20[0],stage4_19[11],stage4_18[11],stage4_17[17],stage4_16[23]}
   );
   gpc606_5 gpc3993 (
      {stage3_16[47], stage3_16[48], stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52]},
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31]},
      {stage4_20[1],stage4_19[12],stage4_18[12],stage4_17[18],stage4_16[24]}
   );
   gpc606_5 gpc3994 (
      {stage3_16[53], stage3_16[54], stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58]},
      {stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35], stage3_18[36], stage3_18[37]},
      {stage4_20[2],stage4_19[13],stage4_18[13],stage4_17[19],stage4_16[25]}
   );
   gpc1163_5 gpc3995 (
      {stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41], stage3_18[42], stage3_18[43]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[3],stage4_19[14],stage4_18[14],stage4_17[20]}
   );
   gpc1163_5 gpc3996 (
      {stage3_17[19], stage3_17[20], stage3_17[21]},
      {stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48], stage3_18[49]},
      {stage3_19[1]},
      {stage3_20[1]},
      {stage4_21[1],stage4_20[4],stage4_19[15],stage4_18[15],stage4_17[21]}
   );
   gpc606_5 gpc3997 (
      {stage3_17[22], stage3_17[23], stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27]},
      {stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6], stage3_19[7]},
      {stage4_21[2],stage4_20[5],stage4_19[16],stage4_18[16],stage4_17[22]}
   );
   gpc606_5 gpc3998 (
      {stage3_17[28], stage3_17[29], stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33]},
      {stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11], stage3_19[12], stage3_19[13]},
      {stage4_21[3],stage4_20[6],stage4_19[17],stage4_18[17],stage4_17[23]}
   );
   gpc606_5 gpc3999 (
      {stage3_17[34], stage3_17[35], stage3_17[36], stage3_17[37], stage3_17[38], stage3_17[39]},
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage4_21[4],stage4_20[7],stage4_19[18],stage4_18[18],stage4_17[24]}
   );
   gpc615_5 gpc4000 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24]},
      {stage3_20[2]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[5],stage4_20[8],stage4_19[19]}
   );
   gpc615_5 gpc4001 (
      {stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage3_20[3]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[6],stage4_20[9],stage4_19[20]}
   );
   gpc615_5 gpc4002 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[4]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[7],stage4_20[10],stage4_19[21]}
   );
   gpc615_5 gpc4003 (
      {stage3_19[35], stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39]},
      {stage3_20[5]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[8],stage4_20[11],stage4_19[22]}
   );
   gpc1325_5 gpc4004 (
      {stage3_19[40], stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44]},
      {stage3_20[6], stage3_20[7]},
      {stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_22[0]},
      {stage4_23[4],stage4_22[4],stage4_21[9],stage4_20[12],stage4_19[23]}
   );
   gpc1406_5 gpc4005 (
      {stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4]},
      {stage3_23[0]},
      {stage4_24[0],stage4_23[5],stage4_22[5],stage4_21[10],stage4_20[13]}
   );
   gpc606_5 gpc4006 (
      {stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19]},
      {stage3_22[5], stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage4_24[1],stage4_23[6],stage4_22[6],stage4_21[11],stage4_20[14]}
   );
   gpc606_5 gpc4007 (
      {stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24], stage3_20[25]},
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage4_24[2],stage4_23[7],stage4_22[7],stage4_21[12],stage4_20[15]}
   );
   gpc606_5 gpc4008 (
      {stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31]},
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22]},
      {stage4_24[3],stage4_23[8],stage4_22[8],stage4_21[13],stage4_20[16]}
   );
   gpc606_5 gpc4009 (
      {stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37]},
      {stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28]},
      {stage4_24[4],stage4_23[9],stage4_22[9],stage4_21[14],stage4_20[17]}
   );
   gpc606_5 gpc4010 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage4_25[0],stage4_24[5],stage4_23[10],stage4_22[10],stage4_21[15]}
   );
   gpc606_5 gpc4011 (
      {stage3_21[33], stage3_21[34], stage3_21[35], stage3_21[36], stage3_21[37], stage3_21[38]},
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12]},
      {stage4_25[1],stage4_24[6],stage4_23[11],stage4_22[11],stage4_21[16]}
   );
   gpc606_5 gpc4012 (
      {stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42], stage3_21[43], stage3_21[44]},
      {stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage4_25[2],stage4_24[7],stage4_23[12],stage4_22[12],stage4_21[17]}
   );
   gpc606_5 gpc4013 (
      {stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23], stage3_23[24]},
      {stage4_25[3],stage4_24[8],stage4_23[13],stage4_22[13],stage4_21[18]}
   );
   gpc606_5 gpc4014 (
      {stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54], stage3_21[55], stage3_21[56]},
      {stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28], stage3_23[29], stage3_23[30]},
      {stage4_25[4],stage4_24[9],stage4_23[14],stage4_22[14],stage4_21[19]}
   );
   gpc606_5 gpc4015 (
      {stage3_22[29], stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[5],stage4_24[10],stage4_23[15],stage4_22[15]}
   );
   gpc606_5 gpc4016 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[6],stage4_24[11],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc4017 (
      {stage3_23[31], stage3_23[32], stage3_23[33], stage3_23[34], stage3_23[35]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[7],stage4_24[12],stage4_23[17]}
   );
   gpc615_5 gpc4018 (
      {stage3_23[36], stage3_23[37], stage3_23[38], stage3_23[39], stage3_23[40]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[8],stage4_24[13],stage4_23[18]}
   );
   gpc615_5 gpc4019 (
      {stage3_23[41], stage3_23[42], stage3_23[43], stage3_23[44], stage3_23[45]},
      {stage3_24[14]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[9],stage4_24[14],stage4_23[19]}
   );
   gpc606_5 gpc4020 (
      {stage3_24[15], stage3_24[16], stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[3],stage4_26[5],stage4_25[10],stage4_24[15]}
   );
   gpc606_5 gpc4021 (
      {stage3_24[21], stage3_24[22], stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[4],stage4_26[6],stage4_25[11],stage4_24[16]}
   );
   gpc606_5 gpc4022 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[2],stage4_27[5],stage4_26[7],stage4_25[12]}
   );
   gpc615_5 gpc4023 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28]},
      {stage3_26[12]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[3],stage4_27[6],stage4_26[8],stage4_25[13]}
   );
   gpc615_5 gpc4024 (
      {stage3_25[29], stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33]},
      {stage3_26[13]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[4],stage4_27[7],stage4_26[9],stage4_25[14]}
   );
   gpc615_5 gpc4025 (
      {stage3_25[34], stage3_25[35], stage3_25[36], stage3_25[37], stage3_25[38]},
      {stage3_26[14]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[5],stage4_27[8],stage4_26[10],stage4_25[15]}
   );
   gpc615_5 gpc4026 (
      {stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18], stage3_26[19]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[6],stage4_27[9],stage4_26[11]}
   );
   gpc606_5 gpc4027 (
      {stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[1],stage4_29[5],stage4_28[7],stage4_27[10]}
   );
   gpc606_5 gpc4028 (
      {stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[2],stage4_29[6],stage4_28[8],stage4_27[11]}
   );
   gpc606_5 gpc4029 (
      {stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[3],stage4_29[7],stage4_28[9],stage4_27[12]}
   );
   gpc606_5 gpc4030 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47], stage3_27[48]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[4],stage4_29[8],stage4_28[10],stage4_27[13]}
   );
   gpc615_5 gpc4031 (
      {stage3_27[49], stage3_27[50], stage3_27[51], stage3_27[52], stage3_27[53]},
      {stage3_28[6]},
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage4_31[4],stage4_30[5],stage4_29[9],stage4_28[11],stage4_27[14]}
   );
   gpc606_5 gpc4032 (
      {stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[5],stage4_30[6],stage4_29[10],stage4_28[12]}
   );
   gpc606_5 gpc4033 (
      {stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[6],stage4_30[7],stage4_29[11],stage4_28[13]}
   );
   gpc606_5 gpc4034 (
      {stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[7],stage4_30[8],stage4_29[12],stage4_28[14]}
   );
   gpc606_5 gpc4035 (
      {stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[8],stage4_30[9],stage4_29[13],stage4_28[15]}
   );
   gpc606_5 gpc4036 (
      {stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[9],stage4_30[10],stage4_29[14],stage4_28[16]}
   );
   gpc606_5 gpc4037 (
      {stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[10],stage4_30[11],stage4_29[15],stage4_28[17]}
   );
   gpc615_5 gpc4038 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34]},
      {stage3_30[36]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[6],stage4_31[11],stage4_30[12],stage4_29[16]}
   );
   gpc606_5 gpc4039 (
      {stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41], stage3_30[42]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[7],stage4_31[12],stage4_30[13]}
   );
   gpc615_5 gpc4040 (
      {stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage3_31[6]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[2],stage4_32[8],stage4_31[13],stage4_30[14]}
   );
   gpc615_5 gpc4041 (
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52]},
      {stage3_31[7]},
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage4_34[2],stage4_33[3],stage4_32[9],stage4_31[14],stage4_30[15]}
   );
   gpc606_5 gpc4042 (
      {stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[3],stage4_33[4],stage4_32[10],stage4_31[15]}
   );
   gpc606_5 gpc4043 (
      {stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[4],stage4_33[5],stage4_32[11],stage4_31[16]}
   );
   gpc615_5 gpc4044 (
      {stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23], stage3_31[24]},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[5],stage4_33[6],stage4_32[12],stage4_31[17]}
   );
   gpc615_5 gpc4045 (
      {stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage3_32[19]},
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage4_35[3],stage4_34[6],stage4_33[7],stage4_32[13],stage4_31[18]}
   );
   gpc615_5 gpc4046 (
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34]},
      {stage3_32[20]},
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29]},
      {stage4_35[4],stage4_34[7],stage4_33[8],stage4_32[14],stage4_31[19]}
   );
   gpc1325_5 gpc4047 (
      {stage3_31[35], stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39]},
      {stage3_32[21], stage3_32[22]},
      {stage3_33[30], stage3_33[31], stage3_33[32]},
      {stage3_34[0]},
      {stage4_35[5],stage4_34[8],stage4_33[9],stage4_32[15],stage4_31[20]}
   );
   gpc606_5 gpc4048 (
      {stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28]},
      {stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6]},
      {stage4_36[0],stage4_35[6],stage4_34[9],stage4_33[10],stage4_32[16]}
   );
   gpc606_5 gpc4049 (
      {stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34]},
      {stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12]},
      {stage4_36[1],stage4_35[7],stage4_34[10],stage4_33[11],stage4_32[17]}
   );
   gpc606_5 gpc4050 (
      {stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[8],stage4_34[11],stage4_33[12]}
   );
   gpc2135_5 gpc4051 (
      {stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage3_35[6], stage3_35[7], stage3_35[8]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1]},
      {stage4_38[0],stage4_37[1],stage4_36[3],stage4_35[9],stage4_34[12]}
   );
   gpc1_1 gpc4052 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4053 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4054 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4055 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4056 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4057 (
      {stage3_1[15]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4058 (
      {stage3_1[16]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4059 (
      {stage3_1[17]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4060 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4061 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4062 (
      {stage3_4[39]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4063 (
      {stage3_4[40]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4064 (
      {stage3_4[41]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4065 (
      {stage3_4[42]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4066 (
      {stage3_4[43]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4067 (
      {stage3_5[42]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4068 (
      {stage3_5[43]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4069 (
      {stage3_5[44]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4070 (
      {stage3_5[45]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4071 (
      {stage3_5[46]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4072 (
      {stage3_5[47]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4073 (
      {stage3_5[48]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4074 (
      {stage3_6[39]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4075 (
      {stage3_6[40]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4076 (
      {stage3_6[41]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4077 (
      {stage3_6[42]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4078 (
      {stage3_7[63]},
      {stage4_7[21]}
   );
   gpc1_1 gpc4079 (
      {stage3_7[64]},
      {stage4_7[22]}
   );
   gpc1_1 gpc4080 (
      {stage3_7[65]},
      {stage4_7[23]}
   );
   gpc1_1 gpc4081 (
      {stage3_7[66]},
      {stage4_7[24]}
   );
   gpc1_1 gpc4082 (
      {stage3_7[67]},
      {stage4_7[25]}
   );
   gpc1_1 gpc4083 (
      {stage3_7[68]},
      {stage4_7[26]}
   );
   gpc1_1 gpc4084 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc4085 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc4086 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4087 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4088 (
      {stage3_9[66]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4089 (
      {stage3_9[67]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4090 (
      {stage3_9[68]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4091 (
      {stage3_9[69]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4092 (
      {stage3_10[18]},
      {stage4_10[18]}
   );
   gpc1_1 gpc4093 (
      {stage3_10[19]},
      {stage4_10[19]}
   );
   gpc1_1 gpc4094 (
      {stage3_10[20]},
      {stage4_10[20]}
   );
   gpc1_1 gpc4095 (
      {stage3_10[21]},
      {stage4_10[21]}
   );
   gpc1_1 gpc4096 (
      {stage3_10[22]},
      {stage4_10[22]}
   );
   gpc1_1 gpc4097 (
      {stage3_10[23]},
      {stage4_10[23]}
   );
   gpc1_1 gpc4098 (
      {stage3_10[24]},
      {stage4_10[24]}
   );
   gpc1_1 gpc4099 (
      {stage3_10[25]},
      {stage4_10[25]}
   );
   gpc1_1 gpc4100 (
      {stage3_10[26]},
      {stage4_10[26]}
   );
   gpc1_1 gpc4101 (
      {stage3_10[27]},
      {stage4_10[27]}
   );
   gpc1_1 gpc4102 (
      {stage3_10[28]},
      {stage4_10[28]}
   );
   gpc1_1 gpc4103 (
      {stage3_11[39]},
      {stage4_11[16]}
   );
   gpc1_1 gpc4104 (
      {stage3_11[40]},
      {stage4_11[17]}
   );
   gpc1_1 gpc4105 (
      {stage3_11[41]},
      {stage4_11[18]}
   );
   gpc1_1 gpc4106 (
      {stage3_11[42]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4107 (
      {stage3_11[43]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4108 (
      {stage3_13[32]},
      {stage4_13[19]}
   );
   gpc1_1 gpc4109 (
      {stage3_13[33]},
      {stage4_13[20]}
   );
   gpc1_1 gpc4110 (
      {stage3_13[34]},
      {stage4_13[21]}
   );
   gpc1_1 gpc4111 (
      {stage3_13[35]},
      {stage4_13[22]}
   );
   gpc1_1 gpc4112 (
      {stage3_13[36]},
      {stage4_13[23]}
   );
   gpc1_1 gpc4113 (
      {stage3_13[37]},
      {stage4_13[24]}
   );
   gpc1_1 gpc4114 (
      {stage3_13[38]},
      {stage4_13[25]}
   );
   gpc1_1 gpc4115 (
      {stage3_13[39]},
      {stage4_13[26]}
   );
   gpc1_1 gpc4116 (
      {stage3_13[40]},
      {stage4_13[27]}
   );
   gpc1_1 gpc4117 (
      {stage3_15[66]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4118 (
      {stage3_15[67]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4119 (
      {stage3_15[68]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4120 (
      {stage3_15[69]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4121 (
      {stage3_15[70]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4122 (
      {stage3_15[71]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4123 (
      {stage3_15[72]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4124 (
      {stage3_15[73]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4125 (
      {stage3_15[74]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4126 (
      {stage3_15[75]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4127 (
      {stage3_15[76]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4128 (
      {stage3_15[77]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4129 (
      {stage3_15[78]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4130 (
      {stage3_15[79]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4131 (
      {stage3_15[80]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4132 (
      {stage3_15[81]},
      {stage4_15[39]}
   );
   gpc1_1 gpc4133 (
      {stage3_15[82]},
      {stage4_15[40]}
   );
   gpc1_1 gpc4134 (
      {stage3_15[83]},
      {stage4_15[41]}
   );
   gpc1_1 gpc4135 (
      {stage3_15[84]},
      {stage4_15[42]}
   );
   gpc1_1 gpc4136 (
      {stage3_15[85]},
      {stage4_15[43]}
   );
   gpc1_1 gpc4137 (
      {stage3_15[86]},
      {stage4_15[44]}
   );
   gpc1_1 gpc4138 (
      {stage3_15[87]},
      {stage4_15[45]}
   );
   gpc1_1 gpc4139 (
      {stage3_15[88]},
      {stage4_15[46]}
   );
   gpc1_1 gpc4140 (
      {stage3_15[89]},
      {stage4_15[47]}
   );
   gpc1_1 gpc4141 (
      {stage3_16[59]},
      {stage4_16[26]}
   );
   gpc1_1 gpc4142 (
      {stage3_16[60]},
      {stage4_16[27]}
   );
   gpc1_1 gpc4143 (
      {stage3_16[61]},
      {stage4_16[28]}
   );
   gpc1_1 gpc4144 (
      {stage3_17[40]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4145 (
      {stage3_17[41]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4146 (
      {stage3_17[42]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4147 (
      {stage3_17[43]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4148 (
      {stage3_17[44]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4149 (
      {stage3_17[45]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4150 (
      {stage3_17[46]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4151 (
      {stage3_17[47]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4152 (
      {stage3_17[48]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4153 (
      {stage3_17[49]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4154 (
      {stage3_19[45]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4155 (
      {stage3_19[46]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4156 (
      {stage3_19[47]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4157 (
      {stage3_19[48]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4158 (
      {stage3_19[49]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4159 (
      {stage3_20[38]},
      {stage4_20[18]}
   );
   gpc1_1 gpc4160 (
      {stage3_20[39]},
      {stage4_20[19]}
   );
   gpc1_1 gpc4161 (
      {stage3_20[40]},
      {stage4_20[20]}
   );
   gpc1_1 gpc4162 (
      {stage3_20[41]},
      {stage4_20[21]}
   );
   gpc1_1 gpc4163 (
      {stage3_20[42]},
      {stage4_20[22]}
   );
   gpc1_1 gpc4164 (
      {stage3_20[43]},
      {stage4_20[23]}
   );
   gpc1_1 gpc4165 (
      {stage3_20[44]},
      {stage4_20[24]}
   );
   gpc1_1 gpc4166 (
      {stage3_20[45]},
      {stage4_20[25]}
   );
   gpc1_1 gpc4167 (
      {stage3_21[57]},
      {stage4_21[20]}
   );
   gpc1_1 gpc4168 (
      {stage3_21[58]},
      {stage4_21[21]}
   );
   gpc1_1 gpc4169 (
      {stage3_22[41]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4170 (
      {stage3_22[42]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4171 (
      {stage3_22[43]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4172 (
      {stage3_22[44]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4173 (
      {stage3_22[45]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4174 (
      {stage3_22[46]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4175 (
      {stage3_23[46]},
      {stage4_23[20]}
   );
   gpc1_1 gpc4176 (
      {stage3_23[47]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4177 (
      {stage3_24[27]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4178 (
      {stage3_24[28]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4179 (
      {stage3_24[29]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4180 (
      {stage3_24[30]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4181 (
      {stage3_24[31]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4182 (
      {stage3_24[32]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4183 (
      {stage3_24[33]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4184 (
      {stage3_24[34]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4185 (
      {stage3_24[35]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4186 (
      {stage3_24[36]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4187 (
      {stage3_24[37]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4188 (
      {stage3_24[38]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4189 (
      {stage3_24[39]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4190 (
      {stage3_24[40]},
      {stage4_24[30]}
   );
   gpc1_1 gpc4191 (
      {stage3_25[39]},
      {stage4_25[16]}
   );
   gpc1_1 gpc4192 (
      {stage3_26[20]},
      {stage4_26[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_26[21]},
      {stage4_26[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_26[24]},
      {stage4_26[16]}
   );
   gpc1_1 gpc4197 (
      {stage3_26[25]},
      {stage4_26[17]}
   );
   gpc1_1 gpc4198 (
      {stage3_26[26]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4199 (
      {stage3_26[27]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4200 (
      {stage3_26[28]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4201 (
      {stage3_26[29]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4202 (
      {stage3_26[30]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4203 (
      {stage3_26[31]},
      {stage4_26[23]}
   );
   gpc1_1 gpc4204 (
      {stage3_27[54]},
      {stage4_27[15]}
   );
   gpc1_1 gpc4205 (
      {stage3_27[55]},
      {stage4_27[16]}
   );
   gpc1_1 gpc4206 (
      {stage3_27[56]},
      {stage4_27[17]}
   );
   gpc1_1 gpc4207 (
      {stage3_27[57]},
      {stage4_27[18]}
   );
   gpc1_1 gpc4208 (
      {stage3_27[58]},
      {stage4_27[19]}
   );
   gpc1_1 gpc4209 (
      {stage3_27[59]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4210 (
      {stage3_27[60]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4211 (
      {stage3_27[61]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4212 (
      {stage3_27[62]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4213 (
      {stage3_27[63]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4214 (
      {stage3_27[64]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4215 (
      {stage3_27[65]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4216 (
      {stage3_27[66]},
      {stage4_27[27]}
   );
   gpc1_1 gpc4217 (
      {stage3_29[35]},
      {stage4_29[17]}
   );
   gpc1_1 gpc4218 (
      {stage3_29[36]},
      {stage4_29[18]}
   );
   gpc1_1 gpc4219 (
      {stage3_29[37]},
      {stage4_29[19]}
   );
   gpc1_1 gpc4220 (
      {stage3_29[38]},
      {stage4_29[20]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[53]},
      {stage4_30[16]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[54]},
      {stage4_30[17]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[55]},
      {stage4_30[18]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[56]},
      {stage4_30[19]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[57]},
      {stage4_30[20]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[58]},
      {stage4_30[21]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[59]},
      {stage4_30[22]}
   );
   gpc1_1 gpc4228 (
      {stage3_32[35]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4229 (
      {stage3_33[39]},
      {stage4_33[13]}
   );
   gpc1_1 gpc4230 (
      {stage3_34[18]},
      {stage4_34[13]}
   );
   gpc1_1 gpc4231 (
      {stage3_34[19]},
      {stage4_34[14]}
   );
   gpc1_1 gpc4232 (
      {stage3_34[20]},
      {stage4_34[15]}
   );
   gpc1_1 gpc4233 (
      {stage3_34[21]},
      {stage4_34[16]}
   );
   gpc1_1 gpc4234 (
      {stage3_35[9]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4235 (
      {stage3_35[10]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4236 (
      {stage3_35[11]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4237 (
      {stage3_35[12]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4238 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc4239 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4240 (
      {stage3_36[3]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4241 (
      {stage3_36[4]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4242 (
      {stage3_36[5]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4243 (
      {stage3_36[6]},
      {stage4_36[9]}
   );
   gpc615_5 gpc4244 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc1343_5 gpc4245 (
      {stage4_3[1], stage4_3[2], stage4_3[3]},
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc606_5 gpc4246 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc1415_5 gpc4247 (
      {stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_6[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc606_5 gpc4248 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9]},
      {stage5_9[1],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc4249 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15]},
      {stage5_9[2],stage5_8[3],stage5_7[4],stage5_6[5],stage5_5[5]}
   );
   gpc606_5 gpc4250 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13]},
      {stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[5],stage5_6[6]}
   );
   gpc615_5 gpc4251 (
      {stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage4_7[16]},
      {stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage5_10[1],stage5_9[4],stage5_8[5],stage5_7[6],stage5_6[7]}
   );
   gpc1343_5 gpc4252 (
      {stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[5],stage5_8[6],stage5_7[7]}
   );
   gpc615_5 gpc4253 (
      {stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage4_8[17]},
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8]},
      {stage5_11[1],stage5_10[3],stage5_9[6],stage5_8[7],stage5_7[8]}
   );
   gpc606_5 gpc4254 (
      {stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[7]}
   );
   gpc615_5 gpc4255 (
      {stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18], stage4_9[19]},
      {stage4_10[1]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[8]}
   );
   gpc615_5 gpc4256 (
      {stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_10[2]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[9]}
   );
   gpc207_4 gpc4257 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc615_5 gpc4258 (
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14]},
      {stage4_11[18]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[4],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc1163_5 gpc4259 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[5]}
   );
   gpc606_5 gpc4260 (
      {stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[6]}
   );
   gpc606_5 gpc4261 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12]},
      {stage5_17[2],stage5_16[2],stage5_15[2],stage5_14[3],stage5_13[7]}
   );
   gpc606_5 gpc4262 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19], stage4_13[20]},
      {stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage5_17[3],stage5_16[3],stage5_15[3],stage5_14[4],stage5_13[8]}
   );
   gpc615_5 gpc4263 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[19]},
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage5_18[0],stage5_17[4],stage5_16[4],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc4264 (
      {stage4_15[20], stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26]},
      {stage4_17[0], stage4_17[1]},
      {stage5_18[1],stage5_17[5],stage5_16[5],stage5_15[5]}
   );
   gpc615_5 gpc4265 (
      {stage4_15[27], stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31]},
      {stage4_16[7]},
      {stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6], stage4_17[7]},
      {stage5_19[0],stage5_18[2],stage5_17[6],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc4266 (
      {stage4_15[32], stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36]},
      {stage4_16[8]},
      {stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12], stage4_17[13]},
      {stage5_19[1],stage5_18[3],stage5_17[7],stage5_16[7],stage5_15[7]}
   );
   gpc615_5 gpc4267 (
      {stage4_15[37], stage4_15[38], stage4_15[39], stage4_15[40], stage4_15[41]},
      {stage4_16[9]},
      {stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17], stage4_17[18], stage4_17[19]},
      {stage5_19[2],stage5_18[4],stage5_17[8],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4268 (
      {stage4_15[42], stage4_15[43], stage4_15[44], stage4_15[45], stage4_15[46]},
      {stage4_16[10]},
      {stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23], stage4_17[24], stage4_17[25]},
      {stage5_19[3],stage5_18[5],stage5_17[9],stage5_16[9],stage5_15[9]}
   );
   gpc207_4 gpc4269 (
      {stage4_16[11], stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[4],stage5_18[6],stage5_17[10],stage5_16[10]}
   );
   gpc606_5 gpc4270 (
      {stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30], stage4_17[31]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[5],stage5_18[7],stage5_17[11]}
   );
   gpc615_5 gpc4271 (
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[6],stage5_18[8]}
   );
   gpc615_5 gpc4272 (
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[7],stage5_18[9]}
   );
   gpc615_5 gpc4273 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16]},
      {stage4_19[8]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[8],stage5_18[10]}
   );
   gpc2135_5 gpc4274 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage4_21[0]},
      {stage4_22[0], stage4_22[1]},
      {stage5_23[0],stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[9]}
   );
   gpc615_5 gpc4275 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[21]},
      {stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[10]}
   );
   gpc615_5 gpc4276 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[22]},
      {stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11], stage4_21[12]},
      {stage5_23[2],stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[11]}
   );
   gpc615_5 gpc4277 (
      {stage4_19[24], stage4_19[25], stage4_19[26], stage4_19[27], stage4_19[28]},
      {stage4_20[23]},
      {stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[3],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[12]}
   );
   gpc615_5 gpc4278 (
      {stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[7]}
   );
   gpc615_5 gpc4279 (
      {stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage4_23[1]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[8]}
   );
   gpc615_5 gpc4280 (
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16]},
      {stage4_23[2]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[9]}
   );
   gpc615_5 gpc4281 (
      {stage4_22[17], stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21]},
      {stage4_23[3]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[10]}
   );
   gpc615_5 gpc4282 (
      {stage4_23[4], stage4_23[5], stage4_23[6], stage4_23[7], stage4_23[8]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[8]}
   );
   gpc615_5 gpc4283 (
      {stage4_23[9], stage4_23[10], stage4_23[11], stage4_23[12], stage4_23[13]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[9]}
   );
   gpc615_5 gpc4284 (
      {stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17], stage4_23[18]},
      {stage4_24[26]},
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], 1'b0},
      {stage5_27[2],stage5_26[6],stage5_25[6],stage5_24[6],stage5_23[10]}
   );
   gpc606_5 gpc4285 (
      {stage4_24[27], stage4_24[28], stage4_24[29], stage4_24[30], 1'b0, 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[3],stage5_26[7],stage5_25[7],stage5_24[7]}
   );
   gpc615_5 gpc4286 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4287 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4288 (
      {stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19], stage4_26[20]},
      {stage4_27[2]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[3],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4289 (
      {stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[3],stage5_29[3],stage5_28[4],stage5_27[7]}
   );
   gpc207_4 gpc4290 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[2], stage4_29[3]},
      {stage5_30[4],stage5_29[4],stage5_28[5],stage5_27[8]}
   );
   gpc207_4 gpc4291 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage4_29[4], stage4_29[5]},
      {stage5_30[5],stage5_29[5],stage5_28[6],stage5_27[9]}
   );
   gpc615_5 gpc4292 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[6],stage5_29[6]}
   );
   gpc615_5 gpc4293 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[7],stage5_29[7]}
   );
   gpc117_4 gpc4294 (
      {stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7], stage4_30[8]},
      {stage4_31[12]},
      {stage4_32[0]},
      {stage5_33[2],stage5_32[2],stage5_31[2],stage5_30[8]}
   );
   gpc117_4 gpc4295 (
      {stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15]},
      {stage4_31[13]},
      {stage4_32[1]},
      {stage5_33[3],stage5_32[3],stage5_31[3],stage5_30[9]}
   );
   gpc615_5 gpc4296 (
      {stage4_30[16], stage4_30[17], stage4_30[18], stage4_30[19], stage4_30[20]},
      {stage4_31[14]},
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage5_34[0],stage5_33[4],stage5_32[4],stage5_31[4],stage5_30[10]}
   );
   gpc615_5 gpc4297 (
      {stage4_30[21], stage4_30[22], 1'b0, 1'b0, 1'b0},
      {stage4_31[15]},
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage5_34[1],stage5_33[5],stage5_32[5],stage5_31[5],stage5_30[11]}
   );
   gpc2135_5 gpc4298 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4]},
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage4_35[0]},
      {stage4_36[0], stage4_36[1]},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[6]}
   );
   gpc2135_5 gpc4299 (
      {stage4_33[5], stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9]},
      {stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_35[1]},
      {stage4_36[2], stage4_36[3]},
      {stage5_37[1],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[7]}
   );
   gpc2135_5 gpc4300 (
      {stage4_33[10], stage4_33[11], stage4_33[12], stage4_33[13], 1'b0},
      {stage4_34[6], stage4_34[7], stage4_34[8]},
      {stage4_35[2]},
      {stage4_36[4], stage4_36[5]},
      {stage5_37[2],stage5_36[2],stage5_35[2],stage5_34[4],stage5_33[8]}
   );
   gpc606_5 gpc4301 (
      {stage4_34[9], stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], 1'b0, 1'b0},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[3],stage5_34[5]}
   );
   gpc1_1 gpc4302 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4303 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4304 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4305 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc4306 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4307 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4308 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4309 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4310 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4311 (
      {stage4_1[6]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4312 (
      {stage4_1[7]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4313 (
      {stage4_1[8]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4314 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4315 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4316 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4317 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4318 (
      {stage4_3[4]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4319 (
      {stage4_3[5]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4320 (
      {stage4_3[6]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4321 (
      {stage4_3[7]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4322 (
      {stage4_3[8]},
      {stage5_3[6]}
   );
   gpc1_1 gpc4323 (
      {stage4_3[9]},
      {stage5_3[7]}
   );
   gpc1_1 gpc4324 (
      {stage4_4[16]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4325 (
      {stage4_5[20]},
      {stage5_5[6]}
   );
   gpc1_1 gpc4326 (
      {stage4_5[21]},
      {stage5_5[7]}
   );
   gpc1_1 gpc4327 (
      {stage4_5[22]},
      {stage5_5[8]}
   );
   gpc1_1 gpc4328 (
      {stage4_6[19]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4329 (
      {stage4_6[20]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4330 (
      {stage4_7[25]},
      {stage5_7[9]}
   );
   gpc1_1 gpc4331 (
      {stage4_7[26]},
      {stage5_7[10]}
   );
   gpc1_1 gpc4332 (
      {stage4_8[18]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4333 (
      {stage4_8[19]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4334 (
      {stage4_8[20]},
      {stage5_8[10]}
   );
   gpc1_1 gpc4335 (
      {stage4_8[21]},
      {stage5_8[11]}
   );
   gpc1_1 gpc4336 (
      {stage4_8[22]},
      {stage5_8[12]}
   );
   gpc1_1 gpc4337 (
      {stage4_9[25]},
      {stage5_9[10]}
   );
   gpc1_1 gpc4338 (
      {stage4_9[26]},
      {stage5_9[11]}
   );
   gpc1_1 gpc4339 (
      {stage4_10[15]},
      {stage5_10[9]}
   );
   gpc1_1 gpc4340 (
      {stage4_10[16]},
      {stage5_10[10]}
   );
   gpc1_1 gpc4341 (
      {stage4_10[17]},
      {stage5_10[11]}
   );
   gpc1_1 gpc4342 (
      {stage4_10[18]},
      {stage5_10[12]}
   );
   gpc1_1 gpc4343 (
      {stage4_10[19]},
      {stage5_10[13]}
   );
   gpc1_1 gpc4344 (
      {stage4_10[20]},
      {stage5_10[14]}
   );
   gpc1_1 gpc4345 (
      {stage4_10[21]},
      {stage5_10[15]}
   );
   gpc1_1 gpc4346 (
      {stage4_10[22]},
      {stage5_10[16]}
   );
   gpc1_1 gpc4347 (
      {stage4_10[23]},
      {stage5_10[17]}
   );
   gpc1_1 gpc4348 (
      {stage4_10[24]},
      {stage5_10[18]}
   );
   gpc1_1 gpc4349 (
      {stage4_10[25]},
      {stage5_10[19]}
   );
   gpc1_1 gpc4350 (
      {stage4_10[26]},
      {stage5_10[20]}
   );
   gpc1_1 gpc4351 (
      {stage4_10[27]},
      {stage5_10[21]}
   );
   gpc1_1 gpc4352 (
      {stage4_10[28]},
      {stage5_10[22]}
   );
   gpc1_1 gpc4353 (
      {stage4_11[19]},
      {stage5_11[7]}
   );
   gpc1_1 gpc4354 (
      {stage4_11[20]},
      {stage5_11[8]}
   );
   gpc1_1 gpc4355 (
      {stage4_12[8]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4356 (
      {stage4_12[9]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4357 (
      {stage4_12[10]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4358 (
      {stage4_12[11]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4359 (
      {stage4_12[12]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4360 (
      {stage4_12[13]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4361 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc4362 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc4363 (
      {stage4_13[23]},
      {stage5_13[11]}
   );
   gpc1_1 gpc4364 (
      {stage4_13[24]},
      {stage5_13[12]}
   );
   gpc1_1 gpc4365 (
      {stage4_13[25]},
      {stage5_13[13]}
   );
   gpc1_1 gpc4366 (
      {stage4_13[26]},
      {stage5_13[14]}
   );
   gpc1_1 gpc4367 (
      {stage4_13[27]},
      {stage5_13[15]}
   );
   gpc1_1 gpc4368 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4369 (
      {stage4_14[12]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4370 (
      {stage4_15[47]},
      {stage5_15[10]}
   );
   gpc1_1 gpc4371 (
      {stage4_16[18]},
      {stage5_16[11]}
   );
   gpc1_1 gpc4372 (
      {stage4_16[19]},
      {stage5_16[12]}
   );
   gpc1_1 gpc4373 (
      {stage4_16[20]},
      {stage5_16[13]}
   );
   gpc1_1 gpc4374 (
      {stage4_16[21]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4375 (
      {stage4_16[22]},
      {stage5_16[15]}
   );
   gpc1_1 gpc4376 (
      {stage4_16[23]},
      {stage5_16[16]}
   );
   gpc1_1 gpc4377 (
      {stage4_16[24]},
      {stage5_16[17]}
   );
   gpc1_1 gpc4378 (
      {stage4_16[25]},
      {stage5_16[18]}
   );
   gpc1_1 gpc4379 (
      {stage4_16[26]},
      {stage5_16[19]}
   );
   gpc1_1 gpc4380 (
      {stage4_16[27]},
      {stage5_16[20]}
   );
   gpc1_1 gpc4381 (
      {stage4_16[28]},
      {stage5_16[21]}
   );
   gpc1_1 gpc4382 (
      {stage4_17[32]},
      {stage5_17[12]}
   );
   gpc1_1 gpc4383 (
      {stage4_17[33]},
      {stage5_17[13]}
   );
   gpc1_1 gpc4384 (
      {stage4_17[34]},
      {stage5_17[14]}
   );
   gpc1_1 gpc4385 (
      {stage4_18[17]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4386 (
      {stage4_18[18]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4387 (
      {stage4_20[24]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4388 (
      {stage4_20[25]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4389 (
      {stage4_21[19]},
      {stage5_21[8]}
   );
   gpc1_1 gpc4390 (
      {stage4_21[20]},
      {stage5_21[9]}
   );
   gpc1_1 gpc4391 (
      {stage4_21[21]},
      {stage5_21[10]}
   );
   gpc1_1 gpc4392 (
      {stage4_22[22]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4393 (
      {stage4_23[19]},
      {stage5_23[11]}
   );
   gpc1_1 gpc4394 (
      {stage4_23[20]},
      {stage5_23[12]}
   );
   gpc1_1 gpc4395 (
      {stage4_23[21]},
      {stage5_23[13]}
   );
   gpc1_1 gpc4396 (
      {stage4_26[21]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4397 (
      {stage4_26[22]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4398 (
      {stage4_26[23]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4399 (
      {stage4_27[24]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4400 (
      {stage4_27[25]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4401 (
      {stage4_27[26]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4402 (
      {stage4_27[27]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4403 (
      {stage4_29[16]},
      {stage5_29[8]}
   );
   gpc1_1 gpc4404 (
      {stage4_29[17]},
      {stage5_29[9]}
   );
   gpc1_1 gpc4405 (
      {stage4_29[18]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4406 (
      {stage4_29[19]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4407 (
      {stage4_29[20]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4408 (
      {stage4_31[16]},
      {stage5_31[6]}
   );
   gpc1_1 gpc4409 (
      {stage4_31[17]},
      {stage5_31[7]}
   );
   gpc1_1 gpc4410 (
      {stage4_31[18]},
      {stage5_31[8]}
   );
   gpc1_1 gpc4411 (
      {stage4_31[19]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4412 (
      {stage4_31[20]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4413 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4414 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4415 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4416 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4417 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4418 (
      {stage4_34[15]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4419 (
      {stage4_34[16]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4420 (
      {stage4_35[3]},
      {stage5_35[4]}
   );
   gpc1_1 gpc4421 (
      {stage4_35[4]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4422 (
      {stage4_35[5]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4423 (
      {stage4_35[6]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4424 (
      {stage4_35[7]},
      {stage5_35[8]}
   );
   gpc1_1 gpc4425 (
      {stage4_35[8]},
      {stage5_35[9]}
   );
   gpc1_1 gpc4426 (
      {stage4_35[9]},
      {stage5_35[10]}
   );
   gpc1_1 gpc4427 (
      {stage4_35[10]},
      {stage5_35[11]}
   );
   gpc1_1 gpc4428 (
      {stage4_35[11]},
      {stage5_35[12]}
   );
   gpc1_1 gpc4429 (
      {stage4_35[12]},
      {stage5_35[13]}
   );
   gpc1_1 gpc4430 (
      {stage4_35[13]},
      {stage5_35[14]}
   );
   gpc1_1 gpc4431 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4432 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4433 (
      {stage4_38[0]},
      {stage5_38[1]}
   );
   gpc1163_5 gpc4434 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], 1'b0},
      {stage5_3[0]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc135_4 gpc4435 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[1], stage5_4[2], stage5_4[3]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc1343_5 gpc4436 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[2]}
   );
   gpc1343_5 gpc4437 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[2],stage6_5[3]}
   );
   gpc615_5 gpc4438 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc4439 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[3],stage6_8[3]}
   );
   gpc606_5 gpc4440 (
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[4],stage6_8[4]}
   );
   gpc117_4 gpc4441 (
      {stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12], stage5_10[13]},
      {stage5_11[1]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[2],stage6_11[3],stage6_10[3]}
   );
   gpc117_4 gpc4442 (
      {stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17], stage5_10[18], stage5_10[19], stage5_10[20]},
      {stage5_11[2]},
      {stage5_12[1]},
      {stage6_13[1],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc117_4 gpc4443 (
      {stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7], stage5_11[8], 1'b0},
      {stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[2],stage6_12[4],stage6_11[5]}
   );
   gpc207_4 gpc4444 (
      {stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_14[0], stage5_14[1]},
      {stage6_15[0],stage6_14[1],stage6_13[3],stage6_12[5]}
   );
   gpc1406_5 gpc4445 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5], stage5_13[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[4]}
   );
   gpc1406_5 gpc4446 (
      {stage5_13[7], stage5_13[8], stage5_13[9], stage5_13[10], stage5_13[11], stage5_13[12]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[1]},
      {stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[5]}
   );
   gpc615_5 gpc4447 (
      {stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[8]},
      {stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[0],stage6_17[2],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc117_4 gpc4448 (
      {stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14]},
      {stage5_17[0]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[1],stage6_17[3],stage6_16[3]}
   );
   gpc7_3 gpc4449 (
      {stage5_16[15], stage5_16[16], stage5_16[17], stage5_16[18], stage5_16[19], stage5_16[20], stage5_16[21]},
      {stage6_18[2],stage6_17[4],stage6_16[4]}
   );
   gpc1163_5 gpc4450 (
      {stage5_17[1], stage5_17[2], stage5_17[3]},
      {stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3],stage6_17[5]}
   );
   gpc1163_5 gpc4451 (
      {stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[2],stage6_18[4],stage6_17[6]}
   );
   gpc606_5 gpc4452 (
      {stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11], stage5_17[12]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[3],stage6_18[5],stage6_17[7]}
   );
   gpc615_5 gpc4453 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[2]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[4]}
   );
   gpc606_5 gpc4454 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc1406_5 gpc4455 (
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0]},
      {stage6_25[0],stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[5]}
   );
   gpc615_5 gpc4456 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[4]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[0],stage6_25[1],stage6_24[2],stage6_23[3],stage6_22[3]}
   );
   gpc615_5 gpc4457 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[7]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[1],stage6_25[2],stage6_24[3],stage6_23[4]}
   );
   gpc135_4 gpc4458 (
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4]},
      {stage5_27[0], stage5_27[1], stage5_27[2]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[2]}
   );
   gpc615_5 gpc4459 (
      {stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[2]}
   );
   gpc606_5 gpc4460 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1],stage6_29[2]}
   );
   gpc1406_5 gpc4461 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3]},
      {stage5_33[0]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[2]}
   );
   gpc615_5 gpc4462 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {stage5_31[6]},
      {stage5_32[4], stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[3]}
   );
   gpc606_5 gpc4463 (
      {stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3]}
   );
   gpc606_5 gpc4464 (
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1]}
   );
   gpc1_1 gpc4465 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4466 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4467 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc4468 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc4469 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc4470 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc4471 (
      {stage5_1[6]},
      {stage6_1[4]}
   );
   gpc1_1 gpc4472 (
      {stage5_1[7]},
      {stage6_1[5]}
   );
   gpc1_1 gpc4473 (
      {stage5_1[8]},
      {stage6_1[6]}
   );
   gpc1_1 gpc4474 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc4475 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc4476 (
      {stage5_5[7]},
      {stage6_5[4]}
   );
   gpc1_1 gpc4477 (
      {stage5_5[8]},
      {stage6_5[5]}
   );
   gpc1_1 gpc4478 (
      {stage5_6[8]},
      {stage6_6[3]}
   );
   gpc1_1 gpc4479 (
      {stage5_6[9]},
      {stage6_6[4]}
   );
   gpc1_1 gpc4480 (
      {stage5_8[12]},
      {stage6_8[5]}
   );
   gpc1_1 gpc4481 (
      {stage5_10[21]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4482 (
      {stage5_10[22]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4483 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc4484 (
      {stage5_13[13]},
      {stage6_13[6]}
   );
   gpc1_1 gpc4485 (
      {stage5_13[14]},
      {stage6_13[7]}
   );
   gpc1_1 gpc4486 (
      {stage5_13[15]},
      {stage6_13[8]}
   );
   gpc1_1 gpc4487 (
      {stage5_14[7]},
      {stage6_14[5]}
   );
   gpc1_1 gpc4488 (
      {stage5_15[9]},
      {stage6_15[4]}
   );
   gpc1_1 gpc4489 (
      {stage5_15[10]},
      {stage6_15[5]}
   );
   gpc1_1 gpc4490 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc4491 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc4492 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc4493 (
      {stage5_22[11]},
      {stage6_22[4]}
   );
   gpc1_1 gpc4494 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc4495 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc4496 (
      {stage5_23[12]},
      {stage6_23[7]}
   );
   gpc1_1 gpc4497 (
      {stage5_23[13]},
      {stage6_23[8]}
   );
   gpc1_1 gpc4498 (
      {stage5_25[6]},
      {stage6_25[3]}
   );
   gpc1_1 gpc4499 (
      {stage5_25[7]},
      {stage6_25[4]}
   );
   gpc1_1 gpc4500 (
      {stage5_26[5]},
      {stage6_26[3]}
   );
   gpc1_1 gpc4501 (
      {stage5_26[6]},
      {stage6_26[4]}
   );
   gpc1_1 gpc4502 (
      {stage5_26[7]},
      {stage6_26[5]}
   );
   gpc1_1 gpc4503 (
      {stage5_26[8]},
      {stage6_26[6]}
   );
   gpc1_1 gpc4504 (
      {stage5_26[9]},
      {stage6_26[7]}
   );
   gpc1_1 gpc4505 (
      {stage5_26[10]},
      {stage6_26[8]}
   );
   gpc1_1 gpc4506 (
      {stage5_26[11]},
      {stage6_26[9]}
   );
   gpc1_1 gpc4507 (
      {stage5_26[12]},
      {stage6_26[10]}
   );
   gpc1_1 gpc4508 (
      {stage5_26[13]},
      {stage6_26[11]}
   );
   gpc1_1 gpc4509 (
      {stage5_27[8]},
      {stage6_27[3]}
   );
   gpc1_1 gpc4510 (
      {stage5_27[9]},
      {stage6_27[4]}
   );
   gpc1_1 gpc4511 (
      {stage5_27[10]},
      {stage6_27[5]}
   );
   gpc1_1 gpc4512 (
      {stage5_27[11]},
      {stage6_27[6]}
   );
   gpc1_1 gpc4513 (
      {stage5_27[12]},
      {stage6_27[7]}
   );
   gpc1_1 gpc4514 (
      {stage5_27[13]},
      {stage6_27[8]}
   );
   gpc1_1 gpc4515 (
      {stage5_28[2]},
      {stage6_28[2]}
   );
   gpc1_1 gpc4516 (
      {stage5_28[3]},
      {stage6_28[3]}
   );
   gpc1_1 gpc4517 (
      {stage5_28[4]},
      {stage6_28[4]}
   );
   gpc1_1 gpc4518 (
      {stage5_28[5]},
      {stage6_28[5]}
   );
   gpc1_1 gpc4519 (
      {stage5_28[6]},
      {stage6_28[6]}
   );
   gpc1_1 gpc4520 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc4521 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc4522 (
      {stage5_31[7]},
      {stage6_31[4]}
   );
   gpc1_1 gpc4523 (
      {stage5_31[8]},
      {stage6_31[5]}
   );
   gpc1_1 gpc4524 (
      {stage5_31[9]},
      {stage6_31[6]}
   );
   gpc1_1 gpc4525 (
      {stage5_31[10]},
      {stage6_31[7]}
   );
   gpc1_1 gpc4526 (
      {stage5_32[10]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4527 (
      {stage5_33[7]},
      {stage6_33[4]}
   );
   gpc1_1 gpc4528 (
      {stage5_33[8]},
      {stage6_33[5]}
   );
   gpc1_1 gpc4529 (
      {stage5_34[0]},
      {stage6_34[3]}
   );
   gpc1_1 gpc4530 (
      {stage5_34[1]},
      {stage6_34[4]}
   );
   gpc1_1 gpc4531 (
      {stage5_34[2]},
      {stage6_34[5]}
   );
   gpc1_1 gpc4532 (
      {stage5_34[3]},
      {stage6_34[6]}
   );
   gpc1_1 gpc4533 (
      {stage5_34[4]},
      {stage6_34[7]}
   );
   gpc1_1 gpc4534 (
      {stage5_34[5]},
      {stage6_34[8]}
   );
   gpc1_1 gpc4535 (
      {stage5_34[6]},
      {stage6_34[9]}
   );
   gpc1_1 gpc4536 (
      {stage5_34[7]},
      {stage6_34[10]}
   );
   gpc1_1 gpc4537 (
      {stage5_35[12]},
      {stage6_35[2]}
   );
   gpc1_1 gpc4538 (
      {stage5_35[13]},
      {stage6_35[3]}
   );
   gpc1_1 gpc4539 (
      {stage5_35[14]},
      {stage6_35[4]}
   );
   gpc1_1 gpc4540 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4541 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4542 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4543 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4544 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
   gpc1_1 gpc4545 (
      {stage5_38[1]},
      {stage6_38[2]}
   );
   gpc223_4 gpc4546 (
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0], stage6_6[1]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0]}
   );
   gpc135_4 gpc4547 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[0]}
   );
   gpc615_5 gpc4548 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[0]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1]}
   );
   gpc2135_5 gpc4549 (
      {stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage6_14[0]},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[2]}
   );
   gpc615_5 gpc4550 (
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4]},
      {stage6_17[0]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1]}
   );
   gpc7_3 gpc4551 (
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage7_19[1],stage7_18[1],stage7_17[1]}
   );
   gpc615_5 gpc4552 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4]},
      {stage6_20[0]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[2]}
   );
   gpc615_5 gpc4553 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4]},
      {stage6_24[0]},
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], 1'b0},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[1]}
   );
   gpc7_3 gpc4554 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4], stage6_26[5], stage6_26[6]},
      {stage7_28[0],stage7_27[1],stage7_26[1]}
   );
   gpc7_3 gpc4555 (
      {stage6_26[7], stage6_26[8], stage6_26[9], stage6_26[10], stage6_26[11], 1'b0, 1'b0},
      {stage7_28[1],stage7_27[2],stage7_26[2]}
   );
   gpc7_3 gpc4556 (
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5], stage6_27[6]},
      {stage7_29[0],stage7_28[2],stage7_27[3]}
   );
   gpc1325_5 gpc4557 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4]},
      {stage6_29[0], stage6_29[1]},
      {stage6_30[0], stage6_30[1], stage6_30[2]},
      {stage6_31[0]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[3]}
   );
   gpc7_3 gpc4558 (
      {stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4], stage6_31[5], stage6_31[6], stage6_31[7]},
      {stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc606_5 gpc4559 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], 1'b0},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[0],stage7_33[1]}
   );
   gpc606_5 gpc4560 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[1]}
   );
   gpc1_1 gpc4561 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4562 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4563 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc4564 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4565 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc4566 (
      {stage6_1[2]},
      {stage7_1[2]}
   );
   gpc1_1 gpc4567 (
      {stage6_1[3]},
      {stage7_1[3]}
   );
   gpc1_1 gpc4568 (
      {stage6_1[4]},
      {stage7_1[4]}
   );
   gpc1_1 gpc4569 (
      {stage6_1[5]},
      {stage7_1[5]}
   );
   gpc1_1 gpc4570 (
      {stage6_1[6]},
      {stage7_1[6]}
   );
   gpc1_1 gpc4571 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc4572 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc4573 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc4574 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc4575 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc4576 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc4577 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4578 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc4579 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc4580 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc4581 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc4582 (
      {stage6_6[3]},
      {stage7_6[2]}
   );
   gpc1_1 gpc4583 (
      {stage6_6[4]},
      {stage7_6[3]}
   );
   gpc1_1 gpc4584 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc4585 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc4586 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc4587 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc4588 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc4589 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc4590 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc4591 (
      {stage6_10[3]},
      {stage7_10[1]}
   );
   gpc1_1 gpc4592 (
      {stage6_10[4]},
      {stage7_10[2]}
   );
   gpc1_1 gpc4593 (
      {stage6_10[5]},
      {stage7_10[3]}
   );
   gpc1_1 gpc4594 (
      {stage6_10[6]},
      {stage7_10[4]}
   );
   gpc1_1 gpc4595 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc4596 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc4597 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc4598 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc4599 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc4600 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc4601 (
      {stage6_15[2]},
      {stage7_15[2]}
   );
   gpc1_1 gpc4602 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc4603 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc4604 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc4605 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc4606 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc4607 (
      {stage6_20[1]},
      {stage7_20[2]}
   );
   gpc1_1 gpc4608 (
      {stage6_20[2]},
      {stage7_20[3]}
   );
   gpc1_1 gpc4609 (
      {stage6_20[3]},
      {stage7_20[4]}
   );
   gpc1_1 gpc4610 (
      {stage6_20[4]},
      {stage7_20[5]}
   );
   gpc1_1 gpc4611 (
      {stage6_20[5]},
      {stage7_20[6]}
   );
   gpc1_1 gpc4612 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc4613 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc4614 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc4615 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc4616 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc4617 (
      {stage6_23[5]},
      {stage7_23[2]}
   );
   gpc1_1 gpc4618 (
      {stage6_23[6]},
      {stage7_23[3]}
   );
   gpc1_1 gpc4619 (
      {stage6_23[7]},
      {stage7_23[4]}
   );
   gpc1_1 gpc4620 (
      {stage6_23[8]},
      {stage7_23[5]}
   );
   gpc1_1 gpc4621 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc4622 (
      {stage6_24[2]},
      {stage7_24[2]}
   );
   gpc1_1 gpc4623 (
      {stage6_24[3]},
      {stage7_24[3]}
   );
   gpc1_1 gpc4624 (
      {stage6_27[7]},
      {stage7_27[4]}
   );
   gpc1_1 gpc4625 (
      {stage6_27[8]},
      {stage7_27[5]}
   );
   gpc1_1 gpc4626 (
      {stage6_28[5]},
      {stage7_28[4]}
   );
   gpc1_1 gpc4627 (
      {stage6_28[6]},
      {stage7_28[5]}
   );
   gpc1_1 gpc4628 (
      {stage6_29[2]},
      {stage7_29[2]}
   );
   gpc1_1 gpc4629 (
      {stage6_29[3]},
      {stage7_29[3]}
   );
   gpc1_1 gpc4630 (
      {stage6_30[3]},
      {stage7_30[1]}
   );
   gpc1_1 gpc4631 (
      {stage6_30[4]},
      {stage7_30[2]}
   );
   gpc1_1 gpc4632 (
      {stage6_32[0]},
      {stage7_32[2]}
   );
   gpc1_1 gpc4633 (
      {stage6_32[1]},
      {stage7_32[3]}
   );
   gpc1_1 gpc4634 (
      {stage6_32[2]},
      {stage7_32[4]}
   );
   gpc1_1 gpc4635 (
      {stage6_32[3]},
      {stage7_32[5]}
   );
   gpc1_1 gpc4636 (
      {stage6_34[6]},
      {stage7_34[2]}
   );
   gpc1_1 gpc4637 (
      {stage6_34[7]},
      {stage7_34[3]}
   );
   gpc1_1 gpc4638 (
      {stage6_34[8]},
      {stage7_34[4]}
   );
   gpc1_1 gpc4639 (
      {stage6_34[9]},
      {stage7_34[5]}
   );
   gpc1_1 gpc4640 (
      {stage6_34[10]},
      {stage7_34[6]}
   );
   gpc1_1 gpc4641 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc4642 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc4643 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc4644 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc4645 (
      {stage6_38[2]},
      {stage7_38[3]}
   );
   gpc1_1 gpc4646 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1163_5 gpc4647 (
      {stage7_0[0], stage7_0[1], stage7_0[2]},
      {stage7_1[0], stage7_1[1], stage7_1[2], stage7_1[3], stage7_1[4], stage7_1[5]},
      {stage7_2[0]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1423_5 gpc4648 (
      {stage7_3[1], stage7_3[2], stage7_3[3]},
      {stage7_4[0], stage7_4[1]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc623_5 gpc4649 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc4650 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc4651 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc4652 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc3_2 gpc4653 (
      {stage7_19[0], stage7_19[1], stage7_19[2]},
      {stage8_20[0],stage8_19[1]}
   );
   gpc7_3 gpc4654 (
      {stage7_20[0], stage7_20[1], stage7_20[2], stage7_20[3], stage7_20[4], stage7_20[5], stage7_20[6]},
      {stage8_22[0],stage8_21[0],stage8_20[1]}
   );
   gpc117_4 gpc4655 (
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], 1'b0},
      {stage7_23[0]},
      {stage7_24[0]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[1]}
   );
   gpc2135_5 gpc4656 (
      {stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5]},
      {stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage7_26[0], stage7_26[1]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc2116_5 gpc4657 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4], stage7_27[5]},
      {stage7_28[0]},
      {stage7_29[0]},
      {stage7_30[0], stage7_30[1]},
      {stage8_31[0],stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[1]}
   );
   gpc2135_5 gpc4658 (
      {stage7_28[1], stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5]},
      {stage7_29[1], stage7_29[2], stage7_29[3]},
      {stage7_30[2]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[1],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc2116_5 gpc4659 (
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage7_33[0]},
      {stage7_34[0]},
      {stage7_35[0], stage7_35[1]},
      {stage8_36[0],stage8_35[0],stage8_34[0],stage8_33[0],stage8_32[1]}
   );
   gpc207_4 gpc4660 (
      {stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[1],stage8_35[1],stage8_34[1]}
   );
   gpc135_4 gpc4661 (
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0},
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0]},
      {stage8_40[0],stage8_39[0],stage8_38[0],stage8_37[1]}
   );
   gpc1_1 gpc4662 (
      {stage7_1[6]},
      {stage8_1[1]}
   );
   gpc1_1 gpc4663 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc4664 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc4665 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc4666 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc4667 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc4668 (
      {stage7_21[0]},
      {stage8_21[1]}
   );
   gpc1_1 gpc4669 (
      {stage7_26[2]},
      {stage8_26[1]}
   );
   gpc1_1 gpc4670 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
   gpc1_1 gpc4671 (
      {stage7_38[3]},
      {stage8_38[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor_CLA486_32 compressor_CLA486_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h400f4356a9050a1f78d54164f4ec4887c41931923e37efc81d7643d358781d27b9ef37cfbfdafe20dafad98af0eded2eaee4a5f56ec026b2f57a669f8f08f6495ea628cb586f39a11090d6dd2d1367ac33bc6c720ad4073d0b46a47c1929e5ac56a9151616838e9585e1bea310bb781708bfaffb661074dbd34e77f84dcb9baa1f134c573af9b8decd1dfa4244ec598c8c89e0dd11613b18ae6b5ffb4318c011904316d01d0c56fba7a60aa16cd1f242c121eded13432e19ea247301f91f351cb2fc9635d3ae83f80cb04e7632d08d9e562109d1321950bd69da5c3209e4314ff5509509d511549a68b7790dca954b3a2d97530726138a3ac335469c7c1714d90b357039eacd882d0ba382c9c61c53f9f4000eae5910d2984fe89cec435e6b30765692a7c91f69bd421d5e7306bd976721ed5d499db95a4b7cab4efdd9d945e1c999796efa2213ab9fa8a07145c3ba56d14bb8b6d1597976062ee4005acf6977c9a74ed6b03aeafd87d44450b9e388061defb7bd835d6db2f521be4fa0526b01993a13247ca4a80cce4a2714a136d5e120b300c9cc527d38c676e22eb566697a35b730f6628a7719d7e97dd969138cdb348b822d689a85421b73d9efaf00bc8812e29c6fd3ec02f02c68f7e80b83c40cccbea016b95f4bf789a7f7a7a9bc7a094be48b9f8c39a9ef40aeeac1f6635ee9aeb14a92a2a29c7fdf8d8d8e31c8daa6accd60f04e2eba287f5d40195d8bc18d36e9631329824ea3d8024567fff853309908f5a07e85a27c53428d3429929155823f7c28a1759b671497bc03621ac0beb210e4c24911a14367805052a927baf499e95918ebcfceadb9f33addb1e7a913d5c958a28e64ccc44a91d10f614b88958cdc8c7556d1eab9509ddff1bd4e8534a3cb89833407f1c8e5134c07e0ea966843a972efab247491dc6a1bd179cbd09977565b2c522e92be01245484843f2f1c4220ec8b736bd2134f5b2e201310da355ad9c73237478b28c5b834534fc589e87fc346b50384b193001ac3f669f55dd58146743cf280e2970cb6c66adfffc467082a5966804088e3965eafa0cedbb6931fcc54ec8de608e7e7d7ae6abe396642b3e242e465379e309e01c213c9df869f1655c92785e823ab5a0e1264ef943f12d14dc19a819f650c3f409c64e1b5ed9879d0c328a1759ee5307034367c4d1f416f8c3f0d6cb7a922d0c4b537537c172727c60d03dbfed085b63c2be5eb68b437969c549ffe01a282bc5c373bb941811c121f97f79bade7bad81c150abf34f8b2f3ddd4ba5db70360314b342ace0a46605ebae44000b6a19d8c5406f358c8fc2dca6821c62d62554c5704ef3f5228e0119c96c5e68955f9300d33405219cc3f19c0c89f23da1c0f68b983e6c75ee8a4d9f510e896643ef6838ca999ffd8a86665a5958f441f4495e1f19744aa955a0f0357a8f64d40fcca588065940738d81f615c7bf5ce357172bcc1a6cafc40309d351e6fc27d6fa37a49273e0f97e04615e5e6115eba69f2a5ecce0b219feb50105749ebeaf394542f0842d0d1a42df50a4b067d5868e57d486ab43780ebb3d064d9666bc8332d7d1ebcfd6843b9bc2a41618d207b073ab4b8f91775126754d15377e98f504fc5a73c8fab012a4b618232989fe570097b84119bc3d62bd177414454b1964ee3663808fa8e52e1c1667ffa533b553c646da41deb7f10cf1547fdd34c505f16a587cd2d373a6703bfde0675b1a83ffc24bc5c3b454f4f1ca5535066439e747b07c6d3d2df0ab1fed7fc819fae63023bf2834cf3e8f0c2e0325e8fdc6e7fb4d428e80b256eb7ff8e5bd635322c71399f11ca0ec31e009f5b960aa241d664f5cfe0de9e71f735a4bd3b2ae0c52e5f990fe293366c028f32e0fdd01d4bb03fa469feaa81c4ae7a78a9e901648881fa1e31e5d260d5f301bbd208cddb3f659128eacacb8425b4387f4fe9f2674edd335671c609a4f1a8c877b3e41e071c85dd3d89984bd5ed5057b32ae055007158e677f6e398371961567738ac083a817be80a98b563dd56dbd69c7ccbf07a92a6b151ded4a1a8c70f3d3455a67f2a5df21c4ca06fe5baa0e2d7bc0ab6c561ef93502975c4d4f247892d36ba134ea700dd4fd309e8c6807be8bcf8953cc6ab4eb7782cc539ba16935eddb73954d6a008fb21b4231b1de10e5c7ff99c3cc9229ed369718b0443c1350f44d5b161d8d8a6996319fde971bd2c6ad3c6354771ad178f1a204b7a5f7e70683eb8202749bd247d84d55d0f257fea8f9ab132371274f073abc953d13d1479978dff831086abe7ffb33efabe171d568c9b59be65584ce6163e27a06de083b7033a173718a6750feb5e8ec5c34b915729e40f066bcc0211793bf1c8cc4e4f81dc5e82d4fe0b999a553f78e0b1d9ff34a25881981328c64643a710f343170d778bf6257c43092167a44c555de73327f8d2804df26df3d729efa5f6461ede1b2cadf10a1df99a6bf2c2c90f4a52f0bfcf8546782e1e06d25c0ecd254bbac3ce57272ebecc1c333bdf6f8da2006ab65f8a43c6dd0b79ae54e17e5e769367ea5e199e3edba6ce7007884d6e79792c32f18c2274d39ebeae15f536475ad7f61b72ac8d0751f2d88400b0fa9412afdef3c4043949f8aea032dbbc3054ad7e3ac23fdc5b34fe68b8e47af47683d1e3012b27a053f7f2f4ea74a5fc7a5229924bb356dd439b3c5b2d8c6bf9af9aa15fbda56a4abd40bc1960cd2ca0a6b5119f7e9a5c3983;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7bd19c5d0a12ff039c85edb619df944e05aa81cc2aa73868b5215522776041c9c47efa8c0307b7faf4e18a66398d4525b571b6bcd567f103e60e9354dff4ff196b8baa16a38a54aba99a7bbb5423e9735fb180aefe23de8da9f507ba937672bb020016639b23f7619790391b6b72fd43568829d92f4724acc10bd50ca58de5daa6ee4751b4449f2e097bb274a1fd562a250cbdb7ea0a7faf61c14beffd4b5320d866f715d46627c021fdb99ec4b70beb3f7fd54232e604fd378ff47cbb427e5ce625a6369d01f40b4ef1557d1bd8450491e2b29d4625489da16a63e6f380236269804dfc2269977144ec39af2062760a29c051976d46060c9981bc51580f5c85b08d81d24518237e918120974e5fc005ffeb161f0aca80c1173c15d1c360d2f5607fe82284437eb450a1b450fd3201f90de73fd4bd1d472418dfbca8d93fa8b26c10b9b239137bcad0b2de6041842c14fe876b871ec511a18186dfa6d9d38f38e13fe3745cda8037a2269d1c1a142e2fb86d9c8d92129f30f015da4863fe58d3a5dfc14555e730452f06660dc73959a6a17122f1b3f944b7359a7068b59462585971f5d9721003c59dc35bef22a8a4213bf740000675ad223671b9ae3da95ec7422bf91d2711872a71883169bbd623b175047864c70df4bc8c25abbd2c8e6eecc1dd6716ccc91baaa9dbacc9229e5ae388fffff57890cfb46a0c095e7adb8e0f98c28eb8d6894fd1d725ea3b9b7e7281dc5636da6b288c73d7d277fb3549f0e1e47912c1135ccfb3e33d4c33ad9f330dd1cbd6cca6b8a04caf09235ca534218efe81515bafbfbc18619b8311531ea5ed243478f2cb4332d4d2366fed3652668f847f42476c809f2e523530f0f30379a54e326ea0e345206cb2f9fd2ae5bc0deeac30d078f984e0639c0ace4ab3d9598e4c5b2747e89583fbb1b56f74b76f6bb1d1c1277702d6f54ba6129f1132408cc647d398c3a29f53c8f5416c9ea6c5c9fd39787de5f767bc8d2080835ff2fbdeda7ba9b3b0e451bbfa0f06f9850d4613753f5e6218f5d39ed8eefe9bd38a86b1222d755d7b2de44a55f273ef338730149e35d3ef0d74af846d78b62e06461bd3a1d0886b834eb0b00f0cbaa60c4de70e028cdc3fec73256b241ba5aaba687d26987445de411d8ea361e249601bbb1dfc1af67be2880b652c319c655b72da7c285242bd32b915ee10d973f66057c8b3297109a2f20ea6afa1149d9f9bc4495844c31137e6e504e9b0a962ad79067d0d7a0ae0702e990e40618134832f88a38a6e737ec0bcd0a62003a4aea8984bbcd1dd48feee4d2e6d162375a844c3553a9265dd7769c7eb2247f7967f9391bc1ad77a6458e2e88440c0edbe037887460ed6a4e0fd0894ac6b82e228d2d0c425afbdbb8c81f78af729fcb7d363b5f7316559a34d3c2de5cf6d4e18844ee1b78e97ca5c82d95cf74fedd4d89e81b21360bf66ab466079113203d88bfae334e5511f76ede8092db042dd0452ec0542cb53850b698cb9de36db9aa32ddec8fc34fc5182c6569040286d239939c87d90843c2e0f874a372e9c5b4bd4921e0eabdd9415f332664743007dc225c6a7e4548d4504231adbf5fa0793ad5d5885155daea37aae774249f76497fcdd130f7e70b76e5176a63cb557df0ce56f261fa4f0e515ddca617acc5abe592a813e649caf72bc74a0d6bb5ae5be4110dbb0db60cf676650cfd6203f284a277f4b71075eb5f4acf207a0ce6c87d45bc7ecc002bc3b4d4d4ddd33cdbc3062544ca3e9f9f55802bcc5947fe616bfd30fdeae27b1457cfac33c3fadb6c4c7f48a3836687c588cc13793dc19fb12bfc8020e55052ad9addb8545df923d60d75a761d5f3aa6d3d4054596e2a79c240e57f9a88fb2b31d0ceffd5c3abf72a68f1562d3f4b815a0ad58f76a783829ba8db68b5a4426f9f054fdff56615ea4e5146c6b4982e23a892bb2a6c2585fe4d84b9f304f139fbdc4a71e06364e15312995c94cb8df90a9bafd94daaa341976cfe0b11b0c3ecbd1f57dd7b2560bea52c8d84a0e8dd5187dc98bda505816c1de70fe225cdafeb382b4bf2d17ae823825790b427a07c1a61d4040c0cc44b30a0aa8f6bab28c5d9ed119c1b8afbcef4323133c4ae1bbf092c1d47acde457bc1fe8f0a04755d6d5914d537478c43ee4a56d495e849e67918ce213a828e003853e1fe295b31d1186b9433667f80764426d10f5a8723c46292ebbfd5241ee3a12b05a719c8bb28de25afe0cdfae79bfb3b047996296d7ec21b0fd298703efddbb9b51f7ee35da33b6456fab75ec3726e4f9fa459b96d5349599e0730d6d089600a9a4d5ca95215c900f9ad2b46cbe46032680e27e443da81dcd797fb45680e12bf15482748ef3670065425ab3038944d816dc304f4f5ec1104df7b30916ebf2dce3ee40894401d6ecbf93dd4eaef15b1f5fefd3d69882b86d862176b9b8f379e5862f3d2d8a00bfbf8effda4955340d4fae45762c218941d6252a9fac257d8feccc7f3b5630f8625aaffab8c44ea80ffb5b6917e6a7950f974dd9ad3aa7b4cab878b0fabdf2a89841ac476fb6f3693c60753883df042907df52ea90d8fb563872a77e2b501f22a48cab8bc270a4404283debfac1c35534ded900c96098de9ab845c5305051ca24066ca00170c78580ff75c437dd838daf99d65aae5b3c3668bf51505900f543df619633ba19915b9cb2e91ea535c0d764131a4198678cc30ab2ea5cde68cb6430da45d3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb741e8286a1e19eea542a54ce1d80fad3f36f03dc9d3c26cf4281c1a2eafb6d05fa9cfb32afc6566843b13ca6fa3f2e0f510bdc1aa84a77c453a126690fc55492253516a3e9b07219fda99d2d7c7ac182aa4ac074283f991b6e694bd98ad932e527ba15bf1378ced68e3037ddd2a214d752ecf70064ad5c2620adffb5f3f488cb4ec5f914bb48991c21b1b01d0dbf96464daa5411ec9cfad9aee80ee3ddda6354c1d149d2b0d78aac201fb85b8407fc00aba566d1c01eb0ebb8b88f19245b238c11405dd80ea4cf146f4d054620d489634de5d16048fe926aa2710edcef00da4f6ced2ef38721e22a9d5008169b42d93d58f1b50fd3ecac334939f18f1274b67845a39a777dec63301b41daf43ccce42acfe0c56e3a0602f0c4c32a716a4d8bf051c1e956a00c69dd3f2e11194ad52bf56e428ff9bbb55eab8568aa2db75c62eec08c9b6668d79d5cf88348e7e36434ab35ecab324804bfaf781e2359f300120f492082b4f9996f170c7ca656ec5416f449786decf5606822978da7d5d158bb3ad8984964dc20cab09c0a9f75463277d7dfc1a339c228a84d8b10e41059757a62f38ac6480bc1964fbe9da97fe101652b9662b8d2d710143d994dea86c5aacfd89477bdcfdb8cad8ae62abaf9ac3fe1e2b211e46d0dea5e3c57d17beae1d7ee6a23db34c14461da6691fcf2ba88d88063f36e3521d6d34e42c7cb5c48bcd1e73dd692b789541a2dfb6699be9c7d5754be42595ed1e501d20a4babd1590fdb0609165d3752fd667661966a85d890577b68132e73e979cc8f2ec1cd552eff80bfc14dd754bde124e40cf3da91f22a274f9017e713afe303f1a7b953d047e8cbcb6e85d7fc7a5f2a76e855ffd2a4034d2e76e79b0f6b30039d186f0eef34fefd7f0b183e2c81a961fa6aa963dad5b6d40c24314d0ce391088613004c4bfe94e14ae78f0eae283682c0bef89f0cb04947b537206c213c40ac849d6634fb697044cde9cab3260ee9bebe1891de0e7789cf6ca37561ec13ed562e165a6257aa007823baafc5b086b34dab2b9fadedbe76cb2cebd7801574cd1c901572ebf18a53a900921f108025f2bac21edc993a368190a2623f5656107eb0c9e827d5ae48641d0d385280f19786971f23e925f564fda45f3befa8e7892a506b29a65428ee76c1c98ffb7968d45f3e0fafb3ba9a085a9da87368f1500865f09082f95d9879bcf36d99e1582df454359a2607fff827f24be52f6f460f3cf51d386a19daebe83e06f691e2f4abeac813acbdb7b7218211a0d914b8b2d39ae66f5b2c64247b70c16202a63d5d49cb3dbac299ec85b21de08912f04eef8d9dd09b5fd2cccf22e0177e5e7e133e1daaa2c895a5f8ce2917a6f77800db2486cc842f6036a588dc4cfb1379d700e742cd99702ab7753b2d14dcb5344a518232e6ec3f3185b45332345976d36c7574ceab24bfb6e36cf3c0c6a55807c7c1283078d9756e8290147f0085bc273fc4533791f2778fb9419b82bd742921e118436eb3a3efdf5bf1b436da99729c2e1782ca7942c3a733ff04d0ee94868ed9192f0795bb54b7b50864d3599a201930ef357669c50682eed244b786d833940d4516d40e3c9f79a60cf3257e066a4f3242ee5965e269fa4169555bf0d5a014aaa7513ef4e18ecad3f994ed4037f4757e68f33e5a952b7e4013f21771dd6b2acd21792a5a215aed470b0759e3affa772b6bc3cfaa6d84e9dd7bb3df3f828ad0d5c8a6b8225120df0b2308b08cfd2d98db6272613aaee0cf8e9210b09781cf44382b5b0f24fa1a9a1bbbc5339734857d028d2f63c8824f39a7ad7b334f7d47b420b50d85ebdd9a15339ac75f279f10f21197de0d9d3490ada9c4adbf9235128696008eb479f49e473cece3c8f33b9254d5e3251f7d67774110a6390cbbaf957bf38ca191b38bf0cf64c86e70bf334ec21310b1cf484ff0d0c846e14c214386f08aa63ce5346479c7b4b6c2238bf010ec96ea22c91b8e99b2fb2469d022f503bfbd5fac9678bbd04148bbbf3b745e64d82045916d0f5336f9faec9db763fcd16e8555ba8d2f11f5ea6bb17785f13ae3a18c6a951434129c9c9625a22d02c4a6fb16771928fd2ac351a67c269c139207b1b9bf2eb032dbb553c9cfe3dd7984ee0364492052a85a640a4bd378cd7b0764a193d3cc4fce8356e5fda050cc7d7c2197623786ff6033cf8ccfcfc9d6615eff8450c6b93405873c10104c5ea058e5dacffe97a94a5c76cbe7b326c890ac32c802dad7723e3e421178ebb9efb2586329323b7c3c1d6ab5c5a4b64b3030901160548574e740a4080e9b420947f0306d40b569c343d43e281e68f1789d1714f23079e75019ca31eb32208c7aaccc1985ab7893122751b6b1fc6ce0b5e8fac781c6066c532d46003b42349146c682fbc5a5a2ce41efdd216760d488a1cbd509a0996199110d322dc0f4b61e84bf7cffd64f52eb4c6b01a5aa0a5f9c7d3a120a740ad622d60d9bba21d04b2388def914268e95d686c7d6fd5ade3cd985ac2b0a5dbf8c08481909d0e3869610b6bc6a3325571bcd161f837ded75ea325c5338bdfb1fa8ff5accc9e1e91fd9fedfe50d2f159876aedade44b23e52904230dbf34acc34e1c41e3e8ed246b3aa8169e5211c3691292d374311b5be0763e13e2492087e52a07e33c12a0b2737ccb6843ab42e2b6deef483eadc28e524f5ddf7ed516654cbae7f07517ed78bba49387b1b2f63a43d4cdfc411b34ac17dc2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4e37ab59f29b114f58c0fb7eddf22c282c3f1b71d788c561d625fb67326fa1c847d13f3f837c3b5a14d3eff5bd89650cca70dbfbbaac4ecea1b56c6b004019720b096a31aed84ba5b1bf365825f5d68c4b68926559b90ab9840c205f7ea990d924cfd225a8e2e83266c1d2428b75bbd6f41d77abf8dd43372e66c6a15ff4b4756bb83c6ac9a8ae0754c361144d6db974d045fcb940029f03415ae21aca758dea97ea12335a883dc2da665817f43313e5619fde23a9e1f8b21dcea9ad0f5b7e398b60ee4d8afd3a19274b63d96f54befb82a2c4e775b436e14c3240461cb7851f7af83b0b5cecbaeb26f8b7725a2960eb636c0f2b96781381b8d1034be76b0d585193cb9a79ff0142651252a2e4a9d78dfb370e7161bae6ae5efc3b9356b26236d679489781234d8d0e821b5f33254b591c8669f0340d6cb74da2b58dd3a68e36af4c16746d78d88521d710e317c68bc690048e68d2d0c0eb31b5caba52f0932c3dd7f92a41a225bf8e925172eebe32c414bab2c52602909503f0367ead9a68d2f5fbd1f3909e4ea9ac84d29b1772c4334e8932f4285918ea5eb776b4e40e05f80bd102c461cd716a492be98d345c5a5b4d63f93300ec5743fb981a69575783335a129801c3a6671c499337bd929fef74479cb98782b9f366b61384702738d1ff02da2d6b4a84ff0bd6f8f6e341d7ea9613492c907ca8991d487ad853f9afd26614a6bb71e0a038ac91a0ed99839176052eaff44b45f7531804489c24a399f9f2cfa5c6e6e86f38a01a77b7cd6fc986728624a26bf594fd9ef44af660d85e531af3778efa1a16709e1a28f50ea8ded4ea649c6b125afe1d11db02edd0f6f85ba5a010f9df923eedad582c0116ebe7018737fbb55ee607b6949137fe3733052efd71dad32faada5f9a405872435bead1d5d76b5ebb1c8c4183820737956ee6a6c79601f1726ab9a3f58a13831fb594772dd228207b32ee7df64ddd7f80c64c1e8abdfa794a3be861a4ea80e35a912560b33a60c1e89fea2cce155faaa9f88c434ac9cc9b51bcb8e8503be5f733bbb38d807d9e1af0f0b9b9412eda2dd953feab17c64eeae9dbbc1aba4fba61d7661d1e8e194558bd0f22ac81048c01a4718c1ad62a5479caa9ae93829d050ef6eae7ff6e3fabbfdaff0a7a7278c424803fbad2850b79b8c0de6c17002c18bbcebc8781ed879b7fba1bed55130e0aa4a4fbd11bbf553ee12b7e2be12d77f003ecb8f21311e1b1c4e5822b8be9ba17faf36732f8df19fcc94df6fdd14544c7c9f6d023eb037f8e0083ccd8887ab605c1ee545a3a512469ea53f40cb187634c7848333d52730bd65492ad5338fd7d565f53e94e92c62d5e9bb06f5f9661e8acc2cac6038f9bebcf1969c0202c08f1306f01887e2f14dab291fa9180e612dbbe7b593a8c1ae1c77b9f95910aa434a4c73f76fb60e1f85cf3d527f323b82facfc8289428579cac13abe0b9725dc3927ef56266980990196e5a6dfe6b07f77bab8c096f477d0f14bb3352621777acab7f9bb68352652ce5494244527c39de72c217a335df47bba5d958775dbb8f8bed64a653fb89328662a6c34048df4e4d76bd9b5a74dda7e35bf2cd26711127aa06825ec7873260dbeac06c2ac863e5844422bac69d651c9830b7e075f8e20a9de87cdc5160693107b1c23994c9c8b9cc5565c006c719f3897d913c2c218f68cf52d753d32afb414e4bac5de8a831077907616f28686229a0268a0944353ea6fab9610bfbe4425c447cd9bf6d9bd773ea62036ec15404f2d966e8afe40b9cecf4642de4ef7790eb7cc4e4c181a68103e557fd7f15f31acebdbfe2155e0f89efd14e57fa2a644a3e1469198fa055d69bac4d87994b85e879eda81df4cc65799c818da3a64c600b75a8f622109394a47fc7ec604cc563bd69da78303099bf11e7a154830a10da38d48fe15c5dfa4bac5693c153d5797f02917c16e2460dddbedf5f0fdf710aa6eb25d2f94d25885fdd43fe0b52b1835f5861d0dab720c08bd9f41408de157fec28223cc6c147c5d29a8fc80c0b3292b8caa1550b1e8a83499eb8ad3308f6075a5d730903c2104b812097333e16312682dea27b0b068311ccd2101dd149f62ea83abebf50728b5d0bfee78d9358ec8c4c50f46df7e96bbd1873a9a5e0258eaaf90875cb8fb69a69a78af28488412c0fc36c9830127728b61aa4394598b1a3e0c75c0ad01bc2d4b8ad3397b83941a1dde58dd6a661095e62b215908839766829bb3c72e500a4589cf16438eec1b9cb5cb9117933cfd4773ee4697f5f6858fd4f2cdd8d4a03a00e8d0aee6cf2c267211f4971ff2e19df6cc0aee0454cbebbb625050eb892141f9ae0aa3ada241921b668091b92dd7aa1299d5134d105fc0077f5f67ff9ab80a01d110146c4f026bad1506661ea06c363c75a0c4c8e56ce006f45f5056c7f17bf1ce60027f48bbf0be657bfd96f5e97852511ff21417a8975f6ad1b9ed47cb6d8323b41243764ef7d63d33776c4b2a1c6a4677b988f932f60b31783b7d7d53d19910b83af9936d1e3fd42133a139b94490407707a2104dc204d28e0627746271ef0e07d5fd839433fcf548c2057bfc0f55f61983aa4cd2877790b97d8f2d24372952fb04335552bf0d1c761c70acc498cbc56493fe3c234f85e7a84a473a8ca6425436efe808b3e74bd3921ced5c3d7cce63e84a6006c4e601cf48414010c60cf6df8a8a85518a1c686b257fb5d4127ab7148402a11184;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h663499a6030837edba3e9bf329916330306e547ddf3ad3f4a0c7e0499579e60638a5f29ddbd89b20b2920f0717c0a513bb1f45b4392f4a3dec93f6490a4b40aef560bd8356d8457007c0dc786672b5e8f870f87da028d56da1988f18e3cec852764565b4a9c4ae450745615858086e2ad1ec1313a3e44a815c6d355687ec55c6f9e045c14926f277ee48c215e74bea990c1e5232ab84e356109fc7a115657da4c6301d395526f232564a0dca07e91e079f2650747d3ed99a5b32abdc25421f9664b2be4cfea3b45602308bdffaf52de34ecbf44cd50119fb9b81fd152f2258aaf0159f9e422c1056e1bb9137ac0bf11bac6d414c4cad26e2d8559e9377e7d52494c91ba93227ee27565c2f4eb5999dc60bbe6c2adb0ea8b4f3ea0ff35c3a5fd4eaee19056c5b7f17f51ad7dd3cc261db8fb16ff3b53793971ac14286a36455816e60e7346285ae1802fb2cb8d8c544580a9e5402256332c045785740ac99ec7231649ed30cc4b010d7242428fbf78afad618232b2bc650d00830ed18fe1990c88e7a4e06882d11510b661375f12ea10869029bbe983bc1b73f93ba410477a8a127f20e39ab99589f352f3dd06e00e79f6e15cd5fd55602d78fefa604b4c7ddf8363f5d78d2695e2964e25bdffb4e22c9becbb6e206c895fb1cff4d9f93d30b25177f2af4204e88ab63450082078751ed673cf83a5e2e8c258e440324ca8072ff9a032bb69a1dd4e27b7b8e8d6d0a1a3ac8361da2dd181c7e19cb876ee9bc81f145cd2c3a18172f19711b3ddf601674134ee38ccab527318952a9e19fe97019c6f89a1dd1b24f319b9c331bda2dd3d30e9521a7a69522ae432a6de3c98e11d5c8f4db9d4cada614b976f2295b197d14e1e3c6b10751cb7c2574b9a428f34d9998df8766352623f22c41bff5f52cc03dd1f3ab56856cc010c05737719d5884a83bf93201249adc8fdc44282670d401af48f3ca7502644f20f5e59080b630bd2479c0a1fa6aa15b4e477bb64f81add21c7edb14358ee6b58694d9497fefdee99fd216e59dff8012cc71d16433f991230bd33bf14de73b34a7d6c79e512fd7676d0c864c3faa499a53d3a1a4d04c435734bfbd43290ef1cf8f2382feb9c4dd5aae1030eb3aff55b5d7aa7c0ad2e910f25c37965d1ea1d360ba3b4c94d45775f6db67b63845c64d85b23eed8d73fb785f28be47b846f9c8d00e0308b7e0517264dd40d1d4acb998ea3030ebb38f75737a1fd989640da5f19dfc0e05830bcf98baf0856d8045cb5dcf6d733075687d4518df630f4c6c28383ee29281f032a172bba8f0adacb3ec7514ec0417d7956bdce73b5eb0884b706918f46e9030eec1aec381d04b3cefa70e3332207c734aedc8348efb95a28cf6f7545bdae046545a1280e3d8b19c73ca8c6aa090f249502dd89988a669af3880a7644d3a1414777a21443780961599e438e3e2ff877056de063b7987de047fd2d08d59a958042d273d264844567295cd6406713cb5c2f308e2cfe755a88daf778d4c2b767d884b2bef2077cd854caf1c08d5c013aa067ab33836b57cdb828321121fd6f8448d8acb81e1808d3ebb4d2bd935c74f1fd0a62bbec4bd17afed084c217561110382ec74477338b4ab8638cc0972ab595c0cd1c4e5a64b9d6be529aa5a26200241a0c2aa18c7bcecfcb83ac8c5ae137afd0561eef135c77c319ea9a248914592f712b5496c74386506e16e96712d426eafd4b4c8d74eaa4decdcae546c0d3c0dc6b0e15a0ac37f58418c868a0786b0445b7b108a9bec9f68da6b9a0fab9cc6a5e50c0201f9caaa26fd8169e7845901f59d703b38ff66d3a5e4306d145823e6602d97147825209a45d5a5c60dfa767ff27c57e7a3c403b23f407e1c74fdfcbe9dc1f737af730e3f548cdbcffdf2e134e87dbd5caa7d8349bcc2d527bf6fda124aab402c6bb51386b844a0d8da954dd510cb513a95bae2c45e43164bce61fbec3f918fb81a8c12b493f3b227bae20ce2982ee7a75f1087446da231ed44868e1fa55e2d4c4ca68830212ac94848c46a5ecdaf4b2b064a8f6f5a1f0bc115e2d8183b5e975c1065054a3b3f5ab57714a20442bdf99f4522cb31ca42f506e0227e42e8926b6fc821b49d5518008b7973cce790a6c07fce37dc455271d49ac93ab229b301a51c5501c1eb46a723c47d18d9814b0de97b1ea0aa7295a5328392fc6a59f4fd247299ef745f3817beae3251dcd2d0604cd9cd2a3ce13a2341df1183c100cbadca8c7f09e8347f94ab806d9669089c2cd6984405b16431eb9b5d8331112b24255ee1dfb206f0f2d5ff979c34bc7bb2673271ea96e9f878c8912d70cfd23ec89c66c2136c6c207d0e08728958a7e75de0cf815151e25db0f5ee1ac841c1108601e29c6fa71a958076443dbef6739dc359e30aeff3d7cea8274d25a345c822fbce62a3f3f502e61bb63394c6b82b05f1c2aab6b764cd89511a49900213a00455c8be14eabe22c57c0746bca3d4a3157fc5cdd32ba00bc2569bb2e0a5ee64bc360b3808ff9a682f0c3399525c591a872a50729201ed9e026030c4e08d37f784de0681c838f646d4843c493d9bf7ff59c008fb63d2c68a40fd542413d0fee0363e367ff254ddf71f2c93ad56c978c6365a1bf92cd147ccb2160c8b84d6c76d4f39fe8988d3af44cd758b5f7d10d1d3d42a6dea9147150a86cf0d7af66cab5b9fdc84bb54370104bbfd34c7a6f6c96b7ec0099059cd07330fadef7401fc5bcb499c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h51e2d9c98144e5d67151d50ee665146055a6a317286eaa55e5eed47a72aa0a33ce2e6923bd35cca2804c1495ad69f2b4b028e4d1457ad705283c41e1627934a1982f1e6e88c1f99ea1898d05e79957ad663e8bccbbaa84c17014ac94eafefb5b74421df485025e98051b032ef4b15ae5053838ce2452a3cda3a93b40353991707276fbc48a5abd86b386389352cbb4fe906801c23057533380f1fb1d977dcde5094c5339c7db7d72ec4baf21c3134259e1581c8db46c51509db8b2b0bfe2e7be070160964361b6a2f7bdc2cd4fedc2d967260ffa563d22e1339c43a7850269c80cf8aeaa63e5eeccd8e0e217a31d684b6a4f7e0bdb3e536f3a5f0af6d32ae7c04ce12fce669051f48a41f751b752857abba53fbafb08a852a74a0f2a418696b2909c9cabd8cdbe56555292c34fdeac65b4d9aa61b4628d56ed1bf18a1e4f6458ede2a02a52e8e577ff8e664c6be6030136414e8443506d63d7f0c7394e1e925374b5219d26f84fbd423f0eda78bfead9cb5ab8d56ae08eb273c9ee21bbdd08eebccf6543a4c1e5554379d492b2bba4e32646c504954e1141848360cb0959226efe4eb6513c94cfb758917e6bd969283f17bc2e83d302df3d8da85d886b8142e3f0e5cd816e2304cab9abd81367f49daa45592cf8791fa684d2676e6e1bd7fd265c705795ddea73dd3c48c91443bdbebffc5495e561f384e79c97fe7eb1ee974ff5a0af7b8b4852735c640e50996cf4c8078ac1f3bdfe1a45aaa42afe4a8157e38af8c808e8e7243fed9ee6037fc69d64ffce485d523fab167994bdff399dbe731abeb5a0511b0518cbd719d591469df7992ca8d1fa6b40bdd216c2ccd49a1a986ed4b6e526bc018a47befbb4f3c23e2b4bb3c706b4a26318a4085033ceb5c96adcbd0913273143200c39b11579ff491baedb1d52aea6c2da2064644b8989b6b0bcfb2a31990ffc84ec961855f51eaac65fe7813bf63252346ebeab125aa79839af3e4dbfccd919c17f6b31ca044c319fe6a7f7809ec7ad381297916ca6b1c757a34c58ce6885d89fd51488742bf85aae03f1b51f37018340ff601ef50459a18361c8e26290a00fbbd9dc3db56cabcdedb23c5d37ae12fdfaf0897fc79e4a6477ee53c083162226f7ddb7bef4acbae22a3c19a4cf5b5734ec9378947fe3d079c152c69dee13aeacfebea3801760bb65a23538db32f757ae942a4bfe907ff619ff8e3fb5ca0b53b15da0d3003f7eb5091e2b48950d2520a43af8e9ef1de221ebffd4eb06db5baa906ebe2f4e99fb12138ff963b6da92f75845024ce15bfac44337b0f933af4f10a3647ac7894ef93acf034c791bbac21119d00d0b00157f4862c74163feb95bd83c3a59c97ccc5296739ba9dd66c99db4c33c38cc36a6c693473599da525746cb65b326086dab76f8731537b7053b96c2f532d3b2341568af45e6ad183df4a1237e5d6b549f446ebe82339b8ccf8b42808451ab7f8528381c9a6765555946a067bb684bbf06076699c24f3a20e5ad2ef66e97678ee451850f8d5c6f4508ce17e4893a1ff521273f925914423341778042e55a8188fed28cc03954e11fb261099bf6e023a6a8f6d1716e2b6d292d23edb8d30d53a5bfe53beccac85b33e01974725c0ff8c5851a3bcb8f742fdbf8049a58f1caf89111ded6b1d6047c789dda9b96bbf81853342a3822148aadc9a4075cd57b5cb9040a8d96c220f20832a4d3484d38575b2e38ef87a3cabe6a21a77d07fea44b1c95645e2168464187b251097d388cc21fdddd9f4e29a11469237e53176a7db77368208694bddd2da70352aec9f022f865ec9716d2d8f1b9554c2ad27db949870a3a94511486e18878f7d3b0f56f781e69ff02d6aa6454480f316b6686607b47f40d598bb68e72079113a48a9ccf53bede3ce23594dc142668bf30de4c50fede6b7b185183560126927f2972381197dfe84d7dc1428569cc40345c81548a6ef7589aad66c97c737acf82bd1050ab6b470a1790a8cc87406d0b30e7b7f1cc1dd418ad1b89dfc8326cd4615c3a04c0ff7955c5c904ea860ffcb28f6621e5c3222ee4902deec02865a06d0d6e1174c0b5d758790ff49067098e0bc24bd0e75d85a853a72a4c5d219a959bdb58cd491d037519374b2713d3ddd9f5b61d01f7ac0c8b78efaf1d2fc369fa61660e32fe4e0eb1b941519f02141147f4e080bae9e4ccdc64780c4181bdad06843e3542b84f4c0682d4b99697eda2a6a5e376a20b1ce7f30e2713e5dc2d7afb88b748ba5799fecbf51b8547ddb2dcb2acd9010ae7a73639b9730327dbde82e0d903e098ab96376e0cc26a054892e0766d514c5eb8ffc20f6835ae4c3d0e76bc6de141a2ac224486a35454fe61c681c257af31293bf1a944c41275cc737b34916d92615465bd0988ea6f4e1b45784e5c90e4e48560dd73f4863070e1fe9ccd62b4bf67b39fba2a7350992823574b1b1d074cf02ce73ea12f8217bf715bd6592c3c6de2ecacf097fcb1b75dfa2c31eb16f8ed0c11541564bd09635dcf3a45b770333378807be81e7a3cd0153d632ec17020563baae020f499d6256769554a6121503258868bfa7f2c05ec777bb4c05a0ae75e741ebc12fa9b2e63bd5941bf569b0b2360890041f9fb4690733b7a0d7b86ec9836228cc1cce8d059c8bd9d84d5672f709a37e173863a12ade4088a702c1e9850261f590619debd299e696ab03176cda0af9369b976747b05871ae6ce4c631a8d7491cdfa1dbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h29e2c6c98d81759b5c6e2632290467e29fc1534f2e4d8c8180a873e3ab29021a570cc3130257f2b08d7a98e9bdd507ab5c66d6d50ba7575baf762c7157ab11bc69ab4bd2a0036afefb3a60062cb9980bfc2b2d7bba8adbe36615e913407016d7ce339c6203fce147458294c08e067b25cffe4cd65e2e002532f10afadba96731c70130460fe073cead3baa6437204a720504eb84db3b4ec8c5fcebfb3578377609959fd8c42a9c13a2cb8621f2a77978dd0efccc91041a6af21a01f0de64be936f39880c26eaf669fb912c32b65833d72c9c1121fa2e302b60610c6c3d0b2525ee8b9decb284b87aa2614a733a4dbacd2a4f0bbcb8f774759c69f2cfbdd4020b3c20ec2938ec6556172fe5e1328a35a6824a4c118f3b887569cd5b330e05babbcdd9db68846209303274dd6e2da7ef12c2dd17268212e984f18806ecd32b010fe6a4a79a7927098396c249bc3feb282d9b0ff0d200f7afcf88f9a5634b86dc84ff1631831e22821f0b064b240897b95a9e17da9b663f0f97042272d644bc30afe00bc7d4e08b1b19f7f1bd572d9b9ca1fabf880084519e8a14c10f1fd2f1a93bc2877c9a58672f4743eade252994600ea013b7610045ce19090f0ac914ff2d891b0e64d0048eba51d45422938cff1cbaff89c9a8940a3479558b2245b31b7bee4c6f844810dbd38ad915c67c8b0cbfc5daa063e20cf07cac738dba0458ffa8f1fc0c62266373fb500360132aa059372f032a816e0cd227f7e3b0406bde89b539a29391004637dc5e64084abc336087c709d8c9a126c34f706bee647137c8ad965bd0600bd415395757fde93019151f08e4e4fd51348e1aeba4d242fafb7c8e8c2ed5d3489a3314107c876ed16a8553efdd46209db5e6ee258af156e210c71f5adf2a0195f1eaafb2a29a42e04d462df05c97bb37002cfddd4526785837b4c6cbe802cf6bbc9dafdb683fc228dde6eeb5557621c3b6235318f45accfb39ef934a9f8e16879897b4c7cca9606158ff4d90f0ccb2d7febbeeacc4530ecc33fe77e0b1768c23f939538563a47450746f0f08400013ae0f3efed5151fd1641439a2f54386d21411267e3d62292b507cdab053829718a71f1410d51888ec613d7cb5be9e8e98d3d1ed5a3ab1a65297528c8bd1bf99d74603d4dafce6263544e3006cee968f48b6e6085c9496cbbd7e3f690a25ebb519cc0ce4df27311aebd261b73c8ab12bd15f6b772eab47a5ea463386c0f62650b2bb8d4adfd72862b350f2183eb37e52fc34a994fb87f43b5d3606a2c31f6eeeafc39fba4d539e75916bab21bd838469ba7114551ebba3f15fc3aacbd012227f49469cdcc7cfe50ec411cab7ff05a1f69bd7e7aca359032bbd75f23baafec82640a35fdd1ecc3b19193c33b88dd602f1016a414d77320a1e60ddb2b51df4f0617e844b65680501ef883c83903578847955ac7de6c79960b1a17db995239e98e669af17535ff56a75badc470d2777c4ffa0192564457e04448064996440d9e129d17e605fa61dd1e2dd15e8c415d9f4b06a327a3f561412ea9cfe57a620cd949b993b619d1b2f2073c5d2de082cecf803bc6588685913a82d17fbca37707ad135250fb07b87baf0e3a285bf11f8979b5c7e24afbfb25ee0702a4617b87951dd8b0a81a62a3d4f95b0833c19308c7f533c1ceb023b86e85ea19c3c6b70b03d68c1602487c669aca94ef8a7fa58933b1d21cad4b11f514e29c21ffab1827828d427eac4357ec5f686e26d0c72ac2f6e143e4704571c91bb8d96f232f89f92541512804115fc78d470c9fd100354d7b29384ba9a1758f0d324fbcec113c2b76fd5fdaf3c50bf73faa8da62df8360cfb719269af0c1debf1eb1fe27976318ee475c8f6a6265a53f7362356799c1ec0102db0ceb3cb94826e04e8aa3a514d9aed7eebf7983bd96f5865555215c39122b99ab0048c62c21f0d0dace6e2b4919ddf4853b8276ef880dad944c6066852f26935348f94462aa739fbf5106c1f4adbbd9da11efcfabeded6c4bab4c12a28068573ce7eefb9509ee7c25809f8d5237f9421ad8f290891d88dbcde39918de060545927e8e038377b02ee6447a316cddc72a4db75362315d0d888fd943152a881af17bdf4e920cd664ee5abc8e7388588e9d5a17dcdb16aa40ce7ec1cece4d1fa76bd87a54e2265ac203e83099dc466480a1ef7439772339c7f3659e4e8dcfafa68cbfec5cb54396d9cced7b804fb364d27e6a07359ae59ddeb620b6bbd80befc5a5f2890e16f88ed93c6ed1e8f9253a229240d3813c249c18b5d07d19089fe60c48d94dfe3529816021ee3d7000c70e925134f993cf1dc710df58bf0ce9b8618dd1a6bfb4a7c5c877386dc0ee6ac7eb1d7d87c5b20a3d7969b98ea1176d00661e8900fb4b3b8a0714138ac6fd948511d52f5e5cb5d564adf3f90c12c4a1eb5d519665e1896a18535d8dd525fa244971e32fd7dc55e56cd88c93eb17de44caaa452d5b04b973cf6e93f7872752a810515db5b1d8bc62858c800e844e3f3ebca6327e708ae37a261dd01aa0d90cbbf93b5236bde4c3493a0f4520d038f48fdf5d6d864a746755d73ede66f43a85038d9512c8b62a406be3376a3f4cbaa5cacd418817006dcbe15cf78bf324d4e896d529f867ae541f214843f4a5f44386325d9a25daf83fa8870440aaa9bd054dbdc4277ed388e361df7a5a27d886c53ad49775b21eed05640e3f00821996b9184db4c864b2a6d032bc9a01ff97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3ba49f06811c64b3991d3f8ab0ed2070fc9cb28ef3a38b41c88bd9dd13a898812dc3feef582b26d913e4c80b4fe91fcffe2d49b64a6010c2608f870cb7ae507cc0ee957fa2bc9b429e395f08f268b3d06ca7f38326779ae93912580596e3074c3cf154a4a9496c083b1d698fa84f6e5aa367c65f13851fbde5d738f60043d3477ca63d9f8dfb34b57caf2bab9457d82918d7373f9298aa42a35b983d423fbc31214501dd1156abf03c794817380077a2146adf67b31eb8b9f665d3ee492ba9ae05ae7dcb9aa89746cc627ce42675467f86f05b6ab6bf8b570a5906a3ba4eba7c8030cd7e3d99158f8b5184b2a1b2dd55c10adf2f38112f2e67602117f512ada9e3a8a87cd1bbf329e6cc8a93b21c414fcaddb1f4e558525ef3836f05349c6ac204646c82dee93ccc53b94603549643c09f56349ecfdfa8aede12467399ac8417044cf743c78668928e9c4195db9694e7d510b17003c69b10d6334b4f043daa27a83e66cdbb5a37b8d06724864be17c883c3e640546a0b734cc0a676c6eb8dd1185e6bdad69de73b102b9fd2cad047c49ceda527d1fc76b3a2ee275cd7cb93de2a8992d9ff646830c0184454c440e82d9b224ed7976ea39323253fe3c6b4875f7f1d32fb7a71d517ee112470410f5702f0e9bee571cc452603f75476004322fae460fd8b6029ac25d3323a8fc301e04511884e9bc03a3166d5918a05c5f21623da730fded2d6ccba3fec18e6a4dadd83d8dd960239e0f8260a8495fc47cccc1a17e6f8431d6d503c65aff0c08837a79217b5e59320241a763d0778ab8585af3e5347342366eaa259f075472b2d26c57ef2eb9394d9c01b13be2fe49f4af3d9ccfe848c3507be283e69b8be2acbd901c364c400eeea49b883a75876f7accfa25bffd3240988b7266814db0890ae35f9401c25fb47fa548137a9745be3be229b84914b959c7ac77e043a2658e8d01aeeea3663bf9574a5c8c805f286ab7f926032ba01ecb4c358dda5b0860188708853188fc987bcf76440c713c027987cc0a2fd85b2be0dff8dd67be45f7d7612b6367270823c57cefd06c6fb2b4680059ab79f2eec3576387621fd3f217647cda6d6d4dcf8b4753dfcbb56a0c16a19764ffc5bdc2126b4d503a4e19c369b5afa8a8b3ab73b4c09e868f4c8820315e65fe8a0c798622623524748694afdb70ed5c752a22c5fb2069efa7f5e12148bf306ffbb4dea2474b0b5e3bc743572d38f596c6852eedd5b975d6766dec5cf4f0ed2107e07b02c98b75702d5fb6c809d9ffd77611e0b6460e05b4e3a5e325bdf0220127bdcb78623ad19e0906f1a6fa29ae6dc91d1b02f8778da9410905e870cbcfb8f0f77c96008977bc9a2127196c1725cc9b675c8c87f9cbb941476704e6ae1da8b5b861a8a658ba43a03c4fddc535b9ea269ab7382c71b503149667864e72ca7d5df61135d41d4239c25f3bd7751fd0c7d0c47ef33703311a5bf7c53bb83b7dbe992163042f14a71078400ad0e1ef17890b6a7c7a52958999f26d59278494549e8856e4f8bb02514a65c24b058c3781b367c88ffad9bc364e19b32fcb9ed0ccef16fc0db04165acada938c7471e0a152c669a51dd02d8daf3a6a2ab94f32bbe7014baa052977a077c46623fa9aeffb6b2de6ad081d8b51839f0bfa309aba9d21e135097dd0fc44667a488639445616377aca3ba55b069112ad070765ed84b25ff0b0010ccd2c3e2908596553a96276ae37e55455b671d587a8a1dced4bad4e704d4641fd8f0d2df30a87e4dc1bb6255a99f7f75384fd24575e6b1fa8c6521f22172f0233d5d449c046db38eaac782224737ed25381056dcf80415dc197c514e1dce475d47a5315e900ca516ba68828250b222c055ceca37824923e9f5bf798de0403d7c14cd1cafec3ceb93d1b857d7ded6d11d66bbaae7f4c167dd1724487ee58e50dc96ce2dc5dfee5fec4e5087b1985f79fb1a74455f2245044d2b2d0de958876ebef7177b59b912783e5f0d01250c39837583023aa201d68c55dc3fef19f8ed11bdf3c246965884bb48550b716d716ae9ff54ab569d8e21641d81282a27ffa48342188f7074861add0de78a5d6fbc5c4d06bc0399b8a374b9427a82c16f2d63e19a5730ea6c1800b5553646f0b17990d79fe62cf1444c601fb2c4a4e4adaff0257aef2f81f5f97b0b6dc5144e1d2e38ac018286be4f15ff3fd315e5e49f3b28322897b3dbe39a6fe90b370692947c26c02ecd7226c6d17cf80e42ffc4535d249c7f8179d25db3618fb6f1594996c65606529026ac0f8dd1f1c93234d5dde837886f83c04705d6892e7d20c106995997938d5b58549d56c8b8d875d8b9cf8438ced22632b8bd3a6b760300e7b49f0b41f95664a8cd9cb9cdde37e3f91828d54e8f0267550cc03f8c82b2341db579b85c93a8b57f8ad892420d6f83c634c094725179ea01f753948bc90f55a6611c8bfb51c0526a12ff2b858cffdfbf81892cc287bba7ad184d4063f880ef47b65488338794d4e9bd2d89052bfc895ba8797eb701c8c84a1921b58759cd3c32da8da97a21f83249327987c8983921215e1b8bc4a7bf297272c9d0ee0046430a506b0655805b2ee12b3b22f8417ee61721ebce7d1022e71d1af4c17bbc75d97706bd646e249e3292b0c16f2573d946f5134284ecde378e853124aa64e5cb4093517ed73e4b22e51235692556fb3cc5af40808dee7510a0a7345524f6dc58cfe4bc85f4ec90626ba34777e0e97eb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h517b5ef698f9b79b1f373c2d1cd45dda504c9d3e07747a8e4630fe03846baf7f6ba8c5b6a193d72548f69769b99204b15dd39311de05f74d036dace6f1c2b05756736628480a82c1b6d45234bcd81119061ec9d01baafbe99581f25edb2e2ae2ce4e407092fc9348918e43c29dbe47c6b38b36732387e5db66fcca7f8f1a9931701120f3b93154a5df887cbc6a9b16e2cf3fd938098e55b1ec70e9ecc214a6714e9486fd91a5e4c7bb4dbf9e4f2a54b8415b70b64b1da035fd9d8c6aca448605ea172cd42b15077e41bcd1dcdbc357383dd993b622fe23189f873558e560a17135f728ebf7f30b00bf73810e8448456e9c255748868cfad491f2b0d2ba15cbe16d7145e383310651246dc811fef507812f38b107655d2eb0c0d9907557ddaa3c24e42e0a0009c0a7fc8618c1a27eed8b809c80505f7d2ff5672f70747b5eac8b033c3713c5d12b8a350e0a3ba8b88822556651c922ed98ad28ccc2e42116592ef03654ca8a1c14e3991252447faee7025f648a9501f5488131b2be9eab38c25d2aefc117e42aa000537df4a21fa5bc43389224363794dcf13ff9febf69372d96ed59be022e380ba038be505437ed06261f0dcd98d271ab77f61c9e2809b48962c498302822eecafbbb2f8cb42aaf010575a3cd775ac42e27cd9598eb7f7c22a11cefafb0dd93a5b2a9b189c0d99f6ab5b002acb7461c2883142ee2b334cdbca8036892e09c9fa2ffbfac9ef51e58070c5c84a76e8dc47d5c7efd2bffa381f8c569a9d466c9d61e9a7dcb3051aec3bf6f3f602685dd4ea09f85d6d38d1c2cdc57d4fd5c4be34d5c16747723e8343fc069fc4158081fb917fad196ca8b5c4eb4bc32a64a92229950846ba007f2fddc291f624744a2eb1540459d6b25e15aa7c3d1fe7abd3a6f0fb31e4a01eb8ebea4abfeccd1c6f8291ac06f067e44046403110172ad69d668173c5b8d181d0ea4557b64e56436b5347da0f26cd76761f77e185fd7ad267d45fd8433222ab136e732a8935664ba0b7430fb762ad329689ce585cea808b4b3825a880e5404587e643e02c365d95c31a9998d99b2566643d1af9745530db2c55b52324622d9856975cb603017ad703dd9b6bf3b7844ee5b59f021154d06bfd75e1904651da46933469070fd93302a1848a01fc5881c1e6e2b10308be21f5dac076ef7637ddadf20ce63789113156eb2e64c6601da62b5559d3e30780538e8cbbe7adccf9f98eb6f8786d737afd20e98411b777ad9e16feaf17ec74e11ce7ed428fb9b688aa527300632960e1260611dd2fe57afc458578218d00a17849e339429b5b713d603abe32a304998d19d25110179006a2ffaab4b3b5da62694d5095ba0cb2d664c1b1cd69dbab4ad6e5117801ca828341eb9753da5d194b2015b2bc854ce00abf87fb8b16dbe49463e681417622dc6ebbcbec1d549438f37da51b63f6bc62ac924a0f75da8925f41bec1857296991a46886b5a4c3a557cc00f52d2bbdc2b5a891034ce5847b0c05d621bf2c8f3708f786b8b801ebddeabe2ecae5037e1f7a1e4c1c8cae245e15b595b14d4ac1a52dcd42653ad9e8c0005d3f118a3fb88300bd50a81cd4785e3cbaa21ba3fd3eb58b491434d41e95c910a587ffab609af75984a729a76d2effcee0b7bf71e7a26c6acf993c3ea74da459986e7faf6f153ebcfd8acea10dc764f11ccc1e9d52ae259bf3405a33355907c9c7974acb3eab0e1fc026aecad311323b2505f9b56037f502e6679d1e4611ac25ddf16e04c5ff535cf98b480638904a2c83111b81993ec4aab576ceec64b754eda97dfc7178730b03df74209b7c510b3a3e90997f0af4763624fd7d0f9c94cb241b40b488aa4a1e62ebbdbc5fdcb45409a539f1d62fcc068d4e946653930b48fda2479065789fcc8f1d6f07dd0c1934659766dd704144e3c677d64f04050535e6095516f4161f67eada5683964e305500025ff83d4a8d826182b442a2440afafe944a304a56f17810bc55abdfeb14cc76676993e433c2ded9a633fbaeeb45ccc35dfd2598b79e506f948df0fe02470469033ce3b55ffd6f5be430821420bd0e94f77d70588e1c23a3a164b1db300226d89b280b10d550cecdecebc932a3d678cdafe85b7a02175808a1f8f10645f67dcdb2366076d30dd3a08e77cfd79734b45811c9120ccb203333f1b50232fd7bea19eb99ad4ca31037f29f44cfea99c25d018c7e4380f326a89f1641e8df9f1cef0d57b87e3e6924985c593bb63a8d9ce38c5ba504e83a38f52fc3197aa98a2f5bda153069a2810946d86bd93cdab5fab20a1f9fb01b7959591415b96f43e680ff81af5a239c375435d144ca076c3947833e46474c1a0389a4d356334b96c86463f96e09220d8190784b0b4679041553edbb21dec137dc0d90a2f45d94c5882c7a6209b1f6d0949f9243337ac4c5742c9ec11aca63d89a193232d2b748da25754dea1fd1d1e9136bb28e1e224256d0621e42f0597762a92cbc750f832f501be64b946796dcd1306b1d952e41ef04e5722ccef958f82546d12068b66bcd452f02175bb3ff683269ec33b24fe78f358abff5cd846f93c07ba6cc8e02c125d785390dae326b7ffa13ed0b0d05f29180bd8622c2201b8dfbadec518f16c636d64582744b469eb545ae56d06eba6e23605d8ebbbf4667b99c279b0f2d6e3f96288b05d574aacd0a09fb10a0513a8a6736933e8dee70f02cf7ba3a55024494bbe01085ec33ede3cc81cbf931ac68c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9bb9097cac37808ab83dc263022391d0dc1f55162d90ab30109c73ec659d85b11889afa1ddecdc702649ca28645f343deaf0ab12c4df0e0049cafc3559e1fdac73d5e772d620506a02d2af238fb619bef4c279241c4346186adf296b5d95bb8ed3b612d995e4647191fe1ea30494ec9455e6de8a33379141339200acad55002b1a856b9db1238e33d5f93c86cb107f1c40eb977022ca29f1cbbad425c7d77757e33199fc775af53eaf7e5d133a671874b2c7c9bca0087230c5cb5fc65598f803876e82a1e88290e5c41aa97e14d933d5f241e1a1e1dde09bc6e3fce15c5455a1ccb092b8938ace89b7bff194c4d04de53a35e2134f178a1daa141710478c82ff7b5983d3502a8f4c75681f21dfec322183388f8230a4b5b6067679435b5dbf33dbf3c5f12c036b358e1bb917f2adfbe58887765f327351525859f04f7bf72dead047ba25c1e047f2a141d8260827242d47bc0182ceb12b7448a8eff79b58974c6c31e3ce86e95918659c6f0fe0361b1533f32c8a507f506c249efc15d3cd01eebff83dc2712ec2a2236942061c061287971af504ef66de3e314edb7272b5ca57c8d7e5dc74b2d1ad28e058c61b1f53ecf10ebd195d140eb292fbc9b2d12244a9f88e5bc5e32ea51e66b2dc185591badfc27efc89ab24b5a8e5545439d13fce91e84bbb92641c2d5a951630fe69d4f3cb4c78168107a32e60f9adf33b5bf7fe135fdcffb3cba4075c1986cb4876226b3fc3fc8aafcd2589e7ddafd39a36904c555b0874a70775be184c38474672c88d98c3fa7f73b54cc3336b1364d324ec8ea21bffb624c14ef356d43844579b84cc9ec9fd2078ce45b64ee05fb54de2ad1db70cfc419a24ee0e8255f76b116cf497bc5cd6ba4b1268600fef7e0152686f5cc7134dc4d5f46207466a9cc7d860de2f7cb07308f85550aa27264252ef11ef8c0b8879778a46eb7d7dd40f75b6c6b114616d5c47a7e30bb5dde36460993cd04984f81e912e5ad762dd50261326c3ab7535983c7cf5bf7e14af97750c9a9687ee2d3fa21ac4667ae188a65d5a4cfb49ee1d7563ffc73995a04ff9e2ebe8a9a3711ef50a6a1a06cf5929c7992f68d86120ed339abe9e1c1d1acf736e6cb8a4174e0b31d2a0a70de646e38f0bd07b47f7cf9d72cf23edc177f583afcddb5e46e4151eb5e819022153de2d8e2902b708046bfc4c55dbcc16bc97893c727a1ec654225bf219d7a88fe175b76db9be693076f9ccc00f8705d51f4672e9fbbbbb13c73fcdcedd5e8df30a311ceab5d0bf03c91c2f0f37a7fd0595c711a210b33a4b2fc47dafaeb15984fb13896a236bb9d0e07401c1e4ad199ed566353c244859815b933dc906807ca4ca8182a1900eee44dd3024aea93f90a9d31aa7d5c7c95ffdb02ce8a7ebf5b259117d4c8e7239cb681a54608d7b763130125e962a2c459840875034f318ec1e7ac6a1bd5ec6988f294975d903ed242fede8e8ef9236fc2da3fd040a19f7a8887d4e52b217d0319605059973d71a93c102f447af1a94f86e0d3c00420b643756331f869d6030ec9bf8fb0b155bae192b935fe7d05f755dd8eaec34e986547746bbb82615186adcb92e5f788034dfd1950a9c4df3dfefa50b2811fcb8b7bc70556ad99acf9a64d671c30dde0d81466a261673f103b13fb830559f884194401670c5626ff20c8e8620a8a3d639f3380ba7429c2ad44b89c521d542e9d5cda4f0a766763a2b2a228a8dc35f5e28f879447c160046bbf0b681abdd43b9c251a1f22eefa1db35f7de40ec3e25c3d812ee347b12eab45eeb60e7c83c6d89a6ee0bdf301a97e5ddf268f21f68530db1f804b69ec59a8c4b3b0b7fce1699005f87489c6652a14bdaed1d258591fe7c2126cdc7d17353bdc2ad02674a152107188598bfd757db45731a0e0c482e4b4b72abfdd9e6de5c18f40f517872fd69bfca7e9fa2bff8cd18a2f6faa55afcb4a371b1e4d971d46162d9778362e52cd53e027fddd78ffa4f5a6847d07570b594d45674d40bc8cfb3aeaff7e66fd6de9dbc199c8cad5f30f518b2576dc669aa57ed37920013c9c945ea18eda5f25a8ec7e001b3d7bfb55f456e0ab080ac10adeb4c7649ef449b80bc3a0cb024d2d6648d5dba9e0d01f6db3a8ac0187d25f4d4ce7eade48e77d845b29273e207a3fa1a53ff204b3ca1b7498b3be405ad20b5f8cc2d3bba65b1d6e18d5426bcb97ec3ce2c648e402c042991911e0ccbb2ff2fdabaf153a37075cfcd2948bae82b35c2ea289fc876d7e4f3ac3c7e4c23e5cf778c1df11da558b11476cbe0c0775458c61658d99bd1ea766889bc399053a9cd843f13421a0b46b6ea9fbf231e0399528b09fffc4c5c4e907bacb260abf0c9bf41efc935111fcc6c880f0db450712cfab6f4c7945d14e2a300df76dbaabd26074de0fbc0099016eaa41ce5e22672afb5d8c6212c6f599a000835ae8870540cee4c031407e9b4176aa8429942e476b808abbdb9975a8af27a423ba731ce515aef0f50c0d0494332e8d1a307a900b5dc13c501c32c464f5a3926c7da941eb9983d2c45b2fa61abb6b23eeeeb639b2900580c0031fe0df927950b0cdfcd0139cfc16a5691cccff5502eaf7ce4ef2b31eee49661aa6ff6e4b44b17ff6e4b0e3c2f6de7e37c1b440fe8487cc56c70dc6a3e6ff65216b6a7037bb2d0533f9f8e4c844d4aef3daf7ad3f84094281b0d3761e13f9fa285ffc5b6e85634c6912b26ca9ce3e28c09e5c428c1315fb9619f86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hefce45dcb78ae47fd107d22bdd730fb1b69f37de88d4dea0bf1df3d4602c575505efb9ac3abec8bfb4c4dda9513d3de400a5acafe283167c59635c04758540392fe4392dc773cf6b0da3b36f23c388b9bf2ee1189ef4a81a4e92e3d801778a9b92263dcc28db070e0573d528fee1b33d06f9be17866b7b01f238a43f7b703d82b34ec7abd6ed7264546f501831fee63a202636f38dba5818e7b107f04d13e546841f16e4a39e9c79c939a0de27c22c368bedb0969302260885b59d1de0e101316730cf35f01bf5e9888ac8f51480c09c6f239f990c347b7d0907d60826b25aaa00bf5922e2c1269b08d75299f3d55802a297326c7e13b30ee893ba4ae3ee66d5936cfbc136e8accb70b2e1f3364cede74ada92c6ab3a487ba2751d89e65445736d1d1618c393404d83e4e39be7f67703d9f1002fa1c57612d89c59dc60049c682c23f0adc206aaae69ac1b47f424abeac4033d1dd960aeaec6c78f36fd7122945672d1739e8315a034ea645a24b589a6df65aaa52909708e7e46f17c1eb7561c301ad989e6b298fec0e85ccd5e27885f3fb977a12d48b2e7ba25c752b3aec9ee1f2ea8937d43e45983232766579b5e6a813176ca43353f4dfd8f124ea1d52fa0b94b0fdc9dfe7d596d960f2a7bc29e24243c15cc638fb4e03b9e6bea9f150abba1c3145d6eb567be15e0ba8a7a59c81134a404f3c57b3b8707b9160c26d36de15919c05816b2b5ff8b47b7826f6b1d0556426dede68a94af5d1bebdcba92708b77293648981d06952bd9fcf927b02135da9aee4c112809fe53db0a56ec83bcd7bc599dbac82ffe4e48b1f0767daa06f045a5e63b606128e9957f844a234ceca8f6dec3cba59eef25058ddc23b8f513c7069a364798f88450da353ffe50b44b642a3d62f82a371197a6541835d7526701ed6e0aa5b544f2e86279e32cd028e4e4122b23f1ac469f9ef7ecc8b8435cbef1833f04fc53c795ac187a45435874bd2fe5dc29cbadec1fead66740d2210dcea0cc29d019fabeae6ad1712f9ae961c3c603443fc3821380d010b6e417a60230f0567a7d7dba6f3f88535adf127db7ebc3e339f852a6529f9ba666bd9932f5cbe4dda988aa016418dc3318d1f2a951d125ce39ebc8801def04c75f7b968a302f6744f1a6223256fe7d2ab5c2f5761c98a77a8c75b7b39ae0fe23e1a896006d386ace8a437a1f805fb5a64fcac3d4cfd368a6f90505b6cae7bff80aed357f74756b41a7138d2529f60c431752c75588b26dbd8f6c9dbcc8b5ec71a3ecaac35dcd7e9eb23e622a93fccc2608dd8265fa069f2cff24f022487bf2d56b295706723f58079e0b0867ac19f0b166a3dd952b4c6379b6c85d4dd01e6be1b346d21680bd67e32e36425ab7dd833badd62d06d9b4d15dca2127361bedde1e4ba374758b34c4b7c8c28a3782a0754b01e69ec19b51ce954d089bf71dcc11391f7a154dc8b837ae55b76c28a7387db0f2aa456e1afdd28122f8d40c1cac3839855a3520e1f756f9e22d80801d144f0c836341f5350e75d26e47e3723c4c56445f1610c8fedce7ed398c9c5f7b076fe4972961bae4fcd0f0fd73401e3e88eb86386a06a9ddbdfb9df538bb1634ddd12eae62d5f6fe8118fe6dd153471b64ae6e6f1d7656672a354cba8b9ee10073a52c1b775d912239a1f20e2c796a3dc563358885d32084275d01130360de500a32f9d2e1f8b0b021d309416cce8e0127fe3f8ba5f3e262ad3beb77e50d3e5b89129277c3c2a5e174b6a7a0cc90396dfb6d832ed38e9c6d25534cbc5642c872267e3f906fed49b4f1cb182228215784d1cc37c2bbf7d17a2066df521bb22a43cfd2c5c2f645debfb215058ae4c4c76d1d0b26ded66152bc11f17114439f2f0087c7cf167a5ec26f8cc833e0ddda2c06f2d2573e5f09aa6c4c896ac46f956cbc113554cff809f1749d97462342083b2c4ee480c45a1d48c3640d418c1e46517688103b8365214cc67e2ca0094ee71151c753f47b2b2a94c4974d7b7def1e56a5cb64bd3bc43a11b9cdfcbdd313fcf9f9d54fc157ce7dbc4fcb075ac440e795ecf4209c5f2be0ece56fc0d9060fc30384de2fcb94d1113128cc10d8f1a9446c2950944a19a7ca01cc48f7fc93fc9c2d14b73737de9e4126f7caabd3b4f175a277b4c94e6111a98452edd73e12c2e47236081283712c69ef8ac5fa8c51802dacd9115530472df7f34d3eb2c65345811acb67f6139cb46121ee159afd461e3efaa4ffcc2573ebe192835dc61cf3f57bb729d893aa31ea59f991f882b6ee6ad1e03ac58d58c9e266d5f673fc14541d7430230d034560e7bdb0f3d9a5fa24b2aa3d72e8c362435a77e847ca096cef62fa22c729ec3e02be8bee7f5edfe675cf63d4dec0f970370960f3aa4d66aac3f4cc0c4f172ebdfdb66806bdd10a6318b53cfc5ab6ac3aecea73b38b4ab82b7a7517e38d063816777645eb315a6465d677ce6f134d0e1057321efc21daae7968b663d193e16b633f38fc37bc95dc9b19bc6972277765e7cfb3d0811f9cbca18979ada9d3df79857bd12ebc316c2367458d8010b7ab6a1e8ffe61a65ae05276016b30761d93ab1a82e191c6828f51033a2c70e5f8ea4dd0838d4c5e4292259b807f248e7807b36365044cbf161bbfcc23eb9d8211d22048a8772eea52a8601762224811d02e98fbc03e7a2cd01e3465c410634e34771b461b9af0b24fa3d0b5d760417ed0517fbb250ea3d982f5729f8ddb8b953798ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h30800dc7218f50ffe550c26c0c3d8bc9834d2a616c9e872500938239255476a394f89b8ccb70c686cd979b82bc0b2015d2cea5187c16a721c7d62ddf60c5d1e4720c8be94f1d1f5166ee35f9663b6e858f4e6cc3bc4dfe6648d0da65d913c49c62cc435559e9123184cd9277b05feaf7faf049e41ba802a0a18065dcd470072dddb93af408a565911c8b8619972ccd93139e7cd772c335ade517a206c9d5a20475b822e04a1ad7dcaa995394c9cfe64c08365efa2ae2dc9112a2f3d2d7696f2a99b98bafa37d6eec3f8d219b9eb1c663dfa389f36d551bce1efa175a6ac1fb6ad87df934c2e7fd1f517712ca04f353a4e30ad2421a84cf6e19c899602916f53e1daea0cb394862ae628c76219e4bed11b8331066481b6e3aea2eb1141f54399d5e2b6fda58a6d34ac25c64c1fc8020027a9b3065172fc8cfb3eb02c7fa8e3438f095053f8c12ea071f2720d2f91205133ef15084b2e406bf5c84cc3058cb43507dee1f614d9234ffbb12708f6abf307480862dcaa650d6d3ebc474d1cede26ae62b3e2217b0f689324dcb5d97a302bb99c03e3b08fa585adfb82b240b92be19a5b17f88521422aaed8b9ac898b33cc42ad5df94f25aea80880fc7938676283c1cbd524cb7c14815fb0c869ac3f5788b5c4b90bb06d4d8f038b04d11bb9f8bc6502bcf80ca5d0f585c721bdc2cce929fca3ff328a9ffd9123d38fc03d45fc9274a93d32fb1a429a7f445c130c010643f0665f0bbdc09d9101570d1a74c402f37857ea737aaa1f234c5428907c36356ba996da9fcac40726fc827ef790e39194ca647a40e3c37a7372818562f5ba0b6248fccaa4979aad1fa51f21b84d2ffff8b335185027a7676376018e25cd370a8ea7c4241264cea943c72ae20626ec8f18561e5a38629d5295b80a4f50c3202fd301c7251d37fdc2e9b15c90f88bc9c88712eeef5f380225401e745b8349b666fdfb42f1bcc73b60af3b0b4ada384412afc46fa3af0b5c500efd40fa56976979cc40ac3d4247dd0d61f2a7e65e74cb75be993c73c35d31b692c3eb2ff08b8628d4109d0605368f2408b3c10f8311797752deadab776d10faaf0d45b5a45dd9d134b0914e9d22e4d54f10046bc76c0593dfb945d4242bae9c5b930e528f3be907578b0510fd4b50e97b74b7fa56f377f89a9725e4bd1a43fce45d663a08768d4a92791ade94e8af33e638101462995cc7f924027a48db40d32d52af65f13e5ebb5879c60fd990368bff7ff105799455a2d3340e783fc52dc9869af7f826a83e9aee2e7c70ef4672be41c9f96826bbc7cb231897ef3fe82c3d46aa1dc0826891a16939ff1a8ccb688a520f7dcf85d8c09a25791ca1af8ed078a319bdbc8c8e9c92147b302b23b444f9834052ec7d21451ac5909e47367877b7b9520807f886fc502d5e2c57128b2e8d8b44736cc34b6529653555366d4f4f8243f8cf08fc385de4c09f9e65e45a7220534a360a7da4fbdbe128256d98acaa0cdabccebd7639455c69e0c5495af957f2c745b0b47a6351e3355060c29d5f062d18f1e2aa8584a4943b1aeea93f2e36b9e446175efe5a2f08ff2cc64da0d6b0cde35760bdd13e2b942d29eb9d7b742ea4202a02bf58ac6888ea9a475f87f177112c70ff140c1572494bcb681d568abc7b7accc010c3e5755bbb880e5e73542465e29116b02d74c94d70189cd2158a8b32e859ab88e4dc6f55c97037e66e0dd56618a9ae91ac1b910da73fe733e926941f9fcbdaa98bee93b57e3a1ac0ccf724f93675470947c9404a276dab5fd42d290837ca13167df01cb70f1268635f8f7cb580e468c8d646ede263b65a51930ad86ae9638276586c3aa12def05c187b30d8deb8be2d75c184625020c3367658cd04796ff947f8fa6617f281a7ddadc5f16840e56925095b5e48cf4d215c437df9ae63b59e3d9183432d1bb5f5874f9225a794ce383b491cdabd8103cb9c03bcd1375a70567d878351a8735c4e49b93ec12234def2ca2e1733e5fdd2fb865deb2ebab558e10da58749d586d5b9392be72d17e29a12cb836a5f6867211e386cf345c9a73e57316c6a010c05143f3bc5e96fcb595c5d4b3172fe93a4ab5dc260a3ea7f161e378becc9ac53e86daf4542aee930fd24902308865f66066d330ec99d6b90d8f4582cae38c5865d4d0ffa3b581745a0d9a1d3efc9f8b5cfeb58119af02c37d83136bee3d8b47247aee79f5c174dceeaa51973f640d95b3f3116d43ea481462e620e265282e341b5d035e5439e041f16469977c2f283b801e23f18765e17cb68ce17c62562051ac7a152c74eb51a2670296850b1083c11e4d00d90c89304bcedfbba478b5e7cf6675f3b8b65f58b416f14d367f8946a74e2ba912fd3ff370c2dd7b0193b5db3827a34f109136ecf7d1ac90965a6affdd5674a550e04f49bccf4084f60c9224099fd87d3f610991d631e41cd923a10daf0395ffc456b6b25f79013cdf42844eb949e4ee0f448015a1b5661103266bff980c85b8ed13cf0774c3a62feced5b7c5f6fccb8feae1d4c8a00abb5f4da09f308c0154aa72b5dc639a75cec16d9cefa2f02cd4ce43e32f3ae41a27c1325d95afdfde98ce75a4f9430a0589d9871c75b00f62fd51383a95be02056d9e2fed25711f1aba606a8afbf8f9bbe78d320fd4a73e97a7403b397a20e5b050e2a73fa4039346a4e38bb9d62f65f87d109d81b8e4473c4d71f55d089cf6d8d954fc46b1b856a8cd52521432ce55247db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb1792bd5086499637801499e34e5450c8a029667eadc3a3d8c099062065334023d169e7bbf2668e7b9ca0019c46229655570fd0aa18910ce5907bfa1aa8220c95ae502c80475eb60bf4c61f87ab47702a79488c5c5c46f53099abf09e1b8638a141c7017feda42a87f10b30a294e191a5c59d3554cf1e35f9405c173a3e1661709287425765d87022d0975b81cc2e6177bff696c3801819e593bb9034d9f8f041edb59d089b24e0ba77c9359e6edc26a686e8ad55e097a49db45108c86231b01d8582fe37fcdf3b54f20f676a13affec80e4266424c5344c008c73349b57fd8adf19e9313ad7fbb459e93d19b18b2fff0be5d142074913a90a14f6bcc71db7aef47ce7e6e0ba7b3a9d7f84134308108a661a2c35b193bb50ea1fabb9f64e8c557211597347bbf1bdbe8e1e495b850466a61af5f1893f1cb610062194b224fe3d502b28696ed50e11495daa3328f845a5e92669aadc571f75addc85cabcd92528487bd2bd6102a1499361bc2fa7a49222db7771e53b124e8eeb68eeda28e7904979584eedcf654ae647e813c390333496fbe865e976559b1fc8770e9014bb9d69a6e9324c8051258066a66069b8dcfd2f8f749875525a05bbb31c180218061911cdfcfd9a67757be9799098c52955ae7d32f5cf629f6e711b5161765764094c2be63843578af5b46ec02396195564d8658073a529a8ff965115b730297255bcee0060a8190b41bd8335676c4ae90a243872081172da9b9d51e25d576d3ec155ed0486a0c2ee297d521abdd0b9fba42c928ae707018f96405d9a3dff1078aed5e4bc8003a5270e76b90fad668bc802b1294f70df43ae32acb7043aa9661ddfcd2aba6022fbad7e6ab2959161971a1d80f9cc3a46c8ad4dcbdcd75d452548c6f92104d4d06eb300f318d3471bc3649b4726cdb91453ac93f1b07b0c1e1b5d502b8dd544de300252c44d28171e167d3b230bd1d091487d9c778642f06f67a8ee0124d5cf9a270ded2149b9a325b3315361378fc6bb3082430d13b456ce1dfd772850f01495d62f7c088713f87d864cc10eb936a419e05466ee92da0b8c3975e52b02401a8f18e362f9bf6b3374b3d2c51cf19c310665db9b6b05134cd4d56dd249ea2aa00e60dd063167e2c22759a32dcf36b9af8ebbe91939c87b709a8873675d9d544ad3f3ee9b5a6dada46a349b03acec5da80cf927527a9fb665872eb7463b42fbf96ac54b56d51c4747bd354d8d595dff8faed3ccb871036c4cb4de22ad9c93c4d6e796a93ae38c61726cffa4abdaa80fc7ce473f11abe2345de40136a5faaa6032336f91e9b36215139d369530af96fee1b5f06ecee5e4fa9808808b91c39349abee2ab9423b053794d9734282ebd000fd2334d5579a98a00a9a110e5fb94d69e307a9d80763071568458354455b334ddd69077d55f58b9ee9f0353280b718e2986e507c488e8126dcb8c6682e50e15026d623c9dbf6e2d90a08ebc2efbc682e7d5380063035041428af6a6fc4ee80a9170d6712d05be1730c5b73d15ffa4fa5a1b524e61ca3235fbd9f4b489ab94fefc8bac85401b62fcdc41497dc796a65e07c82243636ac065fcd24b6eef21975ab981eecc6027363fc12babb638b9045f171cb0e6fe790efcb0f82d03776f146458903da83db7ac61595237fa8aea3e5136df194748614edda0c38090ab46844acdf2676bd66c5e6ce55e44bdfbe656668575b49db09e3251794e76e5237ea5034fb2ba5b7c3deaceba9c352173a9ab751dabef096a2b1b1aa9c8256f727872d27140b1dd8552c53420bf39ec64fe8eaaaab8d49928873a8e9bc3f4342bd08114445c59672d522d8ad5cd54031570fbb7a35cd641aa9a37704c0fb10f6d4bb790482e0829b464414a8e42b45a159b6050a3a0cc91b64e25375fee8485c3ec63c16191e427d60c55cd62b1f65e6c43a063f12c230439e5af14930f89f0b57e480af26bdda5c0306cc6e54b1910f24c078ef5ab1a948763e66a902b85e56a4ba82340b7b30ff26bef1041bc6c9df67ab7af53293e5c2eff53fe0a13fa1bd0639d7e2586908082371fb532b9fd735c1087e3a7d6266b97cffa2dd8717415d7ae5f622d55ce908256bea7e49a64004dccd36f44bfea21de3230e20a5d32617f274341f5f8f05d70b3b22381136b5161e54bea051ae08d6de5e4effca7a1fc058bfc7e9f6ad71452778958af3e2e2947b4fd4658957c7a94617e29f910e837023b8cf4b7aed17484d67f8578162479db3d999c4d2dfb16c740a7c1bca33cb7c846ad2867fe1657c95fc3e6ed6512060a62bae49a753acc4100fad45bd9b9335a74091d3095944e64f334b649ece4191fc44cff4a96df7e2d8c1854c0577d143ea216cdfaf31c23fe6c4769178c43586014ad374b44fb9485253d73f384b73def2ee3806acd0a8b3c2fe1b8f53bb3e909e898a5cf36f2702b94ae058103086e8e4cdba54dd67832206c0d62b1c8a24088334c39d3a8ac806df3d8fd39539c8b205a6ea66f8c9404c30a131b7b03216105f08ec61a825f3373f481d41a054aa05b21b7114c16f9d2bea8a925afc18bd0a246595b4c3230866da378f1463158b746ff5294566d10794f4b5c9832121ceb2a4935edcc80103663fae095a325f51a4b3722904423c832f4dc891fc5ac6acce727f6babad551d20746f6de58ec56a3f5d054e2144093d94fa7b67a9030f7e1e5a0357672f7d785020ac90ef14054ab6ed53916519ab88c85e91e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2fbd7eb62824107ba5a0bc2a0b8083731ffc66837fe849cc60bd51a7fafc405c6c5e98b0b1b3aa98dc0a0b409630ac7088d51c191e2db171e8f91875a6968615ec4df573fa51015d57e457a069a6d2c480aed428c6f450f1c9ce27d35e8336ddf59c5b299929308f8520c2ca591d16e56b29a1f4cc3d7f9358ef50116da41f630b647f5d2ccf50bd4b05635524a197b56191cdd82c9dd86558c8c34f06d85bb87908e3f2c1b90570acc719263ab1de835285b4a34c9df11b5a1c0b798f150f4b9cc3c75dfc2cf7e27f9278033796a39bd7b024b09a7ef380546fc5eddb4aa62803a617cb25384586d438b1194b11124d9ddfdaac008f71ce7dbd1919bc0511e7c6cf968498bac29a72d6f0e8b923fab04383412974804a5c6a459a8e1d2c2d918c59d6a2104f6e17bbff029580d4ac5c3f19bf43da8f057043c0805b7972273874dbfc8e13c72d2e52069e3571ab98253e7026fcd52f263f299c8b70a5653d7852b560d4199e3f5ff13dbade385b2f5250239f63b2cdfb1df379462d2b6f7c0efe8bb1a35324514ee8d0e5eb9cf9b87c31707e33883e24f557e0037706185dd2b80130e45b50554c5967fd6cfd8179290be65e4deb1ea0a3005177c8cc0e98469b2d8126d26e21a3593165bdbbe0ab95d07746b4b632fa7b8f914dd4a733094475e3167db6b2a28ec988d21e1a99e5c3b21f82c629765fcb5c49ee4a4d2dbaa3256239705133619862e3eff493c05cdfd06b905ae1b1a6043c97d9b780d8354f1f911bd16d3bd0db57cddca844c447ddc20fd7d994a7981825573c6aabb58a260a4df7727c241215c37a638839d4f7d98e0334ab4e41787220f9f172c91e21906f88166ea0886acbe63aab41385b453d4df4aea4e65da66f16d449c6b336783b73ca75fe4117a5dbc94a0de6843414dd16bc3d92b772cbfd2f1b492ae1505ca94bdf20bbce05928f915accd3a51bce2f1f8bc2259ae66f31224455c22ef7bb46a128b7f70168dfa82be576bbd922279856a22512b1348570ec79c520e81b68348ddf3b1e5d7eb327e3f560229e5444827c4bd2034f7aa17609f62dae2de1fa4cb38280ca75e847f547aeccec50d51ab927e6123cda4c68b064a19589a332fe2ab49333ab3e9e9fe3fa6cc6ea6e3faf88943edd417e407697becd3e160f395ed7dffa466446f371f6f7950bf3d3f675e34b4d0f3dd32cdd55a56069d665cb0e8b6db1c7c34f0f5e1e7879ad76c87a5aa112e75d239f2988d3127457d5dfd1538cd874f0b72a71673304271fc08f8c9da7e94dfb1467025ac69dcf3932ba16499649985ea4064cc19db39fd2f1a3b0ea52e7e19c49b9359fc336fb602e6444b95178d82f4fb57c1ca1a297483218315c8a4c176de924da7ebb192c23e88ccfdb389d104c0e564bbacead5e7ef8c4836574ccdf855fbe458e87ac1d979e477b83059ed50ff737571efe3814ee9c0f887128f1a2ce70af72c46a5e01c56e9327f628de3139cff778406fd745d6b96053a4126fb8dee2f726d2f2ecea306a8f86b95fa64e30c2064f4af4ae33d68f801d330ee5dc9796da9d2f1f686a4e92ecd3408ca04ff980f0b426eea154076744ba3c25d621ca9fb6e7c492a4ddc10f3f7d5182cd6345f6d38d6331092399799f5a35a76583d0955f64e114f7250b33ba32a76a81b0e3f1f85d882fdf7e00290dcb50aa51ad3095a190331dd6126e5b4610c5dd66d77e2141102a345369881ec4c141ce33e224e41a4f88796532989b8d54bfebe66f0150656b1a515c0b9e600c6fdd63bf3d502c0764e058c934f37d8b4736a3f9d725ada75a2d2bda6f177931c1eaf9ee083075ac351b2f0cdc2b826abde7255766385492a4077e14e12ee6781e1d29389671af482910e202dea59ce99445ef0b9b5139197cd8d9f4b38fcdf07916cb4093e8e8e8f2a837ed996511cd0da7434dca25b43884e5073cf88202191de73e3a5b07fa6a5ed584bad4e9f820fa5a117471d5eb4c1e9bd045e9886537a82df22898cd1eafd3effa2d884cfb9d716b760239f95e009a330481e2788538d654e1c7e8cad07f5f3d01c038d56fdabcb28dcade5afa3ed448c2ca5efb9e5327606fc16e9ebba69a4d28f094dd9ddfcd5c85ac935340f5ced0916057ef78bab4a18db671fd38cd2edcb1941790bff5272de72b37630e6715c7e2bb1d01a3a80c987ad0c4abbac842250d94554d784db8f167ff8976686870a36ec331ed74fb3552f80a0279d4def8847df690b879421e7a2cae1ef7285ed83efa1d4c10625246b0c11533dc0fe0441e98111df90ca1d1de53e72c51f222e0bd2cdab593d2786ec9d30d71380b1bb183d499ec13f2ddca81b14d8692bbffec7b36eb3c466fa2e214aada8aa26e5fd084f4f1070b662df1a82d9ed0ed3c3c4b847a90971ea0298eedbde342cefa7037d44d2fb253fdd849bade5a51fa4afb6be88823fcff80edd55ea6c4ba59c8fa153b9539c02b2b61b02dcc7544bbe1cb4bc4d4c501b03e5c735c6de0b34474cb63fc68e4527fb9934925a0b251da8e2d703bdcf4938599b7934d241c647c7f29cb82ba1d80ee01045c23a270b6a8040e31fb56d1d0af650d2cccb8204cdd046e05907e0cfa78fc321cc2bc608341e64fbc00d136e6c30ca413c111bea247d5aeffef800c818dbdcbc6d099c59c4d738530a67a16f54830bd9666cc7e54826992c83c45a311e4bb57b109473b364b912063cbf5a677fddf9f69f861f4843c3de68b1bab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8e65bd73abad534b3ac8c1a3be7dc8460a30940a29b155f2e08679559a61c1974f1b0ec6811382622a3b3919ccb68c950001a61f4954135e2133d2342b59f1c39d1b89bd750ff1cb2a5be87aaa087eda89804da802d13ee7f38b37cc70c7f728d9baa1be43335ad164104d2d8e30fd371ae5b135ea14a261c247c654e998b724e6624095487a42af8823ae2e97035bbbce3affdec982a81463ab7151e931e086284dc7d7b7b0caec1b2122f93f8f3a967bf26e4ef6c2bf1a97d1ac6bc784d0d12ece2a24a261e4a23f5ab1c95a4ca4b033add55430e4a7e970165038f80087473645c0719e121ace9c313049aaf0bb08aab5d20eded0d9f9bf2b9f0a8c7a2bed3f3c578461f9ab8d914df9bd730f1f6c284b9889538882ba00d8fcff3ee86330e0312f2c497be5da45e15470969ef4802408b2d6ab830725934bf189b063581599646dfcf84e45494e1d096a5150f55d3418bd785efaa92c44c33346293109d6d2fa188ed303d36166f87d48ea33951af626149f91300f93ff776c4ab867738029c9db8778ec6e1e587a8e1bded46bc0f29d5cb57ddb8a792371fa271ad4a6b48c3bd4420e210ecdd7058d436a73db17867dadde5528b77281d2096c1fbade28efd97041e108415eb6800be4422212a73eb6abbd26580c0df2ccda22c2959d708059aba879decbeb8325a47704ae1a35ad918b2866563a02546078938cdcbda0ab7ed863060a70f6b845301c23646a9cc9606099a9f23ee92214bc832d571ee886deabd4e2191e11c0814c655fa67bd8783182ca9c22d9838d17dee1469aeedd3b2b118506fd86c6fc1657da072321f37d9b5881960cac8eab0c11bb933acc7d72661c8fa6317e552a58e9a2a03ef20006c72f8ddd5e785c19cce0ab42d3091557695974aca1ec7f87e0d361c86f4ef9074711e158e9cd8bff18543201dd7f14e33ddb1d56ef1009db02d5ba668f0478b8a174ae887f4758eda071db30fec409f32f6c3d835b9cd62742d9a1b0c532ccd1c33c6b38f931864f40eaa44e6e6b7c610c31a2a13193eb9db74dbcf52f6e37b8d20115ba9a24ce76bfa38c7feb55acef653095e42920d2d1411cfb643760e12d1af5acf785e5a786465d343fae3cdd2ec1712c4814c643ae50c3e012de580ab261b4aa0cf7bc546b1542f34ec3c4ad152f65f1b2434b65ba741017dd79f9659dca5c03623d2140112028581d39798534c7a78f65ed8ef58b2dc4262f2aa5fca93ed90e16462f581479b57e1de52a347a0a9341ea6f89ca7a7f03663bebe7b71538ca3e08b071d92c468bb1c73ad1da6baaf0b69df7bd364bd5a277cf64f27d45de7bd7a6cabf8254f82f440ab13d66fa45079778bd6bbb18c346df9d280e3dc19f552d316c36917902a0ea27c4cf0d1f5f1b0a8c591f6a03c8b2a7b74d722876aeda563028fff75dbeb3325f4b9f81dbda5a4372f9bb36043cad3534fa475b7da6c6a65f7d12bea18495dad4ae12d07d6abcd91b69d43b14d5f58eca11c3581adf6649d7aeb2a99794e8d98b359a9d921cb4b1131cf0d21756643d3e14686dc99caf692404ba03488ac0c61201f93eccb45e95c84ad6a69220c2da6edf4011858d1915967c109c7454404c12f62a9158133740afe9705c659dbb1ada937ccbd066c5934b345694d6b1d7a8bbd07a9dff7ddd3288f15e0beb25e98b8e95ea81ad1638918507cec9e3c0b9afc5a0a3f3aa97866fd67d25956f88d41ccf7c16363ba20719958d3a6dbbc1f2d6a8fd01ec982e24a11cfe0a1b8ed2e45895ee88d0ba58f4679055c4942b47cf2ed5a5008e09c5b4f8ddc88a91adaf3beabae75ea8f6101c44c984b30e2e494c1e008429bc0892fb38c78e342755c63b388e667057c8c7fcbcd1a70a35992d7f9874fe2082171370891c7019615a4033182a6051959c8a3c528f71d278fbd2cef656198125a4790c39792915b9a3fe310cdc3ac6d08dcc2b4ed12eb1add584217bce084c19a70a03a5194bdee655a2e4de970ec4d9aa2d996344c66165cc5c72074cbfe4de7b712cdd135757ad7ab088d1d490f26fa5c01f4be229123486dbd88618af6ba16be9316db25cd2a4406c86d93549758b16fea951cc9e2fbac975fc1fcc5310a04aa56e1dfbb8b85a0bb21bb3486e7642e9cb1f3d6f75c7c8d9170bfd7853233a6292f724b01dcc83d833790804aefc8dfc9750cb5536c76d5165c8398df142a7d021356aec2cfc9891c38e28317b1b99e39a8adf5652c49258a6d3962c389ce53b8ddecd7cdda4ad0e7e156c5eb192b808e156348b44cb2f602a5a1d912355dc885e09c4dc432e512e60ea6df92da15ee96981093039cff4ee88801fb094086fd0d4034f6c22472cad93f60d4c36eace87c0a22c39968d361975884a42f96c5be66a658eaf701a119ae22e940c86c8158b86b92aa6affa18c875e3b7200db3ca133d0900b0af19b5885141761021ecb2c3de973e5be05ba5618d521cd6e041d9f2bfab535510320d1ea3203d0f3503f07730feb7b9efa0aaa2baf65ce3ba41d51a79b320923971c6da7c17ea19184679b92fd9ee426c91c729b3a75fe325c2b6804dfe73e7949fe32736e235b187ca6a304ab21d6bcd539b67feaa69165e62295a874aae043e0da18ee4ab8bfe143b1f2a9d88a4227999b0a89623358ffadb3da71f622430ea77294e6c280b8c330dc7f53fb9b42e305d1dd80af638b75ba2e27e246907a623d9d15d42fb26080622a509b185aaede64783;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1a63edecc2e6e0928e447f7a7a0984acbafe298f1228d079b08033c7b500b2e8d2e56e26bc20757d535d19f0f24f7132f972d597b27f469009de1bfa702cd70ee1cbd954c3256219f42f840209b26cd5375a406f0a3cc2b5c40206289da1dcd1b5a2462954e7cea55ff94b6971d5b659b870eaaec8459d203f211ebec6c75b9d3317e7b28000f0a6c49f99f0c070df7688125a2be6718dee4b2fdd81ce4ad98d59f1364b6ae2a7f7126c2ef3e33948e516bdc710ea15fb2622ef01a3494d156bcbcbfad477028e418e32f3519d8df4e6ab66d6bd4669245bea6101416bca37834420d7dfb96d758928593cbed3fa92a328303470b16998367b822df9efa79421d02b099c1d87cda32cee97a9c4811e4dc6ced7bc0b0ebe4008f5c69dbd80f46dd38b7f61c2be1075260782aaa6e58be3050ba2f63e4d04f8beccdcf5925c016ed7bf815e0c0a50e67397e9c1052c637f08f73cea9d4d4c97a26b6c97ab4b39bae1069af8c7c8e368e90f1552a4dfd484c7308e7686c44a98b5c0f9ee721ed0b16d33a0546aebc1d313b7b36b1dd4ef02061f946e6b9595e8ba5696a7e0e6630caa686897257420763cb6c009e47080ae92ae7b0802b96baec2fce6af6f333c681807bbceab143ce3fcbb0716d734b0802c905e09c2fd6bf1b2253919675975bbfe4eeb084688e97c7b66a11864bd54dff6b1c8630aca69dfe5c23fcd97a9c60cd5e0fcfe62971e695f8942bb17a57f6e9f1d7a3146cbf467cfdc2654ec354dfbd04b734f2a813408f82e0f7f48f6a36cf956b1543853a90185d1311ba5657cc5b0e9694e568c0904ca67f8a87af20c5f26d6ea23518b34a0a118b5d1c7b6faa70bf23e23824878d919416cc96bcb5dce0cb706f6fc034f36d2e371c8a1b3a57a46b4649f632dfdec694c566c19a8594801074963e3df51b1f156f4d696635a260bae29f2ef2717aca7abf2c9712fae864003bb7b375670192620d92a655492b08f96f628c225f163c54022d911a716fee23f2ac4b7b14613697659d289a1b16a41095ef1e3c61ae9567319d64338f80db72edc7f24afadc3462ff7b14a5f568a2c04bad20dfe4dd66f8017fcb6497bf08334e3ffe0c7f8b6d639da0c15b5ee82ea784158ad4183eac09bb9c321ac2fe160375412510e187ea1ace58bc6fe47f13a8f1e39d01760b1f5efd91b3d0162155c4182510aa4546e3b16da1c8c6132f13d50abfa64884ccc38c301f6f05237441da54f6885717025b6880192fd44a8180a1a96010161c97f178d303cff617c146f8f5d43f907edc8c954b22399bddebca87454225e889f9766ab857fa3ab8c128562c4d1d03ecdce029524902f461a29de42785907c18c888cf045e9f1a20d8cbd01823c31a95cb0084e206d69b6cdcaf9c66c4758e8667e9d621871b0ea1de5824db82d7b82ea32bd9fd6f316c8905191272ae0638a416edafc4eab1d52bc034c832ddfdce2b2d2f646dd9f5721e124458f66728216131f94caa6b6571c7542b2e54ff60f697dcab47ccf0a121db3bce4c0de062270203ebc890da971f04da32446dbcab8c88a8e9f8700da36025b7de931c7f05fc4dbf9dde8aaa00e9911d7b5478e6f0e93a999c44a52b93c7f76966a47861760121c0f19b5fdbe21f378ed26f4b8dc3ef9fa16d8593a654c9035b2c658ffa891b7941fbf4c7a10a967284e55bd0e46ced05213b0a890e450f72338c4a7222c83c514f6a625769c7e9486821aa5ff0ab6103296e3c1d5165357f6abd3cc5a1340e8414e6a353b4a9d5e468681435f223996f3c8a51684598c0d724860a917b9207bb4d0c93e8b7372c612ce457de29ab90d61044d67f2fc06cd5c4352c309ec806c9994d3cc80a3e909a54cc898118ed1b197b649b3c2a5c0b98da8a1eabbd6a2a7896ce4dc40ed180720e0b937bb55eb6a6e88f5ec4b0b3d5a64c53bfc710fa2d08f03eb957328cc1cdc8614ec4e214c892337cdd4b7be192e1bea58648784f0d1fdddcb129e1fff0a320c0fa4215cb52859c7ed37196d4097c02c82f4d649cfb6d899d31e5f50dc2035ce46b5a506812559c9cf431c3c426c45d44139ae5a558a80360622c74b7b9d014fe82c79f6d10b99da45e912835ac0a1d467e5437a88ab30189146f10d0772fca118404f41572d46659c49fcd9da442b0f3902bd53a1829d12f553a23693846cacd2859714e3a6cdf7d646126890aec4aac8d6ccb7bbc3d31ce5f70b4ecb37ff31aec65a183a20cfd48c2e0e3bdaeb1030a64c4f11babb199f51445e9dedee122a78d9904eb9a027173292002662057bf2181448b3fe97165c921274b5757c5da16a683eb3d50cb10957c7617a828964bf108b4cf4e22a1c760badc231ee65668daf17c3c7ae66d5a84f931de172cc3987b304b3214a46d073826598e86cef7e5243f95f73c483ca01ac009505396bc6b46eb78642282a6a22fbb28a3314eaeef32d72539888f696648e4696e2372f649d6175a0a09190fe303b84b14caf06a39c873560308248ef4683291f9704343db11c10ae1e0f259e38fe870f50e9b217ab98c9cfe05b778035d6d6b055e63b48f3d2645fcfa38f180dfe001116f4ef930ff15732f0cbc5d5c5eb313618315953619f490054aa55f90161daf554353fd1dc169733ce61fe07c5951912ce3a3d40943cab41f31f73d77ead5c2be7250d4cb535787911ba77227f587e30931bed5032c0a1a5ea1d1708e199d382f3d777e345b0c052b540b3a914;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he04d4982bf7fbee12ebf9b1e2aaeca4ed1accfef74b5e6801999946ead4f3fdd4e4b7a030b0d74b31ee43e224723e1732c9ed261dd2579168159c7b4dd646385f09eb66306fa61f8ef7b68ca68a945fba97c3f37823895decd7c6bf6225fa1e04193716ffca3909f06ce7d02844b66bbf674d64ebcf256a7cb36cdbad45add81b5467bf9d0842351af496732e94aa4d8400adfbfa8f8c63e124d81082011b4b145ec413722a3c8f95873ffb8eee8750f8f157c0b3926cc61dc2b3dc6d9fe21ecc41b5658a37a26db9fa78c0c370fa905d7146c1a9062d65dfd85c5d1ed8629945f832466ee5f27afddc8da455502a5453da8debf032ed4d372c6fd287524cad2e1af3deb8df0c6173bd8bdf6701c2002f9d4c32f109d5c0821b5434b4894a91b5583c54b4010e5cb2a231ae9af65753a14d226d6b6fcd50adab785740309dfda46ecf8cc42d6532110ea2dff174ed1701d43eaf090e3d15fad1c95e986565e8a8fddf8c10cedbd1807853314420e811c0d5cf370819d73e1faf7fc63641b79bdc7681b82742996e467f21d400cc908558e67c0df7a4a47a6420598b482805042cd538f9614cd358049c5918410640ed815e44012109860c9d638ee3716e449d6e7f982c403157751f0c7284fb4095c703d785b4157380f12033b6861fd5bef7ed795d4a4c4bfb461f8c67b703cb858d83e0b01dbb2fde252945014268dd7e3f778f2aee738017c050da505a954e67d920b0136938dcf3dbe43f07e799183fe2205a91e8a3d5fcf84e1f7467f3d78b9ccb155e02bb5d4a74ec0bdfabc39eb14f5c745dce9a07526df6a9865006f341449c8510df47d35958354a0499f450d5c361d00304ed71d4306f1f5ce919dae841d20822ac7bb7418ccdcb91cd9ccc856c254a119d3c84e076d5102764dde034a437bf9c6e8d18fa98c4e2e4a85d0ca648637dd49126dd373adf326167feeabc646b9a497f756c6310265d4233b714e591ee78e810a1a770abb4436af33070a302b92e0daa4a713abc42924534591ca81e6078fc6f6c67b9f2910510e9d2ca0d970c874b1350f8c8745cd6c2424962ba1cdc9ad9d485b0bce3fad3f184b322032d1aa05c5e1f4bdbedd7bd69f96e6691d56ebc0ed503b4e7016a0916a0a75c361843a7cfa1360e2c4e69c4bd46d969a2c30930456543d72b74619d071fe63c0adc58cfbea0c7ea40729d9a19886fe684a6a5056ff1c3369ce41f9b00b0067d7524c4b015bb103b9a1c84e0468aa0c39d5302834e852322ad97a45feca88670a79e3344dd88cca85f8bd06cb113e722b5d16cfd36a0c22aad3da641d6208582963d431ca5077508d4896a483f6dd7c68acc83399ec2e0d8f000f4be54c8ca085a97cea641de46d3c95b85a406efcfcdfcc114d2aa8f61915a5660237ff52c17a42598c040cd985eb23b31702e992b1088024ae656f5d5a3971a83f76a86a67c85cc1b4d88023d2466ece79d1196181f4f725940c94a46c20bf87bfacaf7ae8399e32aa077e8afe0a09cb20d46119ebf600c2cea4c09af9b339f70b03e2eaaf9f0650df2373ab8a0bc1b4c1043fccfec7f9f7dc5074b5ce95f2bc97ef92ac511248b5dd4001edeb8fc76563455fead150545651b035dfdbecd8bc8540d3a69256af1d288df22998a34bbe1ee32b572e604a6b65ec380fd4b7a9ea1d101d0dffc8db6cbcf67274fd586e8ce20857c3b4158fef3004e058856ece3f53960afabb12e1b074310d8c84cd3660bc0afb317ff330c9bf841a3f9f0e07547b1a6b12988e4aab2f753f8d1ec4e84225cfa9975c2e910d447367db741280667197544a92702c466a6004870f4a8765863e128841071619c84b472c3f666950648fdb43954bdbfad3f4b6ad323e05f3caaf0770a0965f3f25b3ee0b6744f7d27e8e3909afa39d75e4aa0a14c1c41fabef471f3fb0f129a00a9f6968768378c725f7e3fcb1235dddb6739a2ffd5241a2656b2d5706b575a986968983a71ee8a10a685b643f8ea900ebddfe0a99ec7fdf17108d62829a9ce40354cf1d3263db27947c91d5e49e924fa4a6fbceb805c4040dcf621c7f58629178a4296897fd154e7bb1e2f59347b34047e3a37cd53125e577b9e3fabb453435f5f058349779440af6f4fd778f1be8a09759cd3e42ee14fd38391c5dbbc056af24c71552b57268a1cb16049628b1afbf63d77238be1e94b85e94143267fcb0e7a162e1af98e9dd7c0735431d757d183a23d43305babe25f338dd883927a6cebb3fc509d37e56940230422df0c9508b642cc5e7464d687f9dca546d78c863583f7b7c3445cb64acb0c26876fb46f99909b85fd449b6dbd356deff2b8ebf67c17a23d3389a36e524733a11fe7593a110ed151ca09758545409f789b5d49295389a01e72c256b8275998e56d2525a7ca2de689e6dbfb2c1449131aee2f38fb2dd4bc147e5a168b3526262297639a4d2fbd7e23ad2d6105896766bc1c8d7f897358a3292fb0a22546178a21753320b6a84e6c97346137bfac46f51120b236e11cad7216f6ed448c8fef0a6deebd663dd00950ddaebccceec543bdf65b2282e80df1bf924a77a2e5f538896186639fb5a2f5444cd4678a95c2846454611e62ee79a8263524a94d2485871cdad1b061d2d20bb255fad9b40a19bb6a140ca9879d464f5ad7f0b32a8d1e44c9ee51ea97f1bd6fc8b3374f4f15d51280bc5d3755ba45742d8ccc536f9a3ee2da593c55df640d3efd55df15a74fa6d01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8c3282ec89d32a2a380776d32b0d5751fea2918503c28ca1d3b087ec7e01fc0245c8834978bdd39228d4e3d6614b41187ec3041c4325a569a683a192edf0197c85c38873a02ceacc89f4209348877e206df16ff56e59ac54dbc3d6c29e987bbe334bbd459d482438795481d4ddf853ce70626a4b877bf281892dfe5f02915743ee15b33e8291918b9b906f68863ec3ffa1a36faf45ab4bdcef6f693c854df29021cb28e1d2773241808e19c60a24f33140e64dbe46703220ccfbf6e6f88f94c98b1922ac128b978e0d59a0a762c12395615692bee26816cb651d53ce6e3e3ee958c686508e79f7552eded2a7aefd2abda9dd9ba608794157881539c37a4b5c32c706bd90c1ac891a601b83632ff07f94a53b1e2b8cf2ec5ba21ce7245bdde9783dff4ceac2ec8e516e093648bec62151e03db86f3f40ccd3a67b7c0eeb7ec62e54493a1513ebee6ee8272cd3a955a78aeccd23460851ef531dc8ac60b2d9c6212faba8f1fd113a7d65013f3ae6eabf6a159a918fc90824885933cbd0f846e6e11c3d390b6c16075b0e7fcd68979199926d408339e1aec2bafd472d9acb7c7e40fc208ee7ebd0f5efae4334a0a434288df155ba24b717e945d60c1f7e5b2166418afe2d7e28de8297a72e6b20dbcf8846d8b4dc52ea5c2e4cbb2bac0ffba1c21426d4e2e3a4a6cf35d5ea1c26298e742346c7a8f21ff580e57d549e59ff0f5f2ea6856a2cf20c9052e792e4e4512c9f4215ab196fae31ca1eb55e01084a49bfbdc9a71f4803c32c4fdc1aca57ba57149ff107aa3000fd008d32686ed6410e2a5920dfa651c5b3b08de39ef80665ddc41dc46241ba9ad379168fb1219f6677f4948c434df3464f4f78a0a4e4302ec6d1007cb404b269a11c07b22a071e9c8ecfddcdf7b1d2b048d94ac34d1ae7ce0da4aa92f2b3a954ff507ffe7e9045e0cfb5984adda58fc1a180e99c3f4f629697480adc1ff7600466be21a5edd4f7fbfc3793ed98817a8b7392e12858c744ed89c8ac27c984658299aebc678ee6bc12e6054c439e48c115fab3253c264de8363faee2d8c54a882a83eaad86fd15708d708af8340f2748e0ffcfe345d405eb623c6d4c84a8deab6b5537441412b1572bb76363d46e32dd992d8172eeb0f52e0976a9bad2bf471e462f18442f3ace026bfbabe78db5f9f84ee1abc73b788cd612e2f103ad90a109be491c8fca0dff3df9b1b7ff2cc6c3ea746ac2e4ff6332216833fe358de32401db99ab91f0cb52b578527ed2bdeb356cc317a4addb754a1295f182b705bcb6342b2db4551b3ec994f6dd66ab792bba3805daf81e0003bb8e2c0f850c8e544eb85572c5926dbd47528e32cec7365f432dcc6d025c1d7314ac20c35544e88da2d2e9ff6cb18896209bb40927f8972da326fa0c85362fc28abc6963279b57a81a09ca34ef6a9be6ac5aadcd1204346808a47742ce57d7d6e6cdb894c9cf0ce7a9fdcb75f02c573cd6cd1a2f75b24ba46e6707796132529864fde63ef3d65205ab10ee76a585861bf1d3b7e895dd3f2945f67cc7b80d73f18bc07c912aa37c60ee357146ab84872c13e15b661516a324419c6fadfe73b6d47f64c3a5ea487c90f02c0ced70cc0801c58ca24c9d8a32f1ba5a65eb6760a2fedb9ea7bf48f96f76937f2390e02b8350b950329e7144ca6d5d0389e60dd25021f9fe4441c27bc7b4a58e87e3e094e88caa08977c4bc03f1f178c6fff25894f2de8d63fb93a5e3c2e35034e49b3926845e2c3614deb01cac5ecdbf766f79b31393e906fd019a3ce2902ccd5bd4c27ad596e0e0eeaf5e7c53b1f9c5dc0850522fdfdbdbeff3b09635c5a6a32113371c8b7a09643fe55ca95f8763fa75f737e85d8ed9880302efac4ea1dfc7dc9e76d7c8164928d27c406b17d341c2ef6d7854586cdcc5691119b6fdad8b0584f06b56ab18838b79e6c3785ecddf9ca3b3d80aeef05cddffb389841912abb6895eb1af38eaa047503b4a25a6b2a8157a979d8723478736de7771404a23ae79177dff065e81fbdaf6941c53296578fccac89a3d65b6027dcd3427df2d024a7940359c4c8289cc4ec7bbe8b9d7bbe51a469dd6205917e800df9d1e3d230abfc5336eb30d71fb6cfa3e244559212ccfdd396626ce95b5dd93ca496cd213392927d8fff91a4578b56a2385a819444c1a402ddd106898def51d40a750c48d9e2fa17a41acdfe6ec1201400e4d9d81b29ac1f0f50179eca8832371cfd8d5fdf39d569a97e5ed5a9f9533f6278b2cbee07b36cd1d9fada7be630c76a475f1a266d84649e0d3f1957173ee41ba8a9d79c084b7ef502c57b0b5cab0ce03bfdd0db351880cc88a8d056e51e66bb7680f3c7bdcad24300342a9a7d38ec34c82b6e93ef5e55bc0d3dda96335aebbfbc55b8f0e9a31a6e4bff671ae1c0da44d98991b794f585e7b121f449e9e554d8165b8501448dcba4c91233628d88a0922199eca377191f166d56f5b4e064585279d1f9f267c90f93511aeacdd64f001aa629d5ccef2d80df32b56947168a135b0a773f38253342f347ba4f4ce0a13cb00cdc6ae2f8242bd76a8d3c3f6d8b171f073fe2f130d0571c1540faa70238d2b7555782a59000ccd5e85ef02fde03998eec4a4331d5067edbf1e8bcb7d22e7a107fd6a10d00153e98dfbb2760d4a26fc3ad834dceacd407be75f8cea655b8d9cdf2b7dd505fb37acafde30b1ef1cbebf3d5ca50e684a24e177ffaaaab32fa193e7f8b1392bee3071bbcc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6ba4285cfc28420c3fe574d23b1c029f0fac0d983ed99ee3623cd1f9b2d0febfec70665a7620b4f6f19b6dd8a48714b04940980827893aa293492e28ceff4446f7a25e3de0dd0a566d0689bdd110462bca1fbf6115166177847d58caf5b49223429c93f5752d812480cbebc59bf9bbf6214de8f468bbb7a42d09e912079f71fe2bc832ab45cff702f88e04111ed29f64a28acff6e8d718693981185969b1350dfde6bef76f5c2874f124cdd1b5bd69d7d22c6fdd11837ede07796cad625054686528c6b27ff9c54e3cafa451020e77974ec2e6f35299c87d324956ec4cc0909f882eebe5bfab032721d8e933389ca4b8d5bd8182be5c780a12bd13e225f4a8e4854b375adcf8fc15d443ca9b250e6e0e11a86b74e0719c13bf3347a178a431e323667a8e8d84bd1c199e7036014cd4260b45e9bd2f91cb37b28ac5f7610c96ec4251654d56e5aa4a440bf153a53e130695ab6ea316c9e155b8c189a87198a77cbff72aa15b1100dfdb5034cd90d8ee411f6c94c8486fc433c4ef609ccf0e8fcab312b9e9fa0346710ae147b257409976a42b9aa9620c312dd0b99ab8315e5bd0a6d7ec8784cedf27d417e610ac39c743c90cde2bc0073c9533e4fceee449177e4f06e664560cd2e41ef52c2e0642e1ed5d7aaae28d33408731a42740a5aafb2ba3ace0c1da7e140d64af5384c23d17c06649e8df1071f77df394bcbdb2c2b0c4efc24fb5569bb19918534aa618aa4dde3169c02ff736367c35d3d564f06bbf3b5eb9a6427aa1d6f83d3652a5d087ea10bc3b4012be6640079494fa8f1fa9a04d86ec994da41f5707d6e8bf5b26b7f4bd17c825cc1c6af27d753f18b6eb7b9e975de78721161e62cd467e0dc70846422965b75dbb311a9766e4d555f3c44a0f96faa24ed43735ed32e1dd78b38f2e30980a7689cfd2c554e99de7bef6f653e9aab2a4de60b3eecab39d5802c3593253babd7488615e71e826a07a6c9defc107a24df7a29aba1739702359bfaa7242dd6a75a76908b1cb45d3767fd5159acb7a94ff744ff2eaa0be14937e0de9358ba0340c70a74e3bd632c4bf52ec752d603dacaf9591d94017a98518f6c59f7e6f92f41db4724ea7d529043211fa9218c149cdb29bd870ab52221715f7e8dc6a46e1168760f0c6b37c1387ddc8dab1e85e1fdd841de55e72e598529bee648a4bb17eeb407d6a0b15ae6acd967fee19cd52cb5deddff917dd62a28ce3d1de9d3c91cfde20dabedede2d0db9b0e6590ae3a00f39b0ad75a5100e623f04d69e0221edc41eb126cad02246795239f59fa0c60c1dc17ddb22fac28e0cbae306260e28f499c8ee710a52c9cc1bfd791b95e2f799a76f2195293da6524bdeeaf90ecae271f4f85c0892d6ea7aea2ed0e5274ebbb53e4d90002f8c60df1128f834d8bc9839b88270a27ba2bf627c352050e3811881c84d93cbae910d7f172b5632eb80c81548893b1f30b6a31a9f8284f593b32ff3e012d54a0492e8e3668e6d446986fb9a322fb150eaa90876c1acdca72ebf608fc07eaa3646f7075166c87c19db096ca3340a62f0ade1ad0cb909033f0a64f996793a20e6d0ed4fc917625bf47dc911f368777951bc770347ce5b28faca8080647e3da5d0ac61e2d79458d9c442af048d6548c0c5918fe25980dc077e6aa111439ed6861285e53db8a1ac76e58ebf1f3448d9021caa4c2d9de97b4d7e247e93beb3f50fa03ff530cb6e389005ffee8fe4268d2a887267971c1f2a76142cd9eac68e84927a73025f5706ce5d58adaff2c5b166b63ae9a12591a4da85ffbd6441597961c2ae1c4c749e5fedd37f6058cd6368cc5e544bd0703be54382b44accb695149913747494b7680012c2a5614bd489ae8457a9029d70123ae957c70a065fdbfeef2c199d7599c52ff0e03baf9fd89119b7e99238d00e22ecf455113b18b55b1a92faedbf0a3a95681dfd8cd9109ae581ccad99f4be97679fa386a8d8d9de36f7eb1648de822f72aa8539c6929005736ade04062c4818cc9325361b171edafab40a55a355d556e4c58a0e7b2025e9adf6d046f892390d7c0d60d0ae31192b2a74009dd793081d42c96f20642ad0a179d14205523cd1aa21480879e8d3332f2dc93851f6d068aea979dc8061ba9d84ce53982a3dd64838a903a2e64c8ca0aa49d7dc9a160d4b78f98a73c568bca65c2561f01c2cb8e1ac82e09fc06eb23d9e430b7a80122ca3554e3940ce3d2037a4f96712d4d651c6c1e18d23c445577690764b6c1deafd897a814783028c449121ef4e29895640015227da531ffff2ee72faa1fc5498456a3750e6bbde1325cccc17e0c31a75f65b11e742072b09004f957c785a2f6e201909c5044d6b1a63e8cd69d086440a0d96b8ce672f2300bf5402ad8722a9c12607633f3f8054240dda4ce08e467b9f743848384df07acc9fa2a0e31c4c98aab8a10612d54420aaac41a43e66de8bacb54ede5eff5d198fb4574e4d3461651636f5f079a52b04015578e4a394cc1377fed9a43915d177768718eaff1539ef05b56536e4bf6046c463e662a3f17a6b4a01aa65d8b5902c0c0d82e38723f8afe4d5580bb2f5d6aa2b540bf90a7bc0eb1135a884e5f904038aaa5016d8f2897d57c12c343c072ff8d39bab3c3266280d294a049f3234f60030f99a5446682ae9eef37b573ee759497fcf713da0aeb72a327242b413b4e5a5e59672c1cf9e9fae24ebbf86b1b9a4319de6a68d3c4e79d7ca2a254c5a0f93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h43f2bbba166579ea28ea007f720c52ab22c6630cfb4aee2f4dde686b74fc86f5f0626481d89bafca28db7b0891288ecb8a54282352e93db64afa770490c75e9e0af96e08e0a93dc99e4cd7617faefeefda4beaf89b1c1358d3450db80e4b47355a0ddbdeed61d1ee908b699ff954ca54f3d306961472363052b066a5ce17a15cee3b0995cf7c4cf74e2f936a646562f3753e44717b6637074a81b06c168868e4a8c1cea1337776428aeb0bde112dd740f9d45afc5f42583e76bfe65dbd761b104e513890b30b3ce369141ac99583b0b12ff970fa782fc4d46cc8d88ee131c7bd847f0fe86db70fb5f76ec96b2f9a41ace5aaa0feb23cebeb4017742ad1bde161be975621712c455579d514ebbb240c30fee30d5d2e323db842779bc9846ceafbc932b8e9c29cbc47a75586a208d5b0745fc6043a7e2d61562574567accf1617ee252f7e3600c0413f7dd72d5600ce6efb0e01b52f694626440cf02d4519a0d5be362f659539fb2ab38886f4742b4f8d37ece2bec02197e134a193ae1af5e853badc7376f0e86241a77c50923cfb0744d974ebda6eb30f3e949e4c2fd835912b0d57776e089588483be37a69e4ec2839856b8a46cb8b1a598e27b85b407bb3ab534a2e26e2a8c469bfaf7bfaf0f1b67dd15f38206cf53b0798213eda44ee15a3f59462ba1da582b9237a2bfbe40142f0e07df95417066140718a9a02cecaaf9fa70f1b683cad3562a64b381bf7ecedddc9bfa64f24ecd26161e98eb72632e93166a49837e56e094d4bb0cdb89e77424d92df8a9d54cadd645a46e45a433bce99e017dcd5d3baaf666cc6ba537079496bf296d5bb5baf70df1542b349ec5552236b982d402791c85344acf018de507de6152d9937255a94c9c9df2f9e452d2c05e75cccc1d45768222b6ceb13cda20a19116ef9f63981ca812266ae100cb612450a92cfd273d96a69b7e9e206594c31fdef2a38247b0ed12ce3b56741448ae9b40da58824a472eb35141965f141313563d23071b3f99a492e4c62dd3e05aea0a19a9250d1b38eb8b2a2ebeee4c8272a817bec5d7ca2de1e2b0f9f41cdfc678aef2416311036ab61246ce5b2c09ac77718d67e5185b79652d81d2bf60a94b7524eeeb8a145c21a43f6114e6a23115c8449f283195e35ea04a605a11d4fd618b252cdbca37423ddaa6aedea8abe69b25cfc40e36399f0cf18d75f03dda6a397cc80e67943e7f9c1a9d6936df54f5ca889eadea98ba5fccbf83d92f8d64256282a1a992091e554f5d5153dc85ca19a128f7b30a9c5bb51bd35a4548e19f483edb43cc21015fbbe2d644fc8761200109dcee5c6c99e8838ead0fa5845ae456606ada7abe3d05f00ac9b9b432ca94790631645f1d76619b66f5f3630586193099eab8b29aa4c3ef4bdb79351f4aa87eb0c1c453b6ae2aa27b44c20e2b8056c1cc0e18484593532d3b88f1ec4c5cb31875714663eeacf2eed63937ac1e86f679a93eb8a6d4875aebf2d369b0742efae4516ca4b055d1b951d4f54fae55c8da046c1028b4ba1d9df9e0d5d24bb3c8bf2c79aa24b9edd99140de646e0e903ee7bc453af9aa05cd3cbdff6e00beb1bcf5e426052221b72685d108ddffd6d3c91486e8af24a7d265ba8cc162aafca5e206c85f8874c42d6746e64db4a76374dc03cd62b1d20f008a7dbadfc99a8792bb8d2ba987a3e14f3190d0e12e8a44b4460893b1ef87ba9c190788621f16aade65ecd6e392dbeae6281a70c515b513c99fc53fe31d6cd9ef5320c5337848601066528c5a5715538505b91332839ad7e4fedb7a28c949619e55e4680071609c748d6027850617d0e05725e2a73af6f2ce50b5c6830f51d1da3a5fa504f27d6a96000fabe3b9bfff253e5b76e1d1e314f0c95328ba367dec9908e9ae7154550471c65233cc91b8a491ab5c544bf1ecf653149e98bed52ec397cc03a16d2ce6e15c8280d1f7ce28bbbbfd7188fc9f263eaf3588809ac6117f454a13ee94827be1b30fb72dfee4fde693da16fa7dfb7e0f233e09cd60d0f14f01f5cd09043404920cc65182141b631e40c2b29b6cfef8fb00781742edbdb62a5643895b4a8c26c04f2d759cf71e7ce6187258d88d8ecdd4f930ea9a4fb5bbd2940114c0139b68ad8174152c9d57fafd4bf446b8364011418d9e9bfb9aee1c20b4efb8687d9aa9c1e33fd5af0eea6ded8cf8d7a0404ad1d7d93a16947e3415b912e77ea23b45959b605a019362ebf49814b4c81f215056e890a394351c43419416d7ea3f60512f7b6678e7afa4c8d3201c5949c12f3c05828036e1df936ca9bbf33b331c2dbbd6812b9e1a566606e42932db4d0aac6fb0326ffb8ef6a57b1b0e615f7c792aac25790caa9891ced93a89adaf902dfcfe25987160e29b1afb242e96c51c5fd7bbb3d3f6a94e1c8b6d2ed5496ce1d312772c1d7c7958b3b6da4b4a979187dbcc01a61e9b9ff14bff2f67aad623d6458d9d259b636a5f2db6f48c4310ac4bdf0607e79dc9968d87cb8e3cf1b81fb08426be06dd8b448ed68901c45d4d2b79fe623ede05c96ae709fd6da892a7432f8d0ac3f7dca837ca20b13ea017f0a59f0e037ac3b7eba47976fd5f8fd2d20fd75c6de4cecdb7577870859b8d41ed025347ac1b2debf8a801f3116b696f41c81fcfb5f179b5603199037aa45285c8933e3e4bdc3cff68bd2bc0265488b46a9e8a02e9767b461ce748660bea2286b7450c58a4c9e8c9bb427e2728e692aab36e345565e989e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6bab6d8c5b8f7700c33d61a0dc43992e2b4ea28dfb92d638087f43cca912c894209d1a81e789ddf083c23da15e580ed85cefb094ccfcc0a04f9b5515e24e7b165858e5161b1d7c0d57c61154d1a1012108097826cd4113f50f606924a4e7ee76a2341129fe9ff37aca30338fdeaad3ed338bcaa87d9d86933407b3a6e704758b8220b847685d677e21c8cc77679c4a1b7f81c07476a1b623b12a33e004fec047c3d7bdd862e5520f585be2647fa61acbb155b95218eca4e21d9950a8a0064f32b99085363677ff340d3c5c00e77dd265639bb43740c7f328c9be5d480656fa1e3e8a837e46884c69943f012547636fc56c1fb21f3fd3e844ba0b8d3ac1f8f4bc37d02275485f624cf82ee6e7f2f72f7cbe691970886e0c5736b0a348b5c9c24f3ccc9add62ada939c8f3a9fb0f851431df480566ff782380955c838cf334b72611c144f9f4fd6804c7b0539ca16dfd9adaf9fc54cfdee01bc0caba027962ff496decf785fccc27e89c1322f6415e0e0dc9bb420112415206477755f5860b9b1fe3f016847b3b184862d047959e4b904be84f57aba3234d20379c460c7088a5eac5805cecb3fe70c7a86c9533a9cf1723c7597b2b597c47f6ca9c63161db33351d4c06c8152837fe42fd2b8364d6342e40fbb93f859085f4a25f13999f8d1a94480f135a59e99fae79a601dde0f58b038253ee0c96c420c949b6681f52e11b5b2ed77692d6df1844325bee8917da4d7825d9705fc04a2fca24d1cf04f2b3d751b80b4c758d7a6574bc6a4c7a7c6c756b77a2532906e8b621b81fb27e4c63b1468836d9edd944e4777199e5ab9f2e99316699bee11d66ae3a735976e805e21fa6a381b5c588c7419b3593040f1c7e3b2b8de351ebc4e2713c033ff2685a85c19e8a7b997588ecca6d8a3d17eb45728c66960597fb03f5a640c931faaa6c68803c3e1127a755cf3b0597643cae260a413534711a7085472740d59f820c87927a3f34a95c1341621e8b109c8b1027707a6d1de3bb04337af2dd839e46cb5539d65dc342ab4a8f616ec609a0eb894d781f813d6795fc87be5b6f6c68955b1fd388a70cd191cbfdf2b3ec8493e3193d499bc4d36da465142c04da6edfa9c47f1ed0722cd7797959c838144a54db6e6f2963d79d4d550e8901de654de6e682130e353eff66b46fc222e94f8e0973acbd45b39ce87d476d96c959a93ea24dee7942320b6c3382d7aca51c9f275ae1856f19cf32f2a26b9d2a69468578101bec50509444e4260a55f7d61245b30bd06df8a033559b541804caacb51f859f2f7c0ce6d1719e5bd6a84c5b74b217d7f263e8659953132d7b5e1764ee29431fe0a1cf6384b569f99c196e7ac5f9bbdb49d992ff448050be5494a3cfb1acddc9ab9ff8b74ea1b0efaf260ab80de19144690abc834efd7a6d9d114d49c7ba3681104c6cdfdd91031a4f7d7c5630a7b8184c76fec8f915a474145c6ea7591f9979107a6e884f64b6ef0320dfe3b0d048953df5929eee838e739d3fc401ebf8d7d93af7ae0b48c1c4e37ea5254705e6e0e9962044e4e7fe8e0399966bbb35b92e686969e4500a8259ca2959cba3c7879db49dbefa5ef51cad2a6a09ed5fddb5a7f693dc6fc957e6c67551389868d2998fb1e4ddc18e21366f285177e34621339ffbd80d12cad7ebf8d1c53ef380ba8d3df58c2853395f5d322494ca5911335ec7b3c9cd92e0af5f6dfa5099a06fcb85f66aec528e6e0db35fc0b0eceb40db3524a5ab09074b98bf842cbf3ec716f50086691c471c91083588843ba89f7f05fdb0743f97fc43cfc20881ed6899a29f81a13b804ce180cdf467345c17a34d353f0a9581613701ac12c95a1024ee1969467329a1917d9c9f3018ff1e3c7f9cbddffcca3e8511c034f1ec3d674fa40c979ebe743a7c068eb60a804948f40f27b64c3a8f662394ce335a3b9f51cda65332ff97904ec54c12761fd85b11763223f420e2d30adb46c43e774c31eaed24e366d04a40ec601a6debca28c9682d1fb70f515edcd666496d31d3636a649aa088fdb10d996e920f9d75d3f22b382b1b01de666d76b8e3c97aed16935c61dc36e30310fa12d40df5e6793b167fdc820de8592335bd9448ac73140fe20167888f0e107aebfcd6c5779817b3d53c99f47dce0cf14d076cf4e3d71cd72269c52697e78d350e4c93215895ac62ca880d1f8af903d6fb3795bbd60ecfb13fdabf93ee4ccc5137cf5a8fccef81501286f0328888dbc7fec9c005a3dee01837995a8df0b839bfadef42588f635d29ddcf0d5da6ad15287f7d576866e4091bd9e8c2422083220a22fbdafbdfd8aef37aa0e6b2626c4bd6dccaee1d04cbdaa42a650764c0552e7a7876368efdcce449f5c8d358acc642d103feef4114a5e89655b12fe627dc04b442be9b51aa9f8904030b82febd57c9d4be5cc9d6f3e480e99bf9f1231bcd300e0ec5b6cb35256bd13bffaa5d8b45a3840e9abb95fc8fa6220f14c552967188807bbb94137a2201962313d1d40d7f284b6848bba8504d57f217aed93b1b35ef253ab90b2dc6ead15d649166e491bb5fccddd9a97b3a07709ddab3551659c5c4d4c9280b7c0045e8c59193e8bbb313b668d36c1248e1bda748940c140e5bbb4a22c9895a9225d3ecc9638a3eebd0a12d688aa4a3af7a51e79962efd046485c2d6e7cdede2306b71556b0b84a48b6bfcf4bc3411077cbbe8899774b7b7422fefe49d4c7f2423cf8e84d927abafec900a8e8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd009ab97d42833a31eb7309fdf194532f200468ac05ec7c51dc3fe0629e87a61e9fb0a1a5b64ec645b3f30b918bbd993dcbf5e7c94358abda3ed586489fb32e001649e05be4c49496156e2360254ddd81267e643d28d465f91d296fbf10ae4d02a5cc9a4efb37f0f16d7d230da4bd3b9813d6f84246c2dc49d12808cb0ce07a4e2ecf5beb15da41c5333db8f7e7801c399b7142b7faf3fc40a3936b3755da01d6f71c24ab9aea6f236761aa434b4d72954017a74e1d9c38a550373376349cc3997ed9a83a7ca5bf839a5f8945440f393eaf3fbf078ed5eca434f0d8047060ed9a1cafeb629aa95e1b9581921aa46be38b525e9011fef4edf6b669d60909f2f94dbceddee4b52b72ac6d85e2ccf5d5d869201b16bd4c1b0c55ae1f572ea7d9f3a37fed9ed428864de8bf974528a0e0ecfbfd74c4d72db0e33403dcce9f9f7cda2a5abb43fb930d8bb224b9dbbf4ec32b6278b10a6d36b8a95e6074c1d15a2da283f9bf6180786e852b9fce0d12d2ba18d26739eaa518b8afdb58181c73251c0060923af44a0f7f971b1d37cdecf33c15d313aa5015f090ff72068a55d826e48b93afc80b4eca5c6e474d7a74ec91cc6d673adb2f2d5ee9be738f6d9a38a4b03d874b4d4d44bf7c2f5109f58ce67d0df77f19e169cf34139213a8c6d4b9edbe2241dcf624152c1b2ed6e96b2052553f268c2e43b07941b53d2cb83d32845b349fb489b7b9612dfac862d62c321874f0f124b9ba2be54cd65857288dfb9b644e6af31904fa9599e4553cdc004aa38afce99c77dc6b21697fa99daa0865894967931437669649c7d77d0db017020cd87e364d7b639e8291b63bd14302c86ea674a1bc5fadf8cdc60bea2f8292a8aecc47bf7dbcd1639cae4b203efb875ce54d84c02df7c400852d0035eef79fc4fa140943de2653f8de7da814ccaf4798375005a318f43d5d349290d6812d7858de784fb969cf95584b97b08d35f405016928a8dac2db98b480d4f47575ef1d22b92219e9b696c0be8cd2a4b5ef2b4e389162a806293a40e8d226972d45f56d5db1b2cc347ef3e72bd036ea51b005a3e54a29c690c98a8ef53c932440b8b97d77a5fa29fe1c318129a4ee5522beefaaaf260c1a44183ebbc5b3f6f107769ae2d1f5f0ca668e84999b42a335025f26bccbbdff1d7b458c7f7f094eed31d80017c0f83bfc33643aaa905c6f22b9186e00a644c428391d1f33d912b8380244238f5656771f7f99ec98b4ec743bf2a34520353d6d6950a0bbeeab7f03bdb2fab8600cc2e872f0e3e6680bc8c037c409dc8e125d24aaa54d61f1f034ddc1ed8fe582c2c34a595710979ef5c693c82cba73dcf8237ce0f8a3db0453e74c326804cd2e4b03c6f5bb6e32287ffdb852d6c1eb21474222b67dac3c950df324a25cb1c43c8e8c261de171e5024254023a11c468ae5994560fbad392728d88e4e73590c702b114b401ec77dd5781ae714518106c358a73955cee774f97192022bd907010798d56a191b9d8ac6c7eed3882ccaaf93bdf81dc8026a481cf0f2d831561192986107cb1d48aa8eeb0a9c86227bcf94d4f4b10c4948e9998d2e765a3833d1389720cb429ba93d05a94a6f1200a981892d71b6dcc1b0495c1bee9fff7545abc76e3036f9707306c5dc37a9acc0ad0f19c7a258fe0104152b1205335e091508b290abb3f912e9609c9c3cc3892cef0b0a4a1c8a291d540eaa5c79397689fa3dae45792baf9fcb1ffc8a8ae90f10bf9c62d3f9eed086af26d8f31b7b37454cfe0cfc241be176e703f0d69506df766efee775a9db2e8b24794af59e7ce24009d1f6bb5d23c3cdcea81d0340f6daf1bd89f0126337ad7098bb8ab70a37321b1ed1e810f078e57204d6e087b66301dd6930347aa6492b60f55e558d8cffbd3c9e8dfc2094e33fb6d0e126b0fa63dfec8ec6f2935cf09a0fd5fe3511ec9b8da53e9e4efb0dcb641db9c30d8324bee525709e7a4fb2695443f283a50294ba3309f71d5f48b082edfc9b4bd57a15a324372988b6395d536cc9266fe99e7e864045cbf9a95ed078b4a6688d2f78cb7696f183ef9fc35c08d4b50904f658315831635950ef2638fbe64ed1123230e7630ac56d28699ecbedd4af5001edb9a32496d6584d67b5f3bd4f227fd09d69233d65624d9e5efdf11c906e92b2992947616d5ca0166a1aeb89fce2d93cdacd53da73f83df673e4a5b0947e9fb99db8c60b0541c2dcf758cd9717884c72b6966918c3fc0d40e8edecb9cec94bfdba76fe934a7809ff3bea5ddb8dcf7530a3a916e152f6bf17487370e76393899b963b10a30518c71c217b38c1b6bc2f2dc345fe18829563a019ffddd32035202ab63bfaf0b257706fa4119d6ed135dc0ba25862555500095277a9727daa57c511d051e9722101c6c804547107d1ca14aa3ac15bdd49d0158e0f483a782fde4f70b866b6c0bce8cf36ef56b7d2a882164a57a5026c338980d019ad2c8932cf8dbf55d78bc2175b4d5f75ee3ed3a2f505f0486d7c0d249488436ad288314ad43576dd62e3e4d7b05b8c3693f59d0b72520cbaa10c12cd04b74e4444f377400adbc88e4fabd7f2de29425a43b0d947ee36e6030141e575c25a6804656c9a3a3da5e6c1a818e60158b16fab02292b9693bf98cdc058e2e0aec28b694ca4820d1b35d1bfb1e50b3a1e1f5657c8274d219d6e3acc4370acc6c1afe75e8986601a317bf54a231bcff9463d77287dad371faac3d30b0bf30f72a45a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h915da4b5bb7c43e7298af5aeed187aa020726676c6b7bf5b0260cf1783a9c5c2294218c2c9891fd08a77e3a150900cce0e17e643cab44a16ccc40c8e3d89d3012e4a61fed6876c5ba9546d976f16dc78c0756f882b584e3244d21645ca1e1da3075c71686b7e0aa61953b817cb0e15c6da4295c987c92965b3ab9c24244f1570fc39a04c1f6c851895193dae969664ee114d1b4a99dd53a857c5447226d5e5dea4444a3ee48c74406a449b3101209241cf8ae8a80e2974d22b48814b34ce8f86b7b8859c13a99466d0cc9267071a1cb18682584e5597f67fcd2b1ceb88bc0edba3266ccc3f11862a92b8948fe1b0d821f661fec8d80e5f264a47e9a8e94923ac17cb2c55b8a9364313b9c074b9b1852708d027f4f42e3279d597e1c5d10512cd02c60fb048167344574f5950fd3e60e112b0fadacc6c4eb1b27792c026121e64f69627841caabe3c86e2d562b92c7a718b2e8dd385898990ec40d76721c919666e9a6c637eba5b3fc436c508ac2a6f16f39c26aafe9b04f7b4dcf157eec6c0431227adf39c220a5e581b31a66fccda87da30177c67cc14131ba754af36468a932aa56ba456257512112bea30c687baab390f3a41a9e66de29bae956fecc505b38c6c2ff42fbc9bc519eaa4c50c374d1564951d52d9c33389be498e5bb1faeb03181b348ac505ecaacbcd280ea1fee066467fd3daed48dfc9dd53b637e8bbe7b398f6fa90cc68b0a9c6b19eae074aa3727026319f76d6987f87cf4cd70b3b3b713b996aca04082f6a60b0d4ae65f6ba87e24b8892b5e260157a6009e7268c298d9f89331aa33f2229d85c0e8428bec8729e5379be16d1ab231d049357d3876215536ff3d0205ab3bb4b7531d9355d7c0b00b8f60023e8831cc12e88a9b8f119de0a120d447d68d36cdc01edecf06228a071200e817606b6c6bcd0df13f705a0e4404b5a524e11554cf99a5aef399714c58edddb70c101a8df9bdb5b143fae274b5eddfb10f1ccd19214272b683f7f42c1df0be9b0c50d7b8647230dfd1991fc7c06495b2552d54f6f94262132431f21747ba1c9f7e64d1e15cdef27363868fbc5f7173f768e86cb3ebd22d220d3c1d4d0799d96c30b2c9175cebcc88702b2be4a5e6f49113c44ff99f6ecf5b9633791bc285f5552649b2a404d43827197a73908c342f6fb12fff906dab1b01cd7c088194e87b1aea08fc3a3f33d3da7b6994b01c334c8a1eead5490fc0683a726fac3da183f08a78bb2e3740cbe631135acb7d2297fbc469d42349dfb039a5c609addbdd80bca3e97e2614d063178a2ac38c6d36345f12542843b53839abb5c67bedba165de983033e6f6bfe77449312fcca83a8aeaf2f09d9e6c1d78e32e8fe9d90ff466d44897961bfc9ae846cdc5b75d06b97289741cc7d32d0c4495de931b688d1266405a1c252fd0c085c434d6da4f26d96001e0c349914b3fe2432fd77b3c1a8a469e34fdf890ea53789916c5e968448cafe04d602816c86b67ad359d0c39e83db85655ee0cfc445302b52baf85585ec5c9476990f5a905f211a9fc27a0580d5a9276edac7e4558cbb14f73efac6e4a4aa62c3cedecb07bacae332fafbaff86900ac314e70e4b79e2e5619d1add00c5a6aee132cf4e10848e0fbd182bcb983d14320527a7f998dd42280e85006369b052b74d53660bf812da0f9231d5562a6ef64dc5012e7db6897dafcca52e274da7ca90137cb6b2abe781b097b3821841345d2a5b86e980736aab4c488ca150fa5157e9445d4ebca5c0ee6e2276cb02d71754c8676d1c67d650e9a7946334526dc14a7bccda09d075cbc216d5c12089aade5447d386e1a0730a6b8ea8fafed7edc28cfbf5ff512a548f6542ec9e12eecceb9d5aa3a7ed47a484551e493a5b265b6e0ce64093c3cda09d0cf5812045825500f51f1523d798e60be036a474f4372220f2c034097fe356bb9bedfb357795f6f4276849eb0ed6771b67965d8f811de58e89e50c2d6405885c16996ee30f3657dbfdfd4544b49535e203787acca955b57e5f8ab563713103ee66161d3aba007b5ddf51338e2a7f3d9997f44c1bd56120e04ebde75f3bf8b135006d04f601924d906d55d1593e9b78a5aaf93584dcb5c736db35ef41ff4eba86dd48b61b63fd06c08870d766a2d7316e302aebdddf3999fbba5955a632f8ce3ccc9cc85d85a9c89e48904f8960b428706708ac150f0bbb05dbb33c05b730ac039cf3be1eeb4b7eedd05fca92648abdc37af84ae8c22bb08c56543c67b1abc2f3bebc559ead79d67479ef8d1e9d5dbae293541243b0b0a0cacfcd2e49884462d1b40e269a74f9039295f3a0af951c8447c953eeee69c0e1c8fdf577534ab3213b1d6bfb1a4b9093024ba4be7c94d665c5524abe2c48a232639aabb27dfd1c737d948c64c2350c1281dfd0f1f8c00e70f2ffd6aaf35793f1325f3fd7589bc53a04462c57f242681b38c1bb5be19331f919fe3f22c6d2204a196c396c55340b8bc9f94424b4f5ce1cfd8b07fe872899afe9f22e879ddd444de75af08a4df3ec34375e633ec8dfb3fe540c124936374b89e36f4ef4286ef116c828450852d0ff268719c8e689f1b97ad1cbc27271e3784b4830d419e30ecaeaca9ecc1b0e1739a102d0e326d503ccff0bce58de6b26108a35be0d35b05e7f0e004565c38e922147104789b38ec3c90236fc98f6c3f9f35d4be22d3913855c77fe263fcd12666f1c165685abb0e870acac58c28fbca63b58b1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h92becdbedf6a60080bbeeb9d2a14c1442d95f03ab795f31be1ec4905fe86cdbe19f85cbdb524a6e447bc64c41384cd3f46a800a066819ae06304098e732eb4fb45161dcdb11c0ab9de69fa86922df60fe0fcc5a688d1051f62507b3d5e88db3c3981f4785f9148c5073db5d1b44e999c8b5b25ccd7717f2df031b4ddd187d27cc4b8e154ae39d193c1a9fbd32c5a980069219a65606ef52cd88b976853b5b89d20fd1791214c3d7e79c83835bc3241420d63c81b47b5c578b891270bdf331de15a41ad659005086277b66714817929b2cd064504308f6e9f06fa32e59494d17995090a9facf24b5e1883dfca2b487f896a83a60d444502c8730b158f0afcb104594e56378b5d5f00dce08c161c6cb9a0307b11c5dcfeb7eef63609710ce01e84f55ea13643c23295a36cf654723832f3a20133fb20fef98c35d60b93f51bb7ec555b140716dbecb77ae380e9e8d758f024634c88a68d41f6cb0618133a8bf0c44024d3313b250e02bb4b34a403d9ab06dad73efa53889927f00f7b5e6d3735471329c52fb2d92978f9e5f49aea3fdb64319a0bd040dfc111861aee9a56a624934d5ae8bb564505522db3e2b8796671ac824f3b9c65611841fcb1f28832facb2c4eaf4db5786e04b0b3f16de0b7daf02399b350babd62268041dbdfb109a42da0bf41ca447a0be15dea717d14c916914a6d5f5fc047ed7389e3da5ab4929b8cc8e9a10573c11667bfb7ad3d96d5db49554fe5b9f2b518abf755607b646402a4eccaee16565e4738f1b2c951bd1ec8dbbb8b20540a34bc8d633bbc47b1cd4947cadd127fd15c4392c45b5349aafb9e96c01827188a4e5b1d2cf794e12434f9a29cdf94e6aeace0df87eed282c3ffa2bdad5ced41425ddb32c07a219a8a9224d2694faaa6dd8daa7469a149fc59842f40438c53f9292c32d12186e20fe2c85957245a9c73826cb17da838c68510ff269bfd51b9668007d33bf15ce1a6eda36cef3307fe538f1601303f6ef0c0d28ec05bbe2149a7391d3eb05911d721f12a7bef5d0022d0eb51ae972581bbd204707744d869bd729a0adeafe95d619419d6bcdf2140c415a47e4fbb6ff1c42b1008f6257600dc145f81844343fead3c8d860556d4144e1847dd26238a6c662f320892f6315e5e11be7b8d1f36f7f9899d14c9c9396e2f38c0a67f81f4ac4a83198ded20e406adaff4e4fa1fe33efdeaf6040fa0506f24e8301d1e783adf9d1ed5b084cc3c2fdc5c924d8b83ea500e6f6231f9623e3b4ae28b7703667bbf074b5213023470f686d3c97594833a9dfe68617baff6341c522f485b7dc59386c0bc2e0275793964fe5745e56efff4696204d448b7301fa880f51dd7e47656bdf1ca3b01acb0924d408cf32033a341f6a273e61c1173ac1e194972669a7648738a1643d3ee7f9db2b02d2cb131324c078a18416f535558ff79ba3c0a009419b65b95e2033c7eaee04a5539eb4d2a4e31f4513e4ccbc290eedb4f4c5d0206656f88ee572e4bddd9ab8d4d218215d7789aca639de2d8f6c6149c92e42f4a46dc304a2ee66aac6e021ca6c6d4ba4a9fc3eb0faa6205450dec0683182075bbd8de73750326b1f19974bf29a1e50197a7e45303bb53ed054b29d76ffd16522749d47f8f9b668ca0a0f167a501ba334236f7ec1dfb7e42ab47c2b6bd3d65881a4ef3f1b46ab6c391677df181a328a2f69b8e096e91002f6737b2ec6950bcc127086d10c5532e3aa1cbbafbed770a77f613801a31959af860af7debd33ba4e38bc9f1c7f4e08ede58a017f4c86c6798890b302ee35a2473c2d4d7847a477732c2bea4cd441e3c0846ef7bd9b0153d1ebd53518eb12555f28bc81e29e3858c56f226a79ce77c1dbaacd6c4f66b078b1e3b585699911f7438b22e6389426288ad696d498e0d2aca9c7320874eae0d6e03a3eb49c10b57809f875b2bd05aea4b93364a6e3dd2c0768a72bbce6df7f86187f3e88757eb9c9e48db53824d7a9c4f684d97964151a88c5e4e0bfce19a0546bd4b518c747cb8a5005a4e020588646848d3ff507f262399f61e91fd82f5d310a84aa8961172d736984ff658964baaa477f7b1d7ca12db1f2bdc63499439ed9798753c8bbb1e906845f7bb459c6a35b381a131c2e3cf180f4a0482c19e0bc0cc1abff34f4d2e8ff843869e08a27bc8b111fa194d82adbb0f67429bd2e78837a93ef8e3ad3accaea9e0a17a8e715f168a3c87464dd4e4ec7246e16fd1396fc34f15244c15f57008b31e3f778b9f309d5c18506cb5ac0e2940e6b27aa4304137d1eea90fe755164b3dd83902d4d7abf9bdff45760af34fcafe7b0a588fc6058738590d7e4dfd6fb5f6c7026484f09bf6e2d70e764143e6f40c40527245e8520d07d0197592866ff19871119fef33e8f0fcbc4a1adafe966cc57f5716934bb23cdcafbe7bad35d15be2baaebbe23a62f02a7c6618b9cf03272ba1463e580e700ced8728aaf89ec7f9e4644447cfc9b2a8066bc8c1e2df17bd19fee33b29a9e09f678064930818f0ca5b3c5b042ce0bd139d9ba230951d3709dd5f906af3495ea934f6e9e010be9ea4f98469f168e2c4679c2b6733f1271c8cd80f264d17994647c4a41073b9318c6ba0c961dd4020dfee0a171beade9f7549b25232429c1764f91def8e84a72f61f7df28f6760ad06d5c496985825dfa773b92f3828a17283f383647b3dd11d2da40b184fa8d5cde451efabcaed1f81cf0b34957a8b7ca05cc301ec37e69bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he4ca8ca9a2f759d87ee962daabc374106280d8dab2dd6a36cf158d577a8f4cf4db0ae001438ce4f76b7d3f4a55579d58ac8c61edd9eac35bffc6ab208c49161141b005d948de53840ba940512251fcec2cce197b5bd6bf71d2b2d1a0c67bf783b93df50b41284c963f97a85133858b387c7cb82fa9eb64277e8eb2cf628405c6f43ac37fea50370480362ba198c60627e9b81d13d9fedd6390659f14af1aa5e40cb370c6d29774d9e6f5f808c10d9e9a483ada48d1e8e890470f916c4970a62d677c06713e26c43a2b7bad5b87d59dddc74be487e7b213382ca909e9ccb4be3005f55a484cce791ca8d51667314913e8db7fcc3820460999f6f3d5bafa7adc5ca64f4107a70b2d488addd2dee957f524989d71c811aad77d5469710c547b356dfed68cad181e8ea40d694bab9c971f07afc168f752808c78a83955f715e98d1b0dff5faf8ccce577d61c297cf2ca4cf6d17da65cceec81aa12d1c0cf8539167d25873153562bee3bcb2cb73cfd1ec2dacdf9dda833c8592f835485973cf8c0931a2ea6f16fd796bdb85d5891e4d8e1a2ab431c5ab24050cb99cf3b686dcfe9a8930214aa356cb64fd0a04ec595fab54795f9ca80fec32084b0992a2c4183b2dc1a3c50e420e1270b51fa0b519a6bdf3bacb7b2d063893e078a2b65670ed61d128e9b3ea1e4d7d4f73e83bbe3c8dd0059ccc72b1373c4b150ad61dc028fad3f6823d3dfb97af5173d1f30ccad97d1615b985ead00641034e874e61d817f229de2645250687a1cb22107c54c758160d8fb19832cf8eb156e2db5ac90150308c28526bec441695adc7e545ca033f83d226eeffa58f0ecdd8a6ba8de581474b0c4aebed8144a9574946aabe4d5ebc3466396247376493af2dea77aa9ccaa4eb429514521297bb76d665d678dda713b0e6bd186da24e17b9e1f1761c05668fc8ab97b4e3e4beaaead69e7f33e91fcc423a0db92eb1dc1237350e40ef18ac0e2cacb35d9fa3748d80cb8ce5cf528248ee991e391e330dc96aa58ef56f247c94085cc7854ff45fadadcfc3f98e81723f604b7cc6b134ded84cac3f76c158ca2060c2fcc5c0bc13616ec7d3381b46fd95ee4bd7145bedf1731b5bbb641d985fe93d8707f98b55e091756311d1312a55f656e9848a79996e80a0e013cdc12b0863ce326690821f4b6d9fa1118a2132c994b17f34aaf42b0a70311d3b6a5462f1cdac6ac8fd770a34c64f4cec68f6004d0f64c8c1105c3e4e7c42e04721e8d98546cc0f5b0d52e070ff265db51e21ce3c17b8375043b5eb00275596a381e1ac26bdbef282926aa1e0d51030eb4830fecd84cab31aac73872302c0bdca8a06bddc44cea033cc2aebb1e3089339a85f87e652a8dd23afb6cddbe35a8bbe36fae4ab8cebcb69bdfce612cabca0d7f70fe4c1b488a2b74cda2f1bcae5346e5830a47bf826592beeb5130dfeb39940f126b32addaea46506ebe5134d470c629aaf855b2bc925de7fb13bcd3e487dacfc2aca57df847ad8a26fa9eddfdfecafd883eb151567ba7e4749adfc7a65d5afa140ac61befb554f27818c592bc5e6927a55d285dcf359aeb973a0c353a29bda9aca1f2f2b825e7ff7574980c292f45e905ea7da5ff8e02791bd47e6cace40b2cf6e2c4d952e72787d2782ab5a43eebb38b2467bb672a6571154903ef79ed989c22ea3b45158e8257a444980e3b29e7b7c493184069e0bb905bcf5d4cd167c9440885fb609c715e7073c4984bed032aebca3ac2cd2992ca95c326bfd5c854b39e5ad786a6461bbe91fdc3e0951f5334aa50bc08a3df97634e40753f2f2874cd503e67f4d20688a0f6d4cfd594e5fdb1ff675ec1d8d2e2398feeb9f82b9552c340c4585e54b56d1fefd67833d4ea39c3008528f54f161bed698e61984a2984ef853c34eaac9a17ea9477477c95c30af7b45f4f9241ff4013a446846d0d0493d791d74b787a9d77802bf4db9ff8f0014979df4902cc2ebf9891bed8da50e54645231b009a12815271e48a7a9f85c0e1ccc34d1c8c0d10679926c70fba91584a5dfd0570f84e975c778a0f6ac87b1d5566abba0ee4343b4519f7c48c492393a3598640855978124525bf8b94bf5c428076b9a57a7af2301581dc959e07bbc00e0460562a6c3c0efccd65c1e85aa3c7a20df8fe12796fdff7f041401f2186a81cf1329479ec563c905abb8a489767d32bc8f57bf29462eea77413151931ef9f835495c47cc4fa3ffe5e807c221d1fdb1955baeb070d1b5523d48bbf8098ef67841c9662cbdac768001ad76db2dca1d06b1f7a7f5273440182492ec93f484af026a3b2401054c7134a5f63e5877aaa37c6865795dd810f9f48c05afd6e9f2832610403c85b1e4e5ff2ae7b404115d5ef5c90f154d9fa099f8a859b940e4934de80afe934c7ad1603b86ca6c1a68368ff066abeb22cbfdc62f26cd9deda5cd064e08892f0ca9b86543c6c96e404f4bf9900055c33c0f556099bf8d69299bae037189639c80e65e73ae46ea832d15ccd11411e7d7c274c35e01b5e48f6f35763cee79213ad7ae7d42cb24b6d35bf4515a3962cc239f5fa6db8aaf52027e51ed505c420e05f28d1fd1a689b26b11ae827724f35cc98bd88b973a56a525ad9bc9e58b0602cf7b7f4f7f5ac6283fbbe344b76aaefcfc0a7b090839861a421e8e94ae760ff5b8a622dd1031a8fce68768a8043b3e41ad55c98c9f03cc93e46d6fb44f897d89ccecbdc0fda59acb3347e8b21e9e4c562;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h990a5f464db4844cd042e8d0390fc905e65a3c2bb1ad2ddd2f0d2dc7b5b0439003723fc49ab953d9e6aef792d71da12382ab113481051590e22357ac227dc949f24942e68e42e68c354ca01828e62f8be320c1afa39efc60ed62bf4daa74ec08f66727699a2939862fbf89a729b6cf595d8c1579ed4c7e5b9d5503bbf9abeee60ca8823916151d50cf7448769b2648c8f4b5aa2a7ae6ab6e5ef2bb6b02af3be54f7ea6b000887a85af5c13475c84d020c5376ed87246a278248c6d6f2d0a75ce844ef1ff5503454901ce3ea2bec8f445436d797db9e1d6e5882537ae6f8186657dcacef116a7e68ea6ae1130fb9a38806950cba9a1705e509d5340ad819488be6607a319c1c3f9036d68bd12d34015e54d2243319cd39dfe75cc6d2fc1b89adfc4f91cd04bb6fc14beb116164a9dfe054f497d6b1c82b68a26cc93a3ee7314f74bcd9f3c15528a64363f6fcd5c9e7248541c41cc2b73373542f488d33a0512b195b3e589642e6cb0071970389153bd657829675d05cdddb777601b92d9297c7f2297509b45e1e644342385061ca69c99868ff28578df1c3f9c5590c26c56bcaf7973212f5c9fbcd5d0c817963824e1cdea5cf23806f2b4f95440413e3607bb9675a1a26ca492b9cc1247394a8ad9fa4e114a46e707e91ef1a613e4ea8f8e03b895574057d7dffd04c86816709fc6cee09ae602bc73ba8436193a9dbbac6dfe3353b05e16ac8160dd7d1389efa2ead9e8b93d33b964ac149f4e8ff767043977ac3116771acfee7c69cbec615817ffa1a28a422fa844d818e6783aac78507dbc0781052734247947aa7dfc79d1192adb6d5318243dc98dce04d118e554abf3a0a1a83199e289d180e9408deedc7d66eb3dcfa53d02e62684d4a3cda313f5181509b698fbd03e531a8746bd04cb8408c098b19f7c2c4437a49822401b61a43eabf799a3613689ac7d9e34dad328faaa22e38d018a9f6e5dbd74b87528539835148a7636b8b1b232faae7eefe015489b6bd52dd98209f09adf6780bfc0c86abc83cb6856edb8b543d86630dae83d1ab54843a6dab878be354d10c7f450a7fd5af3380032a4457d30a6f3c25d41ca3e70f95d5a10cbe714baa72f474b20f972b1fd28e5ea3cbf9e3d4424beeae617f3f466515e3a619084d2b30e2e3f1cd158e65d8ea3c3ff03105cf2a830a9668c80cb80bf632daf48d5f9ff7042e11894d7e528701aecd4b962908f424d760a0b2d65f5b8c6226a8deb60a25bd30bb0a9b3daef534d27ed826852dedeab593cecbb5dbf092967692b9a8c7ba4e78c46344a6dfd221caf2ca3a521faa2164324f1f0baaed61160bf48e2d8816c19feb41ed0e8b811b3754def8a0f9f53f132362c5aeb241e6475d32ef3b576db93cbe44d8cb6a9a7fbf93cf91fac5d52d5c875bb79cd3b3d0aec1eb3c25497536aae05c77df8b159eadb913e84674803ada9180a0019f294a29642d0ce4bc214212ee1f5e115f3b30175e00c3592d0edb030345987a93ae02eddbe0e228685d5f9ba4139357a938304ba29c5d010dffca41229c6279279024393d17bfab723561f02da40b7caec2b9410a1ca0e66c358965760a2d217a411b00babfd104fa2a1cf1620c1e4df4b856bb5567c13437386195bb8534b7276da6130b5e67b16bad49ae023bc1c7baac1248738d79ecf63669a556394fed1153ddc9d010edbe3ebc99e1cb7682f34781394ff188cd1f15a78277dd947df3fa5bcd6427943f0933bbe23c8ceb0e35582a60ec968bbe8e414cd899b1b6f5eb9881f736991fa7926f7b1e33306496bf408700a3a64e5555e510f787d4459ccd03d2aa63bf64fca0e137f7b18d56a47b6a279fa8183ec5cccecbd17143c4bd8845789bedbc0a6de3749551b3c0061bc7a77c8ccb7c7e06e3179a48eccf8eeaddc7a72d1981c0875dcaeaf8d2de5ef8f11bdff9e41a122431ffa7ee59def347bf5e04bae28af6ec21fc68ca1d2739c1ae8eac176339da8d7064873b156ddef83faf242a7a9e43f4084c0ebd0907143a5a7ecfa5dd524b25d14add4029398f2167a33540af04d54890c897307fbbd94e608a259a67691afd0bf41f2e75706b92f0516c8d9ecf54b45fd10965da955d0010f74aa6197d878c56b6ede2b81d37b71f437f0fe64584c7ae4d2c8c25b251899534da21128c00af50ab5e5473207af95ac07c6eded4186f1eec07543705bb4cdc17034b761f72064bcf9d5b346af1598ba2a37a41b3f1482cd298d513c5628f0c911f95df63936c35e8126677eed778504ecf72ae1082945d0bc58eb37672cd43322bbe8ad5c2c43620ce8943457e99235ead4704d652bbd7766286ac25c84fc92ef3edf1494b767aedc9d4f3964de7e24084c0518bf1000818a90efa101a5abe696ed900e4fc9002ba55268cb395d68e4c77b12b2966f146f0633191b48237df0ed672ba652d58e691d018d76850ae8c93502bc5ba0033a635f2bdb6176393db3f5fdf815d5127aa693d92aad994aba46919d36a82b0a48d28bb69d423f4944e643a7f73cbc3d1ba464e6a9aec57773d81a8e073b9ed50989855eafdc8d7757b1450fa1f909e4c5770e9518ac1e81e2f6c9de28567349aa894f61c9a5afe9381864a926d42b5af1e4ebd4abf567135b424331a1409427f92bef8db1ca4687cc9b8ecb1dbac7abaeba98fd45a2bd49899e385e6f6d846e3a0b98b2f440d4e9ffd8213d0b8c2f4df62573e15b41e122397f14ed6640995e4769811c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbf9e64359e6777e35c37c87da94589e9649b2267164c880548f1f39e4d76d8648db1e6831ccebf054bcc5f4a958317d7365fa38d1b909a4bda1e5d1cf3619de7e662d31ef87f8d0aad493a8d5ae6a0830d83473d64f55920164abe6d8f99df9659d7a9508973307dc3d82e24398695848db76c26078563b0acad82310e9ba7185dbe3c51d3f60206644b86fbc13c6040f6d0d321c7f02a3064548512eb58837c117c1ab214c7f77d562bbf82b78a6f79ed3b3ecea1822ccd85d01f647441f57457414eb05efe5522df59852b23bb0cc6fe0c00dccdbc82949d71714888e54bd1d7572f94c0aa791ce8173cb1868fc9b6f2169a909de6352bf319eb202ba705f97ebee9ddd56457caa1ecf45291fea9d258d87ec4fb7510714f8bf6f1180d49a5d421ced3767b263b46d56cd10c57f407cacd4e4207834b21ab9766d10dbaebb12dfbe2e8557bc78be3d589ec2951541fcd79f558051494d558337bc2e77bfcbbb46b92df76120d98aace7d0b10f9e70d9bf58d2d2120049fcad982424bd2ffb0a7c49c4cb05cf52c1692b1bfc5321b219dfd2d8488bc84160f1f40317f1c952247b5f7c3739991c21d62da6471fa8eec89c4fa2603c8a67b24057c9ef6e556c1dcf02386b6f2f13f4379576268ed19f46338062492fb2c4279ed6ab1f7a44d945399239db69976f1514e2a71d71063e94a2ba968b8ee1bc715f80a71f732484332b04d5a89da89dc010ddcf65e01fb28acc797fd9f43c77a433553ac8086a50d82f856f38d928a8d309e5a59b2e73ce8bb05285a05155752cd4df1088a71725f9c40d44a6d0c6bb8486abfbe1eeea6d0be302836b392290dbcf188afc8a6056948477422cae3669e656f289dcadabea65c3f3fbf988720467b3823ef2fb1d1e324ac4786f40c5aa45433a86efce35dc535e845e16ef08405158a7149a13f9ac780ba30aa380aaaf2f4e43a6b5df7989e7441b1c421ffd37769f35e11b229e6089dac491e25c684bc56b65586f2918742b6b53ddff20c2f14b70b073ff9de7be87f7b448f4d95f410bea6321794a74c2f2018ea09df2c15df513c537b7d9b0bc82599f6986a331acdb3c796d54370f104524fc74bea6998ff9795711dacd54e6202d132efae96b651f58038ddfbc4f97523d15fef4dcb0dc4916cd56e54baaa32fcedde3a3a6e028b5a917662b1b8fc7f3626f6e1268e13e4e42d8374c2e1e7dc487ed05c846b9d92968b4e261a3f064a42a2f35bc839b51a6a784fd5fc463facbdb6359900fa5e8bad22ca9e2834a4a53ffc4a1e68ce6fb9a85016c9b4e91798a6afd47fb79c8eb35f4c9ebcf64e6544e0f744df0f304df41e0f461ca505990067b677e1957e4cb29c63e717b1bf57d4abbe07cb61f28128faa28a9a6f78a992280c36d1b5a13753895cce5660b65828cfd5e5529ad1e01432cd9220c22abc2f1e07c84ebe1a475ad877eb8b9d1cd702378109f1cbbf501d049e07dd2e90a4b7be2fbff724ca785792ad35fa44d6e0edfa1fee2ce8680bb1df8450043206deccefd7caaf3139b34f694666a670d478589fdce88d65299c7e5445a64f9592223760172eb46b82361efd85ed91c8e062ded524add9ae88f22b3261cfff6a0132adeb01653e27300f4a059fe33cc4e75302a0a90dfca1d0376ba39b30b554a93365cd72b7608f94bb9a6cd49c9ec1acc6d0781459adab7c6d87f231fad1a55e1363d96faf35a3aec5e5c2c3560d100a3f86f076d7cff632bf27d786dbcbfe9d7e827560f5661dee23cbbd4c3f1e68b50f0d8db57e65d1f6896e3596dd22713bcb3e57eefe12b5deb6d27535ea4491b7174fa41dbf0f255e2074fc80f8e93f9fb252f96fbdf80eaf6d58f793d336faa8d6a52304d7aba594e2764a3e09ea3add4b14590ab994cd5f620d36a164974209a6c65eb2fa1978656e3118a97ed4c5b64414da7341d8bf2413ec0e4e9db6d1d1e5fe84cb836aee5761ade17d1ef4e5c48254d3e85ef2f3c9f3cb95065182bbb881d91a006ee39ac5b694e3c4f580582a258b0d3a25563aecf451987a1586477e648539b39b7f26906878a47f5ec4b0c1d2895730f0875af84d77be47bff374398a9caa28b65032361e5a44347f4b3712023478a03cb9035f1ae9c87782edd05a5553f314a0c2e2417d07d04fe881d2349a0782230fcf02cad797fffeed1753f1ad595c781f6fd26d9ee7c61131231a7557448b1d85a9c8b3100a58274d44cf2aff9732ad0a1f9ca7a41896eedcbe9036a8f8e4bde9b199c1c7a1ef879f49b8aad5308bee97867ad1658791574e7d2672370d5f9545c49845afb6be62157803ff2cbbbd69b4bf02894d9373be7d745ed20f82cb9f157b805114fc382a301d6c035b09258aafedcf29d0942586e9a38f8414ba84ec940f0ee295dab6db4ade8e64e7e42f8c672cbab8040e2f92294ab7136927f3f4fcfca60307c2555893476a258eb472757db06a1a4450beb14589796d6dc528d5bd81891ddd7a90bb0c8824f148e4a7b9152b228f7a920fa2d35a1acd1734bb7a65b14f1bc49aa9e57f5360ec21fc12b7f2873660b6690703fc0412e4bf3d644b95de7843623b160af0f1f9ae02f7baeb29887dc444cad499eec808edcef3c5f3d726427d24ed2e136d4d85c32272c272abcc46d3c8d30c30be4ec323fd59bc79822dd020248403152e2311da5b63e572139f65a7ebd5d5e3b73947dd51f9b070c0b05f48788c3dae16c724d5064b6770e266f81b79ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h902915a932770e35cd6bf6f5577945ceeaf1d780aeb88568d382b4e0c3225228e101f5bfa2099680802fb9cce9ff0c6aefae2aab14dffa0e48f6a55f80e3352aa0689645881c5dd183a983389626a795a65443cc7a5aeddb8155a012a7c2e8a546a5918d9a67b4220c0c05f2f67e86054ab85267f05e2f4016df77f12e81f260f86fb9355a3463bbb1717f029565bd9ec6a105e0f24b35cd826cdfeb0fef051efb0059964e23bac8371c5a07c2a2ae5c5f7c8e235e55c17b0789e953fde425630df388b8c23b9c4139c85978e44c8c87d124b1846aee05963339fd76261f41ec06ff977eef531ae3468d39f1828048c29e15ae49d1778aa6cfc288c8618583ee46cfd6a69b2f6e93e1374ef44da628efbab2190fb021583f67bab32ca3984754171c4e3282f40e4deaaf77f5402336012452287df2435d15d5ef0a82be9ad7cb541faf0569c634f3538dec70f67c2dfbdceb6f88e5416eeb8db7b0311c3bd19a66d1fd6fe1cb426f67c0cdfd9b9a0e632859e3362d5b002da0b4f3630512e6f128b20fcdcb91d76a18895286a87a61595a4570c62b5158ab948212541d2063e641d768aafc8449e4b4215bd506456f9fd3224e6cb0c0c12204220970d33c9bb00cf868dcedc492f1b78235c1f9bbddc27dcdafc649b3dcce6557938afc32e05f996a000572a2d238f40121078c789494db6570e2c3051b15d3eae322b9960b2f1fd6b6ec66eb330437569e20348b6579a95c6cec9b6cb9f81d01775c841b1a8044edc6a6f3cf0c190329a5db13fe088f1cda54588b08d5559b23b84dcaa792b78c4078a4f63e641ed21a00f21c2316a79cf5ae5c80f2f143eebc75c20315ffd086ee08033f29769838b1d9a05b1873dc371b6dc7648ddf332b4eac07e678b1b9bccd96e0d72e3723ba4e26556df9e2389ba9513b952d7ab168901c4d535c61ef7c233ced1571d83f14e985319111ee2a48cf196aaa94e6528f1f652b7fb6c5b606562c0dbde5898e6c33fe6ecf1faf388862c63b7bb299e56f1b087d8e5a7b8745c5169a7b888a0ae4826c17d81d9177105abc35bb5b4daf8e1dab98b25c0732c2864c5fc3bbcd53cffbf2cd8775c207db7fdf0eb1393fd770a29241c16b1c981c44a90cbd5f884a28a4bcb7d34fb2cae14ce666b99673a603267d71de15a5dfac48973e29ef77c13b1630e1c32e21152d11f69fb795ea34a8a2f7420faac6e8e3ee6a6b6320b075925d5fbf6675a1a92354d4665ceae80a3f4d4c40c5293b2493912e684a413bdda49e76dee84ba59804a8795b255c7f90a2811ff9337d1c4e9c97e7b51bece090ec539f599dc03a37bea7d8ac826bfdf39ec1b2cef52ebb7ae8f99643c6af8ba3c89a158bec2ac18d80eb41e53c9345bf28992c856f64eb445dd2bfb0468f61de8f4eae8bc53e5a60aaa7546b5b6637287f8e3803ce25a484ac99e4632940dd3e3f6e60385a12ad7f13064ef58d5427629172df3a385dcd1ea8b1bf1b7589155a69c30f2c62a49cda9eb11132336183a21361da6df7f67fd1a620ff6cff063aef971be8e981bc2929aa01cae5c79cd66bcf6083b199f16154b2aa396f72cf9d51a3f5d396fad89b9bf3a59d2d2863376159ba966efbb26e76883345888b4ba1c95472e4e9018bce9b6dd35d52625a41e52f23103b175ee7af263fe57bff872e1044dbffae11dba92f150acdd7a793a26d8b8460a6331b483a854c46abebd616fae6a45db67805dc749fffa25f905952fd517db5d839e7ba7c11dbccd7218c233d2e718a3c38ee830048445a379c5a3ee475a848792e20dff868ff56df5b1cbc8cd92ecad4b3bc7d8b421e1f6bc9b2596efd9312279e67d14a821995ac345e5c165abad78235cbf71716cb86df28539bee5886562cf128c94bcf1a349dddbd4e4df220b0652f92bf90209f3fd32ca75db2eb44b431dff6603dd11b11b40f331ac7b183d978306e61acfdca5b8142fdd3a7a667f8f35a6dd2c0dfcefac3e52507e4d9ee1233e4227d3739956b918b6cdf30312ba13f29922debd5880b17be93236e0a3b2e533eab684e1e67d18365c927f5c5d9e66e9b27e3e14f9dbc9b6e0656372dcceadcbaf81fc41169f3ab77e47c7b38e140459b0b4adf1dc639392520d77c6a5dfb2d54d01d23e1072f63b9af2b7da01f5358f07f1851e681af1389a834c9d3a82fbccc3832aa2603e2a5c82e6b8621639f687f16b15d747bb58fbe1ea8eaa4e1dc5790c96ee6cbbec9f006e1f8bc75fbfe5cb298f0f807296301ec021ce45fdf957f67a8582e7136ab47e96f716dd36b328947ef5ff7e38e4097103703c2b74caa051a5e4cac3c2477df25f1e9b367ef683c52cbb152cb37bad010f7357538da024b17a06c91d6529673e18d8a6ed5b0777258a324a39c34465d5bb3438ecc5d913952fbd164fd477f7409fd072e293a3301205d167a17516b9c798e82cf93bc6a98966fe3de97a897dd6c1c4debda1832e79f20605221a218bc92c71eba0d5b38686a986b3f96b6f0d7b075e9ab573200af5cdcd7969464a34ced57df5d58324983268d18f76240163bd49889f278eed138fddcbab06f9438a216edd0a11afce3474d936d5ccde6280d9e67b2551f6b10d317d5824d8eba8d6de347f2f283bd856afa2f3878a5522aa1b19af1249147e08c9843a1ccd96d6ab475e534dc8a1ba9e27b7ce1f5bca031d28c5f5440134ce2cfc500eb56d82dc0a460a7d735397729337cdcf9c447bc6292554d93c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf7b4ed27decf6b86e16b19d0566bd3eaff398ac0622dc97aba3cab3e47d4ac533633e578fcb80e06243fbef0b8c65e4d83d86d89e01d853fa07934fb97e34042d2565b521bbb2f87afc649050afee79242e101f8a71737a0b10de2363fdfc4e3c59f51fd986bb7a1b550c0be0412d35a7ffabac83bb548f35b6683689f29adcde1cb43829a03bf3755b4220c6d9704664582da147c8d3e8d6589f0a60649217272f51e95c57e521a2d58a9ab49ac0c69ee41c3c3478dce65b468b5059b32f609a76303a143484dcaf639eada7668d6aab0562d684a7d9c0383861fc35a48ee67736498b349deb5df35341110f4aeb8eaecdb19eed58d454cab2373b222ca2c8a7efb71c1ccb07e9c5090daf75682507d4147b2928235559bf9b89349711dcc207eb6416f3224d8b09fec807625f778fab40090f871a6101276437edaeb6a3341471fb211d6298e166b9680690707d3ca6de7169b332baa349ac6f8b38a6846a6665dc0e598402671de42216e116673c857baf8290485f14c6bb0b6d9d882f91b86e42115208a575cf76a3ca5ca680af18813ef9acded95c81316bf0db5bae2c5bbf99daca8816cca14e2a1a2f82b520d086c7020f6cc8907bc2999a2e799cc28577df1f7c4dd286e3180a8df5338fc55178993821e5e9b0d5a3027b52083e52f18e5df1569e33a2d23d15ae3b2411d41e8a865e85ca8c52429bb4b9789f0328d9065dba0a27462939fc77dfc268d303e4e31da51691b42fb27bb82f3a0d7454c61a0565fa394c40b10357cbd9f647eacc761592605b629aba39bb4055d6c94c785532a088867bccf4e69c64eede877d97e1cd117f564965e33049424d6e0dab7c251c5e20d8c12bf30a5840c23befb5a6bfc408ec5e57ab3d92d500f3d5a2fbcf635aaa4cd2bba3959d611effe94ad6fa4bf880f9658bbc6636100058c261b3e1f028aaac523bd83f344cef7fe6810755c714d3f7316642046d11e06145e0759c685b8c3800e10ff7b22611bdf14c26b771ebcf7952b77c527cdec515b1cd15d31c0457a01561ef467e63b6397a278aee217547a00fc3c3b8129ab859193e2295e2e69238b321d2637a29120b4473b27d1f7814f03799a7677707a6369270c071d1b3fa41329f0aafb7be1e7064cec14a2c630ecb46007f6ad6f8f1f50f82ea0c1b10a3abd5dc8122e759f8404c60ccc24d087ecca2dd6fa2a4f70bddd93b932b096a5ee97e407432aca70228111b73161d80a4710b80af6654c6801b9cb0d3294c4f4a0c9328227706fe6483b227348821c035ac440d1f232d802390892b912d5b5096ab7e3ebe487ca1deb4406de789aa5903c568ad885d3173f21c3155cd50991b913423916654c66dedcc29bae70c01c11dd7cf0d8f6c56b0a7955925090bb9b92659375146bfb203b403e69fd0c1e418c681ddec7900ddfbd8aad3506d48015ca387296d5716d0cf95881bd260d5e82b1b9c327caf421c32624ba15ffd9e336bd7c5da252c40506126afa76e8fd9f1b1544b50d1ce143f41c09bc3701a7dab2947d183d5bef2102277f0d163d16c718c608d874125aafc688c8f9e7622a40f6f0e4800b275fee163ad0f5185c2129334de993160a9f7d9809585750a205d438d5b93a60a23e8f0c4c188635287b782a1d1f4a646fb83dc4a2ee6acbe9bafad3a566de0f4ceb13cd9672dcf324b12e7d2dcf1d93d5548a3bda035b6f1f6dfdaa2fdaa56a0d048bf7cfdb0d95b17e21cd25ab4a5d9dc8126a652dfc28ceafac953b94fbc0ac029623ad0930e2f7dc2532cb87e09a053e36669e07176f1494a02ed5a6cf6f4d3f16db6b79e51740d95e66e6538a3bb012181341841c21fe1756d2cc3a1432847bc167672086b47dce1cca79398b73002da7e77caf41269626156137085d93d0cac0a28cca0d30082aea2a70eb2c9813b10dae0a63782e3ecb737bf83a7ca10eee0b80d3a7202136e5cc304054275c14769f47263e03c037571378cb15859710e43f3ab2b49afa8bbcb4fec3d1492f4d1e4a9dcb020b3382f190f53a5ea2702a8aa8173b74bff80af7f139fd199e6f64f5a801b5d088ef760edb0bfc2d45a379d2cfc11c014ba4f237fb785eaff8c19d6734ccebd414921bda3c790de576a2671089e9d324b556f9a20764a132dc7d02274b0f5df91aa5f2dcaba5a3cacf24d3a8f7422b93b9746e5e9e90698188d464498f69a98f733e3af1d982f3efd11c24c8e6733fe2659202d97fb514084f82e59c5d923850000cb394817d58e130423a2cfaf8a0d1cbc506b8942b3ce2bc5092afa539c76c25a8b0667aaa4997577dda2534c03c989bb7db2db55f29a19e5622e493eac634a527e1315dad9f1f1dac206792ad0e916ae30dfe2b3f935ac481eb8b10c31b852e3d3ed978ffc4501787d015c8f4ec83246611031dc0f2dc0167e7fbe9e739a47a953e612432402c29330fdc32e57d3c8765ccee9850db7b43a866f9d2c15a571785f9145357d661c1271a0c0ce707c912f5b0ca5528c1f0d480a5f0b245cf3462108fe1347c291970cd1afdeba1003840a68d75feb1bfbaecd049fb5f8ce57ca5b1cbf91f575e34989c92d5acbd0eb64fe5a4335425cac0e4734ddd668e85d748c90d04ee133bf194f0db34febf77aeb847d96cd13805cd0a465d50df4ab14c70929e947a3f7211fa528dd920c28415fa0b0b0b9b77e24106c12f9f30f76584c2f04b21c50ef6c7b93f16da214d4cabda0d6fff58a2fc33383bad1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he7ecb03ac923b5f39086fe1b3778364a095561ce36adf1c2bd297eb3736994a2b80664de8da22ad5f5025c60a405c27af9dc0bdf4c3fd9d98bbb570ac0c045b94c10702a707c3ac2d5daaaf93e394ed65916c0f2243538f6e16d5e95ca8715f8e9267d1158b2102df336daed8290ce57d644e599cfca4f7531f3e3ce4a975c88995051a5f0856b900b66f1127d15e9551a5176d1a2a5cf23772f88acb162c8dad7a4ba90a4ac4b714c39745330fa0e98d3e1438a30e495313086689518303eb8d7e31ec09de25000417929b848b8d8ddc3d538104404963c8c5fac643205fc4deec3634fff883b22f4e8772583ab4a73c9cb9d8e53fae018d11bb3efcf463f8cddac0da2461091510577ba9978a5a95fcef47c7795d2957b4aee797a9be978aa8f53d827ed11b23a763bcf1cc231bdbe67d0cc52305af562062fdd8a0acbf1d9c38ada7c485a17241784e61f6e5accf4020ab9ad8c2bbc2d99dae38b7cce1b69de89b89bbf7013a299f21611d2278036d9abf5773b16c4e6787828c5a640e47a52027c2c1e7da09683a7bfebc52ed7b0ddacb6e346f776d9e2ee5505c6ea162c69290b42eef155724b83fc7727d62c943df4ee1fbbfb64172831e9fd596709a75e865dc42cd6e34fde1f4bce61ea15e427dddc1245b4d55e986c6c47ebb64c1720df4f2013f908e68e045bb1a66af782137d353c2c895bd13bb7f6666ce525c36747c073894cc4843d386ed052288c7dffff462556d19eea82bc5959db2fde1232b46bbf22bcc79b423083a0362d1ff81b3e8d639261d67411663a890725cda91edad6c95875398ef76fc3705119da25e1286525ce66db21040b2fdd092e9a5ead5c27d93ab86dd86a54a1ba35eb7929b3228503f18fe2b33dcc3ec2f4cefa891e0f1bba183815e0da8bc2993692cfa65aa0f8aa3de3d2e98680daa1ff06e6127fab6e942f6c0af8d11ddb8de19282741a84efec2a5c247c403dd9456a1feff6570bcfc4e4f42c0feeb7164fcf8f4ed8101ec68a537ff37070d0a321ba4aa9757f14b2c77d11a4fa2a4d6f59f0b68a4cc0a6ce58bc0a3e8f286c3d5b848ed1844543edb2b7d35265d586ebdbf237c73ec4d6969344020fa6fed063fa6e6342232e15f1a6bebd9fe54539f239d4b3a10c47d238c1bce6ccc98dd4b027885aa0e7e1dc0f9dea8a64223e70ad77b127ec9efdf88d45e0f8ea033ddefd2eb08ca7de805626c840a6d9c31cfc2e5d874b6745f3397c74bfb9a15103391ef7f046dad95b4b4ac701bbeb17a8add242ed81ab48218887ba58ec50449c06f6d64ae94661b43e274df7e628c2444b52600cecfa3eaa8084c78bcc3f88ab084336c300981180b3f47fd4c36b25b626cba50a933c5c04ab7215dc2ff212381535ee8358ea81643d7951934c55b03be2a3f5e3611c2baaa358e80154754214be1c78ea56a574faa9e9cc059f6bf2ef4b4673e3bb7ff9edd22dbc06b2d4adb03c2f999e589e132a5e1ed95eb4f1d8fc04163fbbf081949e34d98e482232178f75047cdb921d767da7d070326ce67de6b64b43af1672c2cbbbddd71f29389e4f573c45dffca9f1157e6bfc4976fd9fbac1a05f55c11160d83c561b4dce25eadc142020f276900616e94ba244ab3f307609bcae5944b3eaaf2bb9fd7fc269cb1bf7fa1a0f2446a327b56df552d1d8ed1464c49d098610369cb50ebfab2bfe14e6d7d684cd1264ed0481dd88d6777bc65bce98638026897fc7683ffe274d7dbfb9a0714cb30a5fa5c7138e223e519926df34d0c4e4e8f780e7169876b44dea9e894ea7900ac5a3cf1773aa0a3ea2d9878ecaad92838a6ba1674035c174016ac584398e785e43cf3a59be2913ce92082ebda17096d907ab8bf922c73ef61856a9eb81482540cd20e3238f96105e0d50bdc4c53287a055829f0f8d140f74343e94fd4210fac6837355d97fb8ba33d7b41b5832bf0045dbb548629d05ac50fdf29ecfa1c54dc76bedd29edf26dd202b9386b45e2b583313bd630fc499bd41b1a2f2d9af9b45814d4500e61d1e830e180346cd3bebb72ce71ab2e39e6ba0e0e6fde035a2bf2ec361908bac3dfc109db2db23c26222691ce27c8e17f495b6ff4658ecdbd162d79701a66b384c9baad886c2bb9a0c24438156be9d978a76f339fcd7682e5910deec05e6ac0872ebb40e013903babb6e7257a6587f83688ba547e149b68accfdd2b714db44c0684edc2eb0a1aac6b680a4519e055837fe2c198da8d7e67e5747fa7fe8f000583c3107d7650d6838c1ecb6c11c2de1cb1324b6976a76f5eba8e3a5ebd7356c4e9c1f5d8d72e7a2f48e6c6d728d5469bc4b96fc932dd1f24a4c958aac6e9914e8a51bebc1e80adeeca2bf795ccfd55fc3cf4c62c3fca84a0b87ae9c614aa0c72f5c2f7ebed5d0f3a740221c2c427bcb951c2ea0c950b9a3782582e8ba495d2c4ca824a8e0afb62c1b4b37795518646a68273b1b2dbeebaf3bed366343902cb189938146fbd34391172065ada1ece135fdb4b3ae37ad8f68129b3b0f87ac89f7cacd4a89fdb9fe56d96f5abdad1304d59b2dc7aeef4e1810b8b5c2b9c609a8571223c06f3f0f73caae8d5314142ab8e007f7ce29f12dc8f965b08ef379cae27a1bf6718d3bb260972192487d371ea436a2f8462ed2c393c07e8b412cbd36e4c594c9e6823ba678398abf7bafd52908f972374515b542b6297e6d400048ee46429a7d8015d63636b80df40bc9cbf24fd2c0c0cb59d148f2bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1e96989edede1dd40ded2b4830572910454533dbe19c29f430409a1e701127896409d6a9df1cb01e8e10f581cbbcbdde639e3381f7df04c3564297dbf0a18c941aa9d6d850ab1419f323d137e5aeed8b0e2755d10afe4b70f2a0e6c1e65d700273f3d4b054df5101e62403c5a838156d4a7b3454898781769071a1ee92baf363ba4b1f470cf127bc6abc59f48183bbe737aa8b3329c14cfdd7f675419462aef842c1a2f2b09ed5d7d39178086b874b718f14472ce2b35f1d5e05e689f74aaa91d82d42effedbe72ed9157e144fc443f5eedfab60927f3c7760bc37d303a98e210536a22ab14812a46e3b9ff0522b6d37767b40c6582c87becc895d4e690bfcb6d8b0a114e9ea39bcbe6ec094f0fe7d05b7172f6306535555ebc76796d9d3f78c48dd27ea23f3c3c6e8ef3c88a1b531c73f64193ec12ff221806c5814533d699defe0a0af0d889cd58e54be24e164c58ab261de2e286d080810e4b6429454427237026c4623e90bb1998df3f65ec5dde1a5b3f29c089fcbb3d86acd3f2884bdc1539e3d17c8bf7be2fddf19faac20d8d4850b7e8f9dac96ee95c3c9c12dea375d982f437725d9bd277b2c277b6eb120c6acb64c327d3f3c1104007443869a233eb98a9029f97ffffb8b84ba4b2459c80a6ede1ce8c8d2f00119663316db678bb875da66d21aabc7ff7c57fc10cb06abb63d514552b6cd434e6c416007b094c1a6e6051a1ab2e9aa4788f1bcc690297a13c0d431c1500ed3805d3373ce0e038e6f648b805e26e9bf8eb78c2308e02493f92d143ec804d0bb5289302a7ce2acfddb6c452d8f4d2a692b2ccd3176fb98e853b8a5cc977b90cd188ceba7c94b619a335e20e49bcac0cfe043ba4db37bc6f7aea2f8313c12cbfe8b772cefd6aa1f8033dbc851cc81b04014ff8315fa845a2c7873d9d9fc6353fc6424f8e24cca6f025c6c337eb3d3b339b50d78bc3705eb86b44e853878cb91f265ac21ea3ce168f3926ac98f88c60677f58147c7a80417e7c00f402cd2b48b663498e7f674c31c7b604ad10953aac3c8814e329f0312c0d8f1a5afcba2e3f3df58881b704f9f3116eec2e1fd06147e895679c24b2b6c5650982964dcef292985e99bd9c502446b34131ca898709800dbb5584ea241f5d1feddc9ff522305229432ddf479e09dd282b98e0da2437b3240b3bc862dd3140384271731eb584e06a01affcd451e2243ebe3065b5ee476ea37656411fbffb7a27582e66f283ffbc35fd71add541ff09bf538d2d6427dcf92575368338af28d76e6847fcc63ac01c07db118dc4197ad1bc2ce422cfa504e2db95a6e0620318ed1ea565b2488a35caf9b5f89947b0eea11350d5b93be54ee449b03cc6ff1e4833f75c08b16e8726d42472caf04e697d93882a48f7fc9f3cad6e70ee65afa72762f406395b61b0465a00fd87b7ad23c933611662e9c41092a4c947f24e9eab27cc02ccdfaace85e6158820c73ab1557857e1ac0f29d40d69356a368c986014f181e66d4ae04209eb2b0909246f4b2104ad15ca261dae0dfb7507686c3028c9c3f8de089e218167347e951f4459f2f9d062be9e8cdfc33cedfad06aaa895612c9aa3f4f4eea8e2fee9bfd87e48884200bb0be95a90a946cc7eb257c48212df2fb2bbb4f606d253a2f05bfc6b34f5b964eb4ba4abc7256b0d7d7c74469daf7fa504a9369c7203ef3d241449a788755bfac9034762eddce756d5eccae57eda1a4bf5c6c136e909d8847895eee68afae52c2ad220801eec6dd88e255e88010130965fdd63d6c71fb05c52b780aa3e2c0b7774fdf403ab8d925f9d48770faadf140a51c020ea6e32375f26cf4fecf99a9e6f83a7e6a17e5b6af8a5a0862095b296f904b43441f482814f861ec6120ff4e1108e1734104b58c77f18ced144dd4a6404a98ac0f4034a946af41d32a4f023f87099bc9d67e2cc5aa82ab4c4534d0f44007c4423caa8f7ce1fabf67aa12ad6447cc75aad43ffc748272e400ffaf6db5ac81ed08e28fc7b52a7b04ce47680a03ed667ffdc6af054c1532783d8a75b65eaaa61948d50d6dcb4f8a1fcb2d38bebfe27eb9254066e17c7835575c24ea4b922bc63e5d73682a68a0aa909d8cb7819540de73c56a514d9bdf3559a457ba14562ff3f8468cd0c205e479d3bd2d324c7d3e4dc8660f453a0a3f14231867a177d0345ebb295f6d7e081f02a38bcb95bf8e00a3147d209a8c4b3a911608dbc909b336b4dbe9412c0c7ed9231d0ce917fede2d9454961c7c40dd540ed51b59a487563c1177e7eb10c5dcdddf6cebfea4b0283dc050a1992a172d70764182d8cc54899e436bb6da8c2a39e236b46b96564c59b0fca459c9d3d4666c0aeed9424722b66a134dba77302d18499d67c2f1fd69ed13d7b69dc69601d4ea1e87b1b928d1d3e0c72032e1e74244379979d0957456d65fedf8556491b637c2489f51a4583f920bd80a2c138998ec562178cf58fbda59cfd03fad6e2d29a90d272260431994f000fe70d4a0599fe008c81669149a8e1a1455e6eeaf768ee6335f35b272617414a9e9334fabbb0d1c8ef10589493a7b7f86ec677d5bd16a09c3a9a8d5d0f1ccc25e0ed6bdd97779c7972682796dc769c7f677d2c23d5c2bda15a15f3270b676b5d06fc7cc1ab43f45cfb0db103560fac3e6e3b272a4f182eb63e00a208dda302efbf19d7ff6029cbe40309a1fa873e22e6dc8b906e9cb41a54f659395e1c8cc67f6859c0fac3dccc2ab877a93038;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha5f2d80c09fa693610f1bc919a649910889e9e82d198ef2555277aa962e74123048a7e3a995ba9d50d89a682ed9af5edd20b9b267e72b38550631cab7a433f64b65f4decd8b73000e30022521dbf60883e1c2b5a3255ea20e02f139e468d8afb8d4eb13c02f845a2317f3b9b47b6f54c2dea11153d283d356b523a9ac68d35e8bdced31e6c74e2503ee1d6d5af80100b8cd8d8042505a810533abd79788e36c65eaabe620051a9f1556e80643666bff2ae9be129923266e47446dff6149cec1e47303ee8e83d18af1e647386e16e44313ca586e9cc5ece86a0742244d75536dc7b623963fad55a251c16a05494b3e650ab97ac529ed37d4d8bcaab0b1a3099e4d97339de6e5f6e098d6f8f5e9eb459148ed70f53522518433ae6eb458a71360650216aee34e2244f9a61f4c4eecc5f0a56ba71bf7882f2f1607950523deb3982a5bf45ec0a16dd907b6f06dd23b559b2f87d4ce7935e88466b533d188e9d3d391f6b0fe3d39acf19a35937713b659f3a8e648775a4b02ea49a536f8ba65edc502f874248084a9f3f2b4851e762d13864c19603074de9ab15dbfd72c329b7731d6d423117ecc14c9ea4c39430619b96bbe6251ac6ac3c6e164e09653e11a3a9f8735bfe14f0f2cee6de6df422734e72260aa27cdf5504ca9969b43b78da32f7199cde09c506e23e1a20e69932181a762d839f356d678419a7b6a5730ad48066046f3d87d9ec1afe6449445908dce87103e65794f73392bc4c2d8c1a78067bb301c549e0aba934638aaa4e26781c8fe9796d0ecda73a679cd20fe4adb87dd01b245d270aeae7dfea485a817f9af2144dc9ca1f1a617d16280c6de3137c663dc381f2a0c30a9d149a89c69c869c9b57f0a23ab210f789268cd14472a8a8b5879a926bfb9a52ffd407e9af1c05a8a96df99a92a5033040b875f51edc881537bf01c2034a5bbb3417bd9ab648be88b9b2b009ad7d686df0b8e33ef7828df814ee916c1e2ce9114c4d3a03a5407840c09475f41be2d46751404b583188bc4ac406f1bd4ea52373b7c734d407f59cdf7cedc41c04dc5ab76a71a7a5c69d92da544df769a39a793b4294b9afde8d2d58d0ae5645a87d79e12e5d3c3455ba7746737a406ac191a71edb43299907128795669e66c6e30fc1cd28fd0b02671306bc0ecaab82595782103bcd12bbe83566fd415258db27c2f624de6baad72f0d4e93ad67b4020e39f30f69a28d30a220d6b38f8f8fab1207c1c6374f85094e1da93cdd96a084d05716573b56f7449a72769fdab52d369dacffbd06aa3c4c75b68dcc6a20e9c18d5f7c928b9b3b16c27fd47950857ab49f9378e7cf591c1e7f9b8b1a1976b2368e301ede33bd7eff0b9de66f1329007b122551aced126fd59d2b41db03af575746c69c36b48fef2dab14b00eec300e6c4f91793f78b60b5014c990c97f8593a88e617fdadf63ba71b4b894c3d100890d8525fe843756010fbf16fcfbe6312f1073b612fe5e02a5525aae97493ff5f08784b6c038f4a5fefc77ef855d86e8c683d178fcf6460e391af6009197030c3c666a25d8a98cf7b2fae5aa4441d1f2f146cdb5939f91e5e007520608266256e144ce12598e477ad5713fde774fdbaf04dbdcf467f15fb07cb68e5ede39669d3b40dd6f3e91889ac806089ff4521345d7238ac73a83d8ad83c6ab4ebd9d4a7d7343a108ddc4c8d71c4cb2b5d3867f6276d279b184b1014b0775a432ee831486292c71d45373b3cb386b5079f81f9157b44de75d75d89aa3e4737c7afc1f39343874f644c59805f3761d7a774293b462d53823ffbf743d702447c8976ce72c7a0a4433310d46cc7e892f6265ec08be833e7a4f0cc069004df2f48371bf5d2e2f850fe296629c56bec0162454e3130f316bf2dfd2751d8722fb8e3fd61d09a824dc53d39bb71ea983d2ba3e295b4927c09f9e3707fc9ed18306f4a83f0ed2ba0e35e80d5a9f3b96fe9bb0e653819742e991e7c17279b86a8570d7dddb4656aec4381a7c06110a814d975f9bf69c78c307b9c95aefee572801c0b1cc8c3f0ffdfe34d35de9db14ff893678562c69e9ce0bcd65b54318782cff7fe1e63329e4784af3a67df431aff118331fe9514bd8a9c4a9a8abddc632797a5aa50a21ec50ab5c21eab3a45c92f63ceb114535821db852c79dc31b1c77cf32b728d6e0f623e3fa83f409823ca405899a590b1bc04d6a3a9b969cfde9a9a60a3354a5ac569efde6f32efc3fb49038d0542e48840d7e71b241ba30bcd04cdc6a749f4875913c09e101e1dc3a20079c6490af5fa278e6e53190bfdd3590522dd4d203ca056d3b0f0eea1d159630e7695b45c94b843d0f29096b79a0374a358502bd63df2106d1ca2c5a89d5ef1305921a92cebbe85b8a963d56c05ff473e2977b5345dce23d1f5e1157474fd8a982aeec96df351047a0d43b5d8d12f97bb70636b968c480b63de9d00e101aaa56875c90aa90af591c9f9da0ca542316c4fe7ed59d2b29b5a7dcf0df9d0265f5483ca75055179a6c065575a611153e72028149902fcfcf25308947b90d3efb195d65bcb0f924652ccf8ff0986e6d37103252c30596c31d7c03f869e415c40dc70a5ff953bd93de22cc89ff25d1f385349befe898fccb8419902dc202ea5225172e84f5a305b4bc6e447d2fda4e06cbc4bb0b60cccb82c45ea023d33623870a6e204e371ceafd0e27abb0ebd29d259675b82707a1043ee59f3f9a6871c1ffb425853c7b997771;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h23a6b279169b4f8a891fb31dea448075986583b3df060885e8651e8d5c0b4acdddb846b213b92a0a80026a2237c183331f49a175ef74fd19e6eaebcae8cc33ea787184cc6d3d126a6765af3aa52dc33c8388f516bb95a0c34a6107df2971c1ca6037ea20b8d7c93f7f7d974de83c5853959dea6837c40fb2591ff2243af23ee4f263f4e4da38a7e64dd452945a0920420f101223d457dce4b6f1f21378642be3c3bb3099c0ed3954f4954091405694e479e263493c99431ac3bf1c80bf64d2b6d617f7b2750e37d716470833ec8bf61b0b0a03549d324db8f777c976267d081f6ae7f403f97243e03222e4eb6a51a005b045a09bbffc2c59785ceab5ae56c77d9bae2efce9bda7567086b76ed893d233c25abd3c3928fa87fce77ebc3fa3d65a1a001ac86bdc016d4a0c0989ae78ec7dedc062e058be8855fa4a3c39d87a585f330542ec7b9505a32a566698079ab4fb76692f8e77db48e243ecc02e1b2c86be1d1d987caff886a841c99501fac0ed734b85d93126c6b06e3ae980be4aef9669ae9c72cea84cc2baddc46491badc44a91d9d8391576cb209d9ddb7756b28016e06066df1b715f58ae133e3098175e65801920babfbc544e455a6d940b3e012fc498ba298707b4b20e25f39dd0189b07c95a26c4c0ca707b985de5f5f49421e46a6955fe46c50f22830c7386315463c9c945c3f43449ec7d3ca032df8aa33b6910c0fbfb53738acbfac3f398a68c1ad5c3baf5322b8a31ee9ddb5dcd06009be717ebc58f090fed7389ad7321581acde082b5ef86d7658b0c288b30ffabb6e445903fec530f68a251d2a3d57238cdacb36aaef582a1db4c9ecfe7bc834bf70a50c7dff8acef6cef996aeadcc114c55990ec141b53d2d13da13bda0d249534a60645e5ed160712024689ad04e592532756094d663debdd3aaf524ca45d165c08ed76e433c3d1d88870d225f2551845f4a80f81668479d69088fb94907b74610e1ec314df548087afc8e5c622dc60ee0c2d0d280b4510e989fffdcf26f429af30dc274c55796df097b5be27e3a411c1a28c1144b1777fe5139e5957dd1cfbd598b0d74a8dcea9168ad2924e3d7c2fe5971859344833ecb6fc9e703be157b43a0a4b18cb745de22d0a11a69d6ecd9a67d7aedae10a9433ed25cc09ab648c73f9a68d9ba29017746caac6faa0c687a45bd786d351816709a9400e6a39eaea461a1e0d88eacd20ccf695648ce9d1cd597d34522aa5571e10c97a034024db1851ecd35ce4c0a07f7f6591479b4f1a71cc4e7ca4db58011fb0eb3812698578b8c4199bcee85a5412205e1ae818aeedff13943c713314c24d45ab88ba24c366776c695a2e6e1a978b217022da4166fa58722fb8b0fd647334069eda1f8acb6804deebeced45ec355e7cbeac74814d58eba17c71328edfa8f2ad4673c5147a8538d9439e48dad681052d3f030a96faaf2eb03761106d22b81a00317ad5951bd49d9034826c5b87ecfa8b5a517acb693c288a4d9ea6727d4cc60622b3e5344eae72beb796d1ed320ae622e8046977e52f44a5eb7860215a3633b0921efaedab518a81442e7bf9c0f175395a6db1ec9944ced10037bd3811cf9370d71a4e12a6cb29544730f2f75d0fcb29005b225e5ead5908c2ed9858af9a2da1d1144edb5988247d842de2b4827062c96405e2897d445cb92b69f075d4e7046158b931cf2d2e8c49e53d493d21368c6b88a3a5bb624b546e0144bb6bc4b9f0ddaf27d288150ae097bdd8fa916fe1508403933f9747ac09bd92d695ebb4fda43770c1839cf29ff57f3324fb8afcaac62b6c553b03b8ad489ca562616c94b5eeaaccf9c32447267928caf47b86e1894cede76cf3e6ade4781c08a0e723e130db9c59c43e96ec7a1f332a6ba78fac21587a84fb722dc9392aa584363607fe85b696a09432a7115d0d01dbb2c5c19e328cb5804ec22772feca66a29e3a8527c090af6c71d91482ee0d3b567e8962dd638eafdb571f47f5ac93a627e114ae4570f209c11da990e54e596c372489fd5a32d45675d0df47d3ff948a5d875b161676d4f181f8ed07249767ce2de843d55544690f25ab2726e685aa1dda2bb4ec7b07061612b40ee6d443f50bb84fcfc4b905779fbd1734d2198bfb14370bef4eac3de081e8aacbbb8f746d340b47eab9543c3f1a9e0d016f4eb99147a9f6d4fdee55f8ceda2729d569ae60c5ad9bb76f6abd8f4cfdd54b91d6c93a2fe4f99def34b662e09ad71ff8897ae4a87fa7d5e451b4d9a06e32be866e8c0d5c2d4a7cd49f842c854871e433b8d6b7b4601d6a4a17d56cc8f2ca641a655710398e9faaaf4a43c45f364a81fa6a99116a868093cd0a7c26b840d097856b320816e6c1b0071fd9372b5eadeb917c8119873b561689a8e6c9a108bf741a67030a559ccdd5295e902d4e82f85288181c5f57457b9225b87e0d8ff3ce041fe6cf4fb6f489a908eb6d5e958c6f4b1ed81ce75905b3f519943f7c45d158d69d367eb903dc37864bcb3a691befde1b62c3b16ffc0189431de64baf5771e9d9dff5535162ba1bdc90305fb2ce581c2af0081137e75be91e8db479be7b9a2142828554a7e515940eeaf70446b48eeb217e40ab8065bce10ecdd71a0930c29319dcfe2d439b745d4b35f28c27055d6476959975986f898f4315d3690687863e9bfbf7b76f5a48812218e83d3be8cb6de47bbe118d916254ed8bcea199fb7ef01997446b59be561fc08bda120a83dc6a46b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1f63648e4ed88e0cef6f60eb6539b24cca3a85f7655a560eac0fb8c966f1564e837e0d82d4eed9efcdea807d2c1acf6aba3dc313bec46678499d07ff7449d25876678e75419220d8723a31d4b210f907a13c7eeffd93fba655a06f75c96b052c67a1c9bd17e65404b1e962c814264aa2713fd5c3c78c0f33f6543f271a4da2fac8c92f20119535fcab443283c7f91b9e35f6a8b5fd4eb9b36767e43b9ddaae9308dde1d8c05d907f9f6e5475da8b33057b46d849cfb407c00830057e68e7f6e6538a3053d07bb62621c5eae2f57df02e773ee83db1fb7ea2b77f24e3de6da4c8e77fc6658307a9e5a450b4751bb0d80d436a2e4435c661afb03d238dcdddde48f0664b9544acf276cbf6f4023fcdee4f69ea41f0d83b1612a9417efbf6a46d31a93e9c1d6b35457ee345e9ee2fc2ec0ca6b0a13f34b3a810907f98ac0e786a3df80d05f198e4eca2c5a2dff5e679821035897c78c735dbd6e8d6db81bc4c3855ba266cbaba6789b9a24ef4bdbe3a20e44ebf6a50d1f205af995772698e0bc2bbfd310ecd39fcd578b791d9d6bf6f118776cca800adc1abc6f19a034a7bcf2ab471c2d61d8d22113d238d6143fcc66505d43d21986c11aba2caf2af20086c0a242c897593480a8db59827a5d566e80a3e841c4868b93030f39e4186662c6c9e95789abf209125df5468ab939899f8ed318f2b50e02625dde8d3ae59f5681aa513ad8469b2e4ee3c9983dd03cf31287dd4a761e35e79137704a91d4473d80f1706fa42933745feb4314a0057bce137833724f5ed078cac9e3bc6c46644044820ad2e30ce1bfe8f0d7c7c09cae57c908af0b770a92aca486cbdcb3cea3424de75df4b4c7e5e600cdaf842c8b6746566f593631be31ca6331c45bfce792511725b8f1f714a2a3074aa1855650b05e306d3829fc175914d536c4d7e1d74d1d869855b3f10c704668f8aa0ddd06cc8a163680bc666deab8134ec9543753ee0ddba9f9dc826acd3f2ab95d6b9b05f28c74c540f6af45fce707f14e27e930138ee2c6696f215c282e78addaea495255c66f5fca2513dd287e0d039aa16578263d819c7fcef8f0dab21b7dd920b01d38fa01011880715ad97cb0397006147c464f5dbdfbbe63b162442da909fa16846a5af568ca7aafc84d81c68b9ac28cf3dbdb8f6015bc02132a0f7abaa5f38f8f8009678dbbeb0606a791d5124c15ab77fc1598ace9f66dcd37489e22c2192a24112fabfcd93a5b57a19959afcb7c4483ab105cb6a53d5208cf4e3321d07fae2bb7787aab0d817389c4462d766860efe97a85c0efdaf85e85481d66250e2badfa9c6d8e27d878732c070ee3535e5f16fb831bff98674bb3e83900646215dd7d338a628a124d2adf76ee04a6c9e8c0ea19e625826bfc6f2253a682a829db29debadb481794f21e7b97d81445acccb1d78ad0c9172821f88ea60770f26ea69d9a367a0a93b4aa3833f1ab07f7425206af6f06848448dc344733d5cff98d920fede751bdd2b04e29297e4d2da72df54f775a7ae6f81defd589284c602d29c35f38993cc9292492a82ae96c9fde5531682e5db6f7cf5adef823005dbac5086af63e0e5760b4027fd56db4f9a865317bd54e7a3d854a69c5cf5cf58477fe4b8406ae505d88a9caeb91e6165280d5060c6301eeabb9d7e76e02e813484a8af51461fdfa600f3ff35dd7595f837506456e00e7370e8f3f8e1401cef0886daf4608bf39490cb387fa4d06569f75d3cd0c6a836b2a893c6d68b09b1b38e6ae5915cf44b77027a50a4e5bb4e1b27d977e210d9b2712857cda376de5012ed19a38fd41263e65d853de7e4331697e566bfc0b99642ab3c7a1a9eab23934cc89e1595010d1118328807b5d9dea4ff5cfbf35cd10b2aa1dd8075b86fe9a7d809466c1e0907da20cdfe3642bd9edb988ccb6a3c5926bbec5b2f68e59561822f347fceee49e4e8262f93937edd9bef747664af5aee61a5f2347da0717a63c7ee197818325ea8f78aae4a7ad89945820a73943588d3a8d520da55016ea6e0320897062488139341428f5926673969658989927d1dc811181cec090cd34d01f195f641d25d874eb2b050f5f68a3ab63d485232820b812c4a91217c958dfe87d8ef95690ee8033cd3db2117e15e42eef2b0df7588c27f30d82216bd1fb8bb8e3dbd23ee802f4bd4b47aeb8eaea647eac96cdd03c76962e6eb9544feade715bd7fdd0b1daa3776cb8462966bbb56589a92e204ef31bb19395604444f9be8153d85ac358f437dcc9b0cfcedae887b71eed5341f8a43d1999d6ed192c748cbb3c186a65a17af5111305ee80109c58473ec187dc2ced66066b9e339615a18fb31a55dab2af58b55c95322a291c29490bdb81fa05b075006b4f2355e92ca47a2acc6c88f0f06795a987c782d0e4844212f8de23f81bd311e825aad76733ebb81fc812e06b87428ee598c40b6ba4b91589f63b1ae26c842ec6d77d9ef1dd201f7feb0fa1788809afe8d80d65ccb836fc74554be5545939067e6cf23b9a1797edca9641d9f72c3206c3fa8cb848345718b70b6ec58b3c244f3ac577ed974be282bb7aac72481df73f953087ea44dc935a3262d74fbcbfbbdd92dd7e23b9e97e924c393ddddac3f4a4e32fe88f3dbc8946bf0a09ba8afefbf43403191053bfc63a938b235df1da75ed6c1949bb6631c18456561223694e74dda345ad67b9138799fdb3f1b439430fcd614a7dfe76b2f62e02800bd24700a1bfba06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h10dcc71299ce37f7c7cee08b44215bb48cf948a6fd607e2a4b42dfc1f7abbd9a80159fb571196e38d5238e5a2804a3b68ba692a6e3a773a60527a1615d9b8641117e998f67db2db4e9561f73997474272b0fda477862be77a2e6e5876d26dbdae1d9bbe720becbcda2bbc9c31a293db6d77c3036ba67d15905bea32cc464c73afadea8e6dbf81c11aec232d569c1810fe0eca1aca250ecabf6bb6a41d48e1ce53fb636b279fadb3fb267bd151bd04421b3fd9ed4aa3a44cdeea48c9f71e426b4e9c8796209840b527e33df3dac98635e7d6040caf3f59d3e48520efbff0ffb66245756547921580c7a75cf8655011392a888b7930944f18e153db17b1a90a51bb94daf554a37d4d48d43c2ce0409353f2de3c9775bd6c68ae39a3a20c92d86f4b447f54a281673da30a051b15809fcddde4e568ccd1fcc8b56ca17a2f6334205913222eb20043828b044ac899723f6fd7d68842030d728807c1132c0ea9813a8c6b936f9a71f665d10b88bf91bfb1970f109a00d6ce93622c044d2ca008dd81d6082298f4064ee3cecea2728ba37a30f58e5116146e59e285edaac97dac0d3f06679a2d0f964543b81a5ee471ef9dd6e9db9cb3f7c27ce66aa27ad05a37348b6502281fe5d304f68adf8d138a750dd6aefc763c9b4ee7093c2cb291df15e6e9109722836837b12caa21e1346fd1e9e369dfba99a6a37b9131707d1ae6bd95e795c854c4cf9935ca1b72eb9e49f1f31f7eed2067cd9722c72b6d820761edb4d8d6cdeddf7171e56ae694ed6fcca47ea829c915a9511c8240ad806756dbb301d38ae5e83cd8267ee4c5cd5f108c661c447cbad0a9d4a355f664d98793a8abd311571a91c9c2200908c9ec7e78a093942d9e8325e5346b80d747f50f9d74b03ff3cc460aaa311722fdb7dfe85fdb4bfb4e176b99b26028c21e20c5a280395673faffeccf7c6d17daea3f33833c5b33be9bcff44cfcdf2bfd6aa8d78ab37e45ef4e83f3b7f8e6270569a389706d1a250e78f9e375feff1b5845ca94d406674b9c80de306330b11eb7f8f46b6b4b8b3cdd0b1a0641a5117f990e50dd2b520b080dfea457b5e945b85f0bb5bfbc2e3c08e3f9ebb352dba5c7452115797fa614e8841b2f391cd94f2852e498c0652f6a0d8636db68cd3e8a8484c5f545cad3bfa22bdd6d712082637814e5c530493901a26f02d2b09ef6fdaaf7273d504a55f260bf019be0cd9b716237c4b55fd7d24e9de9cefd298ef921d074d862ec84d638cbd042a270b98b3177ce5c702a3bf0e49e529f89ecb0d557d552f8d384879fcfa16c4fc0506aad248a4430e87fdcc420365c24c7251bd7504acb916036887caed51ebb547a774d7fb3af6a888fc397f282edabf732dae17d0fc886617638c8d0f1a47dc5c49b69aa931e684770818efdacd348d62ad72796b3e4f593a1e25e1f5c17f8a6dbef45e88cca92392970555aa1f0d9057f2078bf4d73f04d1cc510799b4570abbe84be3d350d88ad8a8cb6b47db8a5638aa95e05aba98e11bcf02481e6d3c5ba2f576301b7a755c7e96d6894ae75f10360e93db1c64620bb1b63234f65091308bed297496a5acb9ba25932ad58587db2176463f0a289c1b1437f8137b8b2f713411f8f5cada3deae01545acd235933fdad4f9249f1c57a715a366e7a1e2edcdfcffe2757ce820405798e2eb581b0d81a1caa49994000ca1ccffb3d81191b7815fe15f68ec6d7089fc2b80cdf005ebf057ea24e1c79241d8c685a0847f1d90afdc7c92247ffa85aeafea772d016b95490583c2d46de29b811932278be5b9c0a42a87cc8855937f5f6eb0590e91c5e8f81902dc8e56ce19132b8140b6fd0085d5dd75293f9b352f06ae36f0c878a098058fd8acdb5ca19b6549c0015ef1c78f054871621a507227370080a14d47f76cf5b3720c00b386a7f11a962ca0c28464735dc3cb76eb3e2c3b23c91b4fc909887322ee27628f56559ab3be5719d6a6d81765a287a8a77c96ef3233f4f43e822fe60c4ca7e0ec9075def31829eb1c987464ef8342c92398e83539b3623f9ac6f22fadaf45af5984a137cb7080eaf07d799dcfce1b684eac3e59a856c33713d006c463fe84ceebe1646040ea2905c44ba1356245804bcee427d2dde705481f6350c79133abbdcee273b1b0e05dc638115b8edace9535e127c8f60e91bb5c2960e49ae065d88cc1657e14467b81d0a28dfb0829c42ee7f3f4e1b39da16afad0684d9b9d606bd5505b4db510eed656ca6260bd507766142f84e728bc8fcc804ba330f1dddd0754e214c07477ce506d45eb02b333fe8227a657c886209528a265aadd28ce3ba1154566b7a7fa1a0fd78f5e7cd0a7d93897d7d312cf53cfe71c2a7fc07eec7a78e7565a433df949cfeea7a5983005fba05c6a0eb13e021a0c4be4d73b8028d7ac4dc03a05e2d8f5e1af44978b7615784ec71e2ca549c2d09cd0967dc6537b6d79f5fb5e2023d3a783ce278c4ce354346e71399778931a46d310452e6572998568aee427594f42e28e962e23312d6c2fb3732dcf469af5545da596859c0c801ac40b530210d7621769439703e529c09897047382a65e4387af60cde81c383111dfbd795ce8013ce5abd451735b9f1dd8e2c674beb3a80d2d1dbc185ae83b17724af746079fee04e9b1d2f7b2ec27751918be62e575607ca32018c5b180c9a3385b517d8e2973088ccb36b57329b4396caedd9ee72626839aeba35aae8ff4b3aba35177694251;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hfec81eeb66972314cb5e324f1ca35ef260b46e2886ff28b30d093df83f9554036c2792831619c59ae48e490e92c987d1da8ae87adbc6bcf5925d16d285f4c9428206e8c8e66f17c09bd7b910304f2dfb53e0b216919517009d6008118c7a4677883f8f107ec4157617d545cb112dfd951e32ef89d3f56a87d4589c896b01a692a11ac9125169d54e1ddf95a7667126ab2891e88dc9b614f3b136776f752552766874524845c038923c6e716eac6dd00bbc98fb8493bcc2ddfb56acc0faa7581a39c798921ce5b7de73cca4cd11cc7655fc222a15fe7bb1a78684e5f006d065d8864b1e1de979f6970cacf95b0a65e9fd77af83492742f7aec930969951df595382c92b7a5f6bffc3d73dcca4f5412f58c9501f27c943c82d758c38e29204287337c2c2a1d4b43abb0a54c246f2df4d3a8793ba27cf0377396164682769cc3fc873539316c09a29b0bb61d3ec37d2fc9e3a59f266cea110a56967a74ff4040a1df677d85678796615d460378d5cd00785df9645b05a3a3c42c11ff1301e4eb812c9f412a3e55d99f7739adac3c397fe4770fd82da5662b8118ad2a3c093d344b9a832eab3bd5ac5eb3c92d5acdac91b4c9d1ccc9ae0b6cda2c1c249b32fdb29ba2dde55a83749a11e354d9ced8599f9e2771af56e426a60212485a4a8e1fb9ca5244902abe77561562ab193829df1e09631b11143f4535567b1bd40d412f585043dd331fdf670aea637d005e6234734acdcabaaae01eac6aac225361d7d42417b8cc4875ba5621f5044f4da2569d357b4d4ab0080fb835ffdb47e1336178a27907e82dab199b3a23497f0791056d834561b006f444d38987804da686d98a7fd7229d8f50d36b74bdf06bb4bfb6d64382b78bd4137c872844d03742ac62f8716c779f98db3782661ee3e37eea848ec78910b03aeda03899d39935e131ea5a1e2b7e24a23dc4223f420d05c54a683a669d8ac80e29b89214d7f36bd875184d4024675268e8ff9a4b384c7083c35d3ca7b5ca25737e46d31b8860d87218b4d280004e55a274588ae446f90a8aac23907c9d7b46c4ed72c6d014eecb114aa35d229f9f32a665bf8e988e4385db21e77a8b9fac71ddd645a778b4edb7301c350a85833a80ec03bca5c3c5ed15d2a7857fe1bbdaba2f4eb095cdfd79e7527a76ffb26a27edc1203b60d09e07bbb0bbb0f6d1084990f6f6c955a626ae9d5d65e88fda4ae7ccdd636181b3fd3e05ba2f77ea7079f2f5fb7e91b03bfadbd8236ccb4aedeecae1113f7ba48fc7d9248e158972f57f2ed0f854f2a2a658583f964a43b5d5f036388c89b1f9b41eaeaa7d0fc2eeec29c0dbd3159c6c99fc1ba3bf78b018c8a492f39aab69a19e1a4ca49eab9da3096774bdba4e29050772cb4a6a94a0eab77e2a8bf23a7aaa05620cd74ddca8c498f101b9e58235367ec6f72a1581188e9fc32cb34d91e11750841d1d2ed942ac467d60a57e6b60219f513c510b04aa19962882e4af94e1127f656b8dd5a372379e8abb1a32309789ad92925bc247b59ceb329a5583f3c9f68f8dccc0402aa75befee965a74934c1b56ad04c588f91008fc95386f301c8ee5764a7c34f8893648b248192cf0fd762f42d83271a7d75b9f799ed97fe6d4eca70008ba48f490f0d3dac3f048e8d07f2cba0e233fc9ad38774434b9e6edf80c48141b740f808e3adb9824e54c60330b27d0eed4cd2e5a23f0e2f96946722c5cf8b0e13aa88625df560c48056e635472e46a3014fa995cc98b52f0e36464f769ca8785d23dc186037d1898e0164d917ece28ffe5208d9b31110faa224ac8f8bae5aa89674ebe3c7cf2ed7558ed1170e8f7b5e652baff50a114ac74edd03eb9701dd53c203f445c9f73c026fe3a37aaf00ee871335ccb09e4c08c1f8a16962f0cf532eb4fd8a3ba328e2e423efdb415e554f3a72002d8159c22a59cbea87d01867de2d04c27709bb28301a6d973d7ccce8d19aab1bbce207849d08f35fa4d2c200d1d67c51f901fd4d237b0d1da7f7fcaea62d5b99af6a8f3c24afe86644a9a6f3b961ae6cd97db40a8508cd943f4a46329b3f61bb128d90ba9d9568a07aea43a5332c0919268e201c1f06118e50f20d083f1dbb98d927424569476fe5bd2c1849a915779f8e20b1d1c46db22b5d1e0b611471cdc3bd798d67c1656014ec935a6454c309317cebaa6e743675b21c105d564d3b39af9d58075724e766cc3c270d06773aae59605d35a403674fbae4de11a115139e50b8eaa7bca99adc717d4676ce59cdf368ef73b5a56484c2d9f7e2b88f02159ce18bd9853e8c49416cdb318971f77fb45fbe88c4dc2637073aa1f1319f0775b1e4ff18adf62602a27927ef055cb15d486ccab2fc45dadc56f68e8a1195e58592b25e37988a5535a9781c74b2b04d8e52e17125b6b8f8a8cc1bb57971c8b3d0bc9b97d62331a6f70488a62b685ba52291bd42d9acd7c6d7c664b8de7ef1ed38f966d7fbb26dde11f4d03879d514e5a969ce61ae56158eb306338326ad516bbbcee12f21de50a233e6e5259bd99d8888518eb2b94aa152c4f36bd8acb09d5f60748e811e567d7b2730238d69c746bbd426b40bbe974989d2960eb32fd95076c2594d950213566390bf5d88e71458066b12315067ad69da96aae13bcd997b2673baf44453a5c45bc9f3b6a17ed45fb3d6f00b5c69936a09234994eeac2c182a08e1b32c12614e266d0e84419a8936ea45ed7bf761e090a3f830c3fc03c47c6404b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h51d98915becc0e2d51153cf8bfb98ee0cc3e7643ea11e01cefce5143df613f53211b7d1f707bdf87375a036b5d71c67c108a805f81fe425f4ef42b37663536bd4670b63fc40a2f3f7bdada34d0125ad92fff6fa114c7b483defa1337ad4dfd917dac051681e9752d95c11f6b7108cf9421bae189f9a933e5068187b90abd9f3022585b082fbc75ff3469c29ea0daca3b44bcc793dc48cb519c66c5d18f3c700279bcbaae989c4b3972615cd8170b47c22f5240be1f5735bec3bef2bad1ad795c70c20b08da19b2282636ed9a418528cf4a9104ff6d7c7134916a88071e961e8d0b99b55e8b128324b36210ee3246a3a989dee3a6d361aba78c8f62760e578b7a880f4dfd2feb2744c44983999c77bec68932564cca637f58c389c9947960c8aaf0ed914c02d500f01391a564bb0f7c1a61242b8f91caec634ef73c3bf34fd6a9ab9cabe425a0270ed8ff346b8c60d33738bb18b9c609a16871bbccd82780916159f4ad7b21bb0df5b07239e1551f4c5963a87d7670a62d5eab3fe0d8c73bc47b17fec1dd9c5325a0a182af7813b1f0a623122504b9645821353820b8e621ed6924512f7d9cfeec544038447d2e9248d902b69f51327dd337bc5361db94149bfdb5d8f565a83e4f8b5617b46420c31450a1c12cb2199c6789dae87f0907c25c652b27f6f030681f820895fe03f44d21c63b5ccc6519d1a2692817c03bfb87eb3f5e2be0e08f66a3f1f22424e15572c23b0ec88138ac17c651efcc5cf97e9481e79d1d3d58cee509626b0b787e65b872f692b6aed5dddcf615f22c08dd39d5fab32c296d3e93e3f0c976c85641773aeba1960a617541bab6a8c7782b438a66350f45bb125048027fdb961b70b3dbcca2fd0359220ffeedf40bd17e6bc89d6a3a1c3e820a9647abdd3708877a02ee051f29e4b0477eba13f91040e421e40fea142e1a425f8066efadc198f9eadb4b04085a2832daf21715fd3727b34e7a68bb2523188657a96bb4d8ef996d6d7615fdb9753b2718a78b29928f8a4c2f30077a4cd6bea39d3bfca2edfc9be655afe773ed107028ddefc2d69f95bccc7ed4657da094255efa5491bbd38f37f52d63034841b876313f280a20cc2978953b8d104d86889c02e10cbb6d6dc3a7380f071f60cb208a0e213ce6a73f96fa65a1cb2781966d44440f0a12eb0edf6b67a5c5840f49831980a6ad1584d99b51f4efe82867f2179afa150b1ae7e44b724cd57bcc140c5937e9667152d21ed389aabdc44862d3ef716c4fe8080ff0f3faadfb2d3b4c0c4c0d6aec8910590d274c65b1be27046b9192cafead54fc9d92926821a85661b340730e09765a1eda05d2258d597029cdb5be9290d616c8a81c938092bd4c6d628c068da027a1007ce82d7bfdf35a284c11244ad7c8ba89eeaf20daccae12ce5321a796cfc8cbe44479f68326ea144aeb317cbc5dc415191db208a5fad0abbe25567bba6fe3bdec09aed58f9fb6c83d19e7e5971f7ddc672d2eb80a10b6c261797325daae975015da37f092e53a7a707347a2086ec5a91a94af5a70038caf2ec2734dd7b5f9f678a6fd00546bb9a28e7e1e59c219389a417c8e7749c2b5cf2d7832b0336303c8e1250341bee95f1c95ed2c169c00f1d8eb8920f20db620f929fde145ef2ae10523c05d2942842a4b0929038450b75de660993a781a035a932b372ea21c577aba4ea5b082e48e0f5860e8898265535f0be026e2ccaacb11cd46e2d9a09d1aa26358cfb28f6b872772fbd9b62f333ed05bc9a3921c0eb7a1cdaa28959d598733c216371df89b272d261b67551f7860ee5d00beb3e1b0103305894475800f80b1427657ef5eb23bfcac89927937e14530d98696551d124b7990e98eefe18a581819e14397d6c63a718769b565e3d657885767f4ae06d115681235385ab34c57136af2c9d6fd8df582a4ad338b547f7063e68cde0c8384927012740cc42bd59a6323693545bdfba991f19f2404b6c83625ebfef1c6672850e39a839da4258780cf9dcd505242e30aa5398b7318d9240c132b8aeb2bd8007b26ea6ee678242a1dd275692ff38a398c1c427fd2c084a6951cd14b4f8739b3975b054a3f15421e27af07c58622800ad5352be682bc341229941c012b04bf01879e18f22d1a716f4d4b9ccdcb10c1e3fa873f22b74a5c2e0693a43ee1c785bd28e280c4a883ed964a33e2dc59ba6f6c76aa994b7340caf6bdd9be4040862f67ec2efecc904d4a13b10f7d5d3f44bf2de8f5c3b4cdecf03761fec406bc0446bbc2f222c3b4c25caf875275718eb3ade69c87d4ee1e723b89d544d06633624ab9195587722d5623b00ef1750c8c2b36be5be5383c793739955358b1160f5bf6f275b03897d3c49af7e08f2985902c02e4360361b67f63c060206401702242c192324b26439700254e9cfb8755153cbb6064a419d645d70a052e27971f2ebc351ed62ac20e02cd5a7fcf0ab69747aa2698841fa25c441b5436c931e6b55d059a163f6179d7f2dc2f28c7554447c7b1bb0e94fd34af9baa66e2f96f4dd613a90570889b1d332124b25ef58e52a142ef8b92690474ff3508bdf5ee6ff7499bdfb596165bcf5abda7546bbb1c55416c1679ab7db93fade39beebe15f7dad38797169852431f8e9aa3ad9eb54e3583ec141af50b0b991638aff8a03e440a68dd4f8a793704b50480eb4d9cbb64f5e60212b851c23ba9eee6bb532f08d7bcfa20cd738182549be26e92d66b097e34817c66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2a6e66fd5e529f27cc027d61d57f7de6b8b4cead31c0181f5eb5517db35c33e1c3426a9c136b558e3931d08910328f06bab6896f5ae56045c2734d88f257f47715267cdec61ebf9bf0fa1a7ac0f9728a2fd23c6d05c58c2a7fe1d40823053e0a105429fab55d83571dbacdbdbdc6da74ae9272d00e6ab3117e63e92f2e0fc02116cf03ab7dae2546b542de03ea11d816460efce26df877471cbf8fc3bac28b55c4ba7ae849a1068be81a6f51e036adffcb67b9658110b5c67adb4ea69d0391ba67043ea569f99432e27bde10e1072483631557911406007d043be8b3a6f914a2736f17c7b3e7244250c77a43b9126d50f5c28965a5addaa441dfb72e9668f746a3b42e9d16066a11c259a933d8d19ee93511467f60b84868a5acf69bec8b069b3a0273aaa8c2c544b43476641e58d675c7fab4d50ccca9073d1dc93dfa5babe206b1d7139c884d1d8b05ec2cb55d6e998592260e2b6e37c0ed9b897cf74a3aaffa59b107ca5b27be4275da2ddbc2485f6994a60da423a7e5fbaf51cfd581704acc37ad879c62ba55b2ae9c0060347258f4125c085d3b493dec801919fa5658575b3c7fb79b08478033ac5b68be1f4619fb7aace250ab34cf66b612bb3fcce42f984ca4f8ba4caf5111eea49213c2307b0d1aa3353d8ad0aa240d10d14dd527870aeba5265625ae00ffb1a4d9372b52d8a2003142f1f843909bf78c7bfc49b5d83ba47533b67520ed0e1c5572062cb65ac763fccc43db5bb02ee414ab0059d130d799389d71c5c0ad7e7271d2fc2431171d1ba8d5cfcbc246dcb5cb1b3f6151bb10e1ad589b01778cee755c1a1afb645d469a7f4d01f81bd4e7c824ccf8d93003c49301e238f582dffb5edddfe977dcd09478c63a7db8ada4c819847ef565ede9325a78310228f98fd005a285f71bb366fcefa420e787ecb4ec3977ba4c23c8a71e9ddaaf48564db503ae63cd9be924385ed4bd6ff9246ebe1eb3b9a713d661f0f6e0882534a318fd48c6b547bd6be69a1b923bcf40d4360877eced762db7654df3cdc1cbb24c9bcc503057ae8ca0423f2c84ff3a106f5a78aa4a87fda1571c2cbd5488e2afa84565a828d3ee23c68bd22376ccb2fd8174c7581b1b6c29848c670c0d67922db77f0160042d6c4720e8a7dae1c9791315a5b98d9aaf99c83f91511bd23e56ce9563b6356a3266feff8b64825c50f98b0f7f88a8a01a6087c7d4752f20dd6f2d5cd2e71b446f56f907e753f94295b6db2a721e778293fc83805b26801a38b6030f2457bbc54b12c7315079b0e3590077a6caa59ad9771ab7fd4a10d25d2901d765920b66edba966a769c8d225f929088e812368463e4aba85861608cb5b60617c01ed0c04b163cceaf4d8bec8adf3ac2deff5d9e8481f5c1f3f198b6756d3f1bab7c7e306cc43bfe5ad02e12b464baa5b8ec7f1c6ee8d8b47effbb8376cc4a192fe746b2aed54c6962e5952d0072cc1ef43381404640333fd095ed98fe0afae70f01a31ed5c130c689b60a15bfb729b8b7223edb14d283f5b0c794469b918fe96ffcfb1158430b31d2f6925db20e51f8a74de1c530f09cbd501710514fbef90593d8c2520fb184302c027a2b84155e2e16cfb637d9e6d3deb41cab4522973d9810fe7326a5f8def8892dde185de96cd9657fc4f98ceed7fd0b55bddb52cd7fdd403d689a53fc70f5fbd9f151f75801f4a0914831f1045c674086edd5c744738137ed4bb0dcad82b0c449d727fbdef1388ef21e9744c498f9f70a2da5ee8d5b05a2d8ece284bbfdc1c5032ee8f0f00c13c7dce55ed672fe8f5e5d1e1f5f4ac0a5eaf74874d116af36585522a40ff6dee268d780e615c39f63ba2e8ad98b78a0974debd3770caedc60c5806c9a58781628d922921ee95bd8913eba141cfad03375e2ddea6d5556d96631fd099fdd0345cbaa51fe9b7598899543ca132711d2098359866b7f2d035c6b3b51980c34b7ec290cec7650e3b63c575cc6efec09aece8450e04350a5e5cd1f04954c88c05024417228268825fc41e9d2911f101495f037bbe354f2e91c1a86daa55a55523266eea7f218ff4827dbd0384d868a2c01725a67b9950c7b219dd4f77ad4455cff8529902ce41e1906717d6968a7a1ce0b013ac731a570d816aba9ad6a65e2a5b766e2b572ef78ff99b4650cc70b52f34b80c23e91aa8aa672b7c0685c833b6138c2bbc21ba2a8bcd1bae2bfd5d197040d71707f8f68c401de21fe19a4196f43f202236c79ee79f32deff8516cf8de8bec63d678be7ceb324f9ec7b5db6ca7b572fa897ed15f5205114fc1da9503ac77bfcc039ae4416ac7fdc425bdfd161a2b3e409a45f2bb2d38ccb63cc88f9e447e6af21612ebba771887236edfd4721fc353f709de1a385359fdb800d4898b0705141069c8bc51acb103f55f9e0f471d8053d8da83b3e8e211d77507ae2102ec6f158309753a478ca3f87521e620b32019bc7558e90970240f62c27a12327de3503fc3588f9482d615f731ee7b79d61d45edf530c4700bc3108c40e6e92ec7e5dd081edfc0bdd02af978bfd648f8c5af7f3af1ae960dc567437ee351b83dea5ece113b3344fd06b7ef70917d07227bb726bf5ffcfbe3ce3dd697eb38138ad737da6b67851df43e243afc2f7bc1bbabba0ba077ad450d580d706cd769ec38a14b3e59aeecbb9d198001d5d264683cc0687d317112a0731e75508140fcdbb91ecb60f3f1a4f70225dc0c684c4d75dbdada68f36473917f8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hfdf4bd9a8c789f58533e19c78f29b1ae865947709bf682061c96ff3a4a5077e6e4699a6bf5c5ef995a108c03993266579e219b53856e7eda1bdaab29608c89e474aff4fc2a58a3f7408d22e8648deedc5b8030a56b162fbbdfb2b8159ba6ff82eb3d2efc37fe16ed3fee6daf37de2f792657de0a28e8f1b16714b2b5ff6c38a869967df18a5d70704755735d94138b73dcc699d236b81cce1183ff2860706bd67b719997d7b67aa2920fbcb85305115b3a53962c495000a47edfd6bbfadcd99308005fd9d25db77981247302db898183245aa382c4f2d6c7441f382d72d1bcfa36d96f04a0e6b8af0c98826861ab9faf696be949e949f1970cc427efa96a42bb7dfa3b9e88a188b172e2bfe0391b123d8b5c4b72911952e8103481033afff97043fcd3ba982da3d80be585fcbd5756c2746489433995fd89da1e561f151e494d0cc271597094871b749b15ef40b1453e5173a9876a38e2bf957098bd0c037fe4f626e26a1f00211c72c81178a6c80ad5b9a131f5da2d0ec701af232bd61aeac2ae1b810938cee843237b6c81fabf670a6b937161169793e7c8f263f239f33005fcdc2e6bb2f301e153bf61d7a52f2110648a1f4f9b1ec583fdde36c343a5a829091f844965218e88fcb2468cfe90ee70720bb9251263d767ecf1709e5f66bf008da3c2931c83babb9f2c616266905a7445f0ea1468a1040ffb235256f1612398eaf878981e3a1418ecb069aa7e126f97d15257d3721ae8155c11bdef5d3ac1d9d57b28fc2ac54a39e5dba00b8e24d4bda3d8a9f1bef4435183560f618d7905f9e486f71b6c3117e6795d75a13488fbce1af78da7119944a01be6b4d476cf78c70fb1e8979220091c51f013ef6877b11036bc8aa3e0bb255694c93702af97db7b23e6f423efe1d474c3dce6711afde5a3e2fc3498076e3b74be87995d4d407c17a6898364d9ad4bfc8be67fa1b963a8c7609f13d875fb7f0315dc6a12cdef6ea13064f234155146f7faeee9c53dc0339c526a94081028a7dd0e8f9326a31aaed911f3e4ae0c1e1762f9181fb01348365185165d73076b06764afb7e7840fd90a41ddbf09cf28df9134b4607b9bc082a138aaa5ccda1804a32473e0b9fd5e3ff6db9595ec8245b646557913007d430169a7e4bc4c9f926d2c3c01a53845faa8aa8c20814ff0f30d789789e21378f20f041d18d63a1d3a2e3f880e955b4ef5c0e06f42fb63aed7daddce29c3a248d126fc982850bb712b60e8934eff7b18a655676340d0a41f127610fc2fadfdfc7f66d1c471ad3483533d15d227716e9daae86fdb919c17b36eed17643fb8cae247f0772e3a22f26fb8ebd373b2736e81498e853b287c1799192e74d84b0737ef4aed9967827bf5a747eaf646611296473fb93810cd39e88a4f4196e5f21602f80b3bd4352a0afc8a0771ede02d9f07e1fd40c5b066ffed93ed12cd5cb6e28529d3ad70ede02399e0a2b8cf22a0d1650f40cf2a8290e960da61287f7bd9eb3e67b6c779183b7ac3e9fc075ebc816b2e5a3e5942b5f1b2828b8521e00e9b624479c77692d5c66ed4abc7a23736660d1a0ee3564ae61cb747af270d0832f9e7e0f9640e697f698a510f02e3f8c0606b524e1eadbe2f7b28e517d36f37008205f34a694acdbb57a2a73a51c027e64d716d4537746a40eca9515fa82403025dd5fe0277dfb480ebe7a7908d416827a8f6c99b58946fe3294b87b70f5046a13a9ff6115b89bc9fe1a92583ad1c3deaaae65ac8af7f6d314d05d4161191cfad566fae72851fad3b5575bb8872a119829db0be3ad2bbf54eb4e620b837121b686c09057e59bdafd160f41630f0576fc9b5e5ad9d99af90f685fc64f97db0f5ef4034d3dea9d4c673a0a596600cb4b8bec2d537d0f6d9bc135685641525c4e33f160846bfdb3d6bd5eb5b73cbbd1cc3071101e762d73bbfc89bbcdbbf586aac97756bd6e4ce797302cf3d46166558036e321c3e9d1e3577acd686ec020f4babaf0895e454f2ff8d04dc5cb0c016a5ae069cc881fd0c8bf76f8e8512786296fd4fa93864bdee1a1c205f56bcb745bd155b875344bd55fd720d9142300e8beffa370cd57e53d6c8136e642257c7ddfd1049ec42929b4f729784c03591126f971614b3cc2bba1292096eaad26127ffae84d0c9b761be8d463b6539edd9bc26959b2777464d995d2105564797481d823bd46dc5fce6f958188fc4162be94ba6d12712cab95a7fb886a560fbb21f9259a4536f4aa573ec2dd11b76e9bb3f36b209d0277e7383d12989012c82c4c9e786bb913b33a7574907c2ee5f5d6dfa798355394731534312a5a80e552dfcc4412e781b0f286d1af52651e9f3b6c3567a1d63ee2017777b5ec5e44c09dab37e33b1f2fdb7198a19d27be2fad97aa65a055ce001551e870a1affca3ccc1fbf45eff94002b838e4bf024002a56a114d91968966294d1c89670f57e737dfd39cdc9dcc9961574afd7148057d369bec3792b45a82e54e57de5f89e3b2f7d013f45e25a09f7a2126272c137abc51c66642bd9496e26a9675622d5e151401f1b7f845f85d89ab191c5081198c2fe97b61067329a3cc5fff69f1e2ecce390d5670f494c91d85a5c9bbc6199f42f0cc355e3e933aea3ff4678ddbcc726d7aab54d80deb2b4abacc8b5007dcee584b174998d3031680465ac93f4a0a2b6065cf12d68e86a9620ead13b1de53e13b58b3850334f4c936571f9cd82f4e00eb39c92b543c4282ab533d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbd1ed49bd55cde3fc113fc2e59803ff7fba17a2f6248afc21ca89e159c73b9e818049dee9ed4ba661867bc39cb48cf67bd04df72a19886e0254eed0d0f4a972d23f164e9360fe3f863bb250047302343cfdee82543eb2c9d329e29bd467d74b15e155d79085876d5f661502031b9902a11b3fd2a8e2a9ce7ac226d46e66401d85ce52f44f1f58726793e728c1bddfdefc01be2a690e95ab2e41b2383a6339568cc79decd105e39fb44ce0e9020d9f4e4e16779472716f1506f2be3c3ae4c3ac3a7947d2c36b46f9051d351692e16adc71e4869bf7cc5612d03d82caf460ea76d7d92aecc1aad232e027300a405e00e4815a3715d1a4b7466d7be98e91feb89d1545ecee676ae51eb0ed57d42e929dd6498c56a38cf4941ed6977cdb04fb347a67573b7458f0e90587e0b5315c1aa037927ce2697680b38e4d0505f96e5571be5b892f43817defa49bb49be5d5fc3f0efe850c37bf50f530c0cf664860dd06f019a08ceb03d07ab25ff1b0ecc02f10593a934a4c17cb4bfa51b2126a9ea4ec848c99e46dbc5037f6a0b325c06d32d5a212d29fe15afb9b9e3ee800708b2e868a73573899e246d6a3cf13343aa84dd3f91dcda0f93d5a103b08e59e0fbc4f77b2528b4a672001504662f16e7a6e57ac02dbf000d333fd4b59c9f6b5ccc02551e0d95a511c6022e6157cc19f863f560410668125e6fd044369b1fd9f9e791c6ded418b55eff9abbef5f189c752be571578cfef82c675dcee2430290ace3ce8c569280e933b89f24dd026ab596fd09c4e74eb91ea6d30a685b690cbaa9ba5f31bbecac65dfbbd6aec1e65e8e6983cf6ad40a3af2ea27ccd0335371470a5b3cae2ee4a8b51c66c53403adfd4fce1b6cfa9568d493e61bdfb37a081e94c26295458627636038f92cfff3bd682a482fafbc03f32c76c74770071566729eadbf5933f52d66d2e8d1285c4be863a20436c8000af6e95654f6016024e4973925aadfb9e2b52ec6814b6898e84e3d76e34796a1777a8541e1ee36f320e1e3642571c80b2ab030864ea8f2e0779f1afc76fe8c7e4e04ce2b8c1063522562c77cf12abc032cc8d7460c0dc849f112b4bd369a591165d490fdc672fde0b86091013402bab8176b7f60924109e596260958a653ac0f5f18c239dd5c867d2d1038b516d71932b16e53d43c1d94cd2d89dbb600515b7c823e21bfd7f95dc6f4afe26493c0fa9e24ec2adfb5fe1e15335abf14b152f3b6f56bf728b1fb4683d4b1fc4d6289388b012accef78b7996846f6e5e40b0f206606f39211c78a279efc712868128f4a4f1eddde1ccf8d50ae1c86754a0deafe7ca2e73765409c61be7341f96bbe251d3c13cdbc656b154d9af7b1594b661e3b379d3e2616a9cf58541c82d666b8cf88fc03feeaac305d6dbb656f22ae8f496def54bd1cc8f7c0b44ac694ffbee3fb3f8d0f10a54f16f79d145687bca3f74decfe548639203e3c8e081de3c3c4860aea7f5f8df7603827381294db1a8169d7eb4086abb154c08f5e29070d332e9dbd436c4fb5852aeb5461b3b3e15505ad49cd7004c48f0997d8ea1b7ce1e6555a2223de2edcb64819b42fdba01f8a9311ea581cee2f8544af530f4934745f4a79fa4f4651468aced645eb1d9e9cc7feaf767bada2304a04eef44ccaad6cf97891b6c6b50fd07476987385db9ef40c6656800745f2152bad88f099478bd9c8a10cd92465276632a6b15b214024f48dbf8d3a4b0a7446a19dbe56c63a68186e4f398b173c89687030d5e2118a74d20fc91bf9bf8ed45dc8f50a3e29dabd1959bfe436518c31dda8c81ba49f1ff105173f800cfb61eb0264838454262b71bb92add4d38e06da671115905e1e396f749207908a06d67b650c766a1e5f1ecbdefcd6869610e6eda07ed9a4a7f0a82a5b9dcec6922f54d21c4c7cd78f70f40a4a4ab9e800a60adf9456c7bab01893f5fd25087640825a07876169231681c85ba1adb8522661dad33359d351c0cb9a1631562a12d74dc2f35070e35f79bcc8d7d4fa7efbdb15237f09f767851a7c9239241d505b1f3e44091666347f2a2a62637573cd9ae3c465fe676538dd06d0bfce9d58fb656a74aa6b870a60533e43341a8be725108126bb44152279f88b5de17cefd77081622c9a1825cc9aea4887a604037344c99a9d40a600c28f0dda178d8eb5ac024a9d13f9aab470e9c131160cabaeeb75fc1f73712ecee6ca90309c4b55bfa8beaab08eb205b697ef9134b57d4ded5c34e9506e8c0fe53e5ce8d1ef4006842dc362f83b12f34d22937ad513f8512e67e34c37df3160e45ccd8bceb492537d4f9641edf8c5e2fa136c28182ce759a0b8c033d83dbb47c98065f153db2885b013b2850889078fd199f925ffa33ce8c3a2da9b157142f3e748c24ae433c3987cf46742ac6eb4c5ab1dc20a2d49b84543f764c4596c4af79176c95fa23d46e6445596655347124c2484c696ce66dc60d67d4ade24fd1cd2bc1a58b80f06542f7dd012ed1317e44209b7a13db4a5e4bf3da1d4d117d9bfd973bded586bce33a919b9eb658e5cf911f9076960db4828224c68f90e599aa103dabcca312937f5a83ce9e88f2125b6b3c7f457a05704f26145f8d71168f5c30c93be0be8d51400f6a0d21b4662e2289a13fc58cbd9d7d41f6f060311621327fcdb432f0795e37f6fa0b04e397cad9dc9ef6d8bd76ef514e38093338c7377c7337a08a679842c4385de98d718246f51aeb9182838aeadab8d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha1350798f0785f787934d455d58fd8aafe136435c5690b556d1e28517ef0c08e076be7ea9d3177b9befd39604e33fd09fa59d4fc792c627e272440cf9b7ca9f98f8c7019bdcd79e84e52d196e5c1eb835d6c02b62038cb71712e6d3364231f23e14ebda3e2cb00ff01928180e4bb5ec499dca3372eb54b2cd017905b51b40f37f53904e102f80a6ae4aa49ff9df75a474462489fa3a6ed7a262329d4a8d03301902ccd9f0177ccea459466769d8faff0d1f97d591b75f0d3abf6fd8305a7c0f0c085d29ca5d3a4438a7cd36729eac2aa02b9e0ff478099b3865fbe8462038b096c96a4d581713bbe9657dec494c24b2a0fcb7599949a860532685703fe480d4c67e682a165cb263dfedc291b4e59703f915b74ad943c041139738af2faa09b78c34eaffcff58b3f16f698d3a576cc5842723d2169627cc72d11122697681f37adc5aae4f61313b6d14803b4c22daa7a90f5e3763be1a4dbd3beb9b23e67869f56a5297d9bd6f20cca3ac986210619acf2e5d65de00a69c36264f22169ed2aaec35cbd3054810a3ddcf464f9302afa51cbc6de40c1f1734efd722bc3540a0a4ac78216238bac370d19502aca6f518f69eef858a1b3eadb9faed703d23669d0573041234e5ed08cb73271c727528b2aa960cfd327d3a05d85ff5f1b1070da4f7658a86e93004d19d05f9594ca2a7efadfc3bf2315f41a66e2a9bc074051e785b1e6210ee1f2d40600d19fca41a3c0174843d9f362ccb0505e1418a1c7172b6444f6f63500738b02741873931352a5eb113d878bcd36d57a2537c3ed843f58b69faaad3940196dfc64ed8fc49cd36a79305256b9a52f9283758eef85257ec6e6b514feb26e9218ea6b252cd2ee100157b42eeb0f1e3263e6b61b40bb4997d7fb942f8dd359b8e31edcdcd124881713e4e84fcf17c3e261b9162242db88bdfc39eb5e8e634bf12ecf5e3780c885a7ee5231943c96b9f9882e6cf14d884bb3bca28914f58e4c548f9eafa25a2bd67d76d48c96e320a226e1cd6efc092214942f3ea68f63dfff83d6c534941ae14a3b58ee69271495a43ad068e848d3154c99763446ad36e2e79f1072b493919a4328c98ebaf2fd0a20b31252354774315259c88dac6fe7e3053278e3e7c8b93ec0ddf9776d912dbc49279b57277e248c47a84c9c1f0c8da9abea2bc988d313b0fd72d01a4d314e5236f2bcc59e3270a05db02fe7f18a5d173ee24c075befc84ff0a72473e2ce80cd428d6dc36206a66b8fab869c0e98c9bdbe91adbac079ce486cbae03d180f4bdd5d6a6d85a8cab87cec10cc3b085106aea5365f1e57eeef14d6fc3d2b1e153aaa1f481dce49004f583c6db81baa75301e776b623d7778626cca15658bedeef378941438ff26b09b8dee6100926ff8ead8c7275cdcf25f3c43e01a60076b864b979ee0e338279445489ffab99dbcdda5265dee330d4132fb89c2fac48dab6e3402282581e3774e743dda43642d3e2187ffe69e8e40eaf0c90b5fb2229d6893252583011581d2c2b3e3ac35b836502a66d4fbff496697ff4a7e6b59c19ffafc727576e34879512451f22bf8046c9fcf2fe71c1108558f565ec8bec628616961d8a91d1f32c67872c1c96c105604c689ce1b863d0e926215b0a84d2042e4936d50755ecc1beffe34e84a8a1f95271c8648ff859d9475bf8e0ad5ac23cb30cc4f3391725e6eba1661edbb587fdb25a0ee5590dbaa5b7095ae7c39bb1d70334630f5d315948d711a4427cfc852eb8a8f2fe3a61dd7682619c0d3ff015d32c2e93bcd1b86f8cd702a66481900034c9e66338be05dc9b840fe0ac83f11adaaea055ddc21925f901ab0e5816c3d0e5ee364f4241312a9212d2babd6ef432eacdb3eafe0358ce74e18c5ccb9be128263bc53f77c2c8fc56e9e3a63ff23c6f470384ffeefd727e43fc1cf2bb50db1063f7c0b188265ac263963a3e22a4762b3de8c1969c2653b66a4d19242acbae41ede06898c5876f514708cc09d18db38b197edf2beda183a36ad06d23fc321eab202c9166cd5612f11dfc0027c1f7b8ad8ec03c7f410b8073c024ba7b14a151507ba5748da26e422eb5486fc38a704efc829e427a0261cef77d387f6f76b0c508cc69a2625a3c0ca00d52094c8389abb5f14bd66f97f55d4e71ef679498596df73b0467e4a2534ec8441f686336b9578039a1a46f320b653fc9f50754121b34d344061c5323ff99779d81d4d73d8e51dc7a8e7c0a1a9cd01a09fa78155800a0dd703a2a5bc63d6bec928ae47f36b3e92a122e4057f20ff302af51665268cf4e3cd54a2275323755debdfcbac06a19b9bf4bd83a047ba7ed4daba8cd0cf5c2956fba9ff0d49e60441553d2ae7b307e39e2ed712657093dc3c0d2042e1cad950d7a9e1f133003524020f6c9f80ae6b3fb44598e983733f00c10e99f454878c098c2cd85e86830f1a755355a97a24c5c096c02d5740cce677165be0f09e2d6b0a20e1f710b50d452b1d3caf29a6f127a592abe49d5f55f325e6d2288a7f3eff6d588e20ec1b20ef6e124a795b5e53be451914a1c71c79035138cd3376eddd6e3e98c0f565c99e07469e898339c5cb78a7ea50b7de0fd3eac48bc5d141805289d940730a02472fe6e6e2efcf472c52be79f5a1ea851dc656af2b98a4524dcbc1a1cd6d49beba8b0f02f526d3fb26d9bf6314a6eec984947fb63fb43b02f505a04a7cbffa86dc267561298619e2bbb7a90105f6f7025dae12512ca7dca97be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h25ecba2ebbc8ecf39e16edae47a14a7499d952e2bff6c44594764b89f447bc20dc1aabcbb35675c99993d583ea3f7f72fa3c941dfd605cda772412aa35973a1126ad11d8f7b902e9087f139916ae8ab398b877a0c920b9dc4489c55af03b93e9e294b1cea22c1207a253480facd10df4a60bbcffdada302de01d1433a70b63254e89fc6e7db3af42807539e289e6c5562ce80c6f00dfb7c012439f7e49240c248c1521596d8197b2e6dad5c74fbb74ffaa3012446f2fc2354e4f194f49ea2eca599d6d433da13380363763019e15adf09cc8a17072f8af3eebb35f96007e3fc98b84ef5e198ae9110545f928595b4579c1f6c9337355762194d372537b16b154e15807c08ed27d62f838c8f0cbc8d040ff54f37089ac6495d3b2c771f3e038f15d79cc33f58c1818884e5511b35aeb9d4f33bab2c1eb4776ead9ae5d527723635b6e9a7cc4ada0c10714328648ae35b7c927b5945555c4038a34d8663dd50c6b481cd8c0dd478a392dc540ab48bd222d3b2d23023ef4797129c94f20b980b9003819822d8ae8d461804fe75505732063ace0827a426e5e49195ea008d76c11ced0fbe64767789e366055cd89e04113f5ee77080aef5d697a361be361dab13fed22648ddf3c2227f14a007e07406b908640f5cb1f846529b893105ee4f0612229f6eddf3ff16d47385c5aa30eb9f8164f45782cbe98fe2d9dd5cbf7b460e58c40d9d39af86e74099211a32a5e00307cb8e388c758b4d38ef9e3bd9edba31f6166ffb0ad72283d64af9a896326ce156110e3c5c89a63db3d66145eead595ee126f2ec1048c632641686f0b781001d861ff13a597141a841eaa8b900bbdea496193599ab7cd89027867c31ae4cd93c6c6d0065c91cc8701257607137928df069c62c7ab49423c1438fe188ba5d6384a6aad888c8bf580b27e66c3233d840b112f09053339d9b26523194d9d31e39f92298d12a6f24c0e5d0a4a7a12ae2ec8244fd9db67d910fa4e0bc11bab821c29255ea0c811d8c8831ad7a2e614cd8f3c71f3a4883d85549a079a4cbf977888616a2206f009097961f0d33f08a5bb5aaddeafcfe052a57d552b5b28adb009e6b3b62c66fd72c3e9bcfeee53e2e7621ef21750c5eb7733acb98c807cd54f3e5ec4189dd59fd0ee2db4531f4baf442b1120e798a3be14d908d04347953b6a7e22e5c798e2b08ef666845d0548ec69af436f91dfd0a44feaabce03bd9fbf351fe159d72fd168308e3daf06272a031c03e7ca4e2e17d430c0cf07d417222a649a9ca8aa6950418bbf9500ee5ead4482a3373bee2e49b7be5b5414d0590637b9d7da82f46e6a30322de5ff145a12a4ff8a94e7becfb05a2de049f06a5fcd31efd6e3bb84c8db0d6faa3db75fb5f8a4ef6a40f7833889e0416e3a12dd8d8b12315d25815690a1bc16c2e919f6df0d5cbe084a46b4b0985644e67835844cdc83ce1abf049e1d616c6652d288d091ee0031843ad198228c434fde9305b94e4fc411049881d53d6022699c63c16572a60a5b9f8ed64fb945df8c05e0b9088021478b307187795348a5493f33f2c7b51090db42b26060191291fa945c831abf3e7723fe471e5e3ab0478135176479fc14a79acb84f251cce500d8980c62d5d6e85259bcf50b439ee9e3f038258df4fffe50961b09c817c2fbd4b714170e036320a3ccec1b491168246fb26e06257fbbd1e003b90bec93c1b8898eedae3dc2b9d769fb5b93a37ff8fc723147e8d5a99bb543b77e262443d118a5c16964ecf7a827f2b7d40ab415df2cdfa4539902e3671bfa9126efb8fa3e827e53c90ce3b287ae2ffbdd4dcc112d02376205821dd4bad3d227307ceed88dfba54ec97ba9f784d633dfdf012da998014029a214666327d97d4f3112fde221e03e8d5903f2c59c1245989419aea3f80b772e1cd0fade6f48dfe201b18e16ad8e7bf18be706f7da21a45272394e835d48b835e3887386b35955dd3c94ad9e0f2eadba99fc5848eea7b03acbce951b6871537b391a06a661304046a364aa08d66ac039c3fe7aa3a19a14a158b1df08ca074eaa43a7c555fc1f789c7def8faf6913bf6eea9278f2c14be25622373c617b1b674bdb19602fe21b744c56410dacd70fa09e99c3e5cd2f490def32e2110bcbcdb222db62e833a30fc25edbe8226621d4445d136734ecbd1eab9716c10310d4512b05c3ae2ce501f9233c40cdbbed9f51c3cf429ed0f2cc280718463a34ae96c853f473ef2accc957c2f3f6c41979487c330d15df5252d6b3ba5d57e97bb4eacd2107db44abc0032b352295c46f0d4e62d00ac22649e9bfa9b9ac8672d4131e2f3fdfc7fa81b743d4ea77a377b7e8efa236115de0c933b49569aed44928066b3543df280ae232dabbc5795470b7a2337a8438a499d07c23969c0374114db0e4d2e752bc8c18c5857c7efbc17b529c29debc21ef5804ed0a19daaf5b1783622fb9b3645af16052772d59a73cc57060f1c22c81362d855faefe25419c946e8dae4a3f4a6aa1d17c6ace39df0669f635b050988c818a43ec4ac87163352add22bb594fb987dc7a96ab8145a90c375f25892f9605f7e795ce2158aeb072657c3e51aea0d784463193f860470e7b3a41f63a2a6317b00b9eacc1524239a7243468df0f24456bca5d547da67711f6e998eb3fc5b853520cd1f98ab590027cbb0c622655f8de87f0a5a1011f10f5400af53bfc7581140be129b96d28f0e61a6c672b42e7d111c1e2e669f400;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb7d86f19c2a3ac9ee980094e6af876476e5a4d4ff31e694db69422a95ac65c53219719538062d9d15178a3fa6d25c2a27b360506027a0ebc9794c1cb9290615c1091468f20631b4b34c6d60816e2a8f89c7fb892de3d02ad5e73e574c5be85562569f2783e865bcfbfa9cb3868bce747e978c8121afde05f1a9dc7ab44666c7f7d095d415010400502c7bc1c42992d93ed17ed63f14bf7d98dd56330909b38459b307b981f471f19140687ca899819556c471e81679e1bd1c1b8dc1cbd39407e0fa9e0b47d21d8cd6253843557f06d9034b9e62f857a53d4e3747d650c2bdb12e88998b19931d53fa4f59ff0d62732a18eba04029b7aaaec49e9152590cc6c8d9ff98604f737e9e38f5497add3c5e238f01e1de398adc4ff250de6cfcaa97deed7f02d144208de4421e93a0ef069f5cee3e6adce65912129c69d87117140727607b7942eff4f289055f03fb5395ccf1119f51dd6406a160cfb9bc616e84489151548683ebe5f1a4a2154fd9d405e9f11308146efd2f09624895e0ca93632ba53e853914ec23763e64a1c707a0c7b8fb70272778e3a592e3db5b9ea2b030e37119f3e4ae90209c69563da836507b96b3469eb04c29855738cb0ed551f3f65456770a6b0b2b6a60dc8a9df3096c916db25dae6b778a244c1d6594eecfef41bcd914112971c8a130bdb5c3e3d00f24d0b7ee5b79be7c2e518b30e6106ba8f5c0fffcfa86760d07c69bab365175dd0a49faa90040649b3e80a7e3ac15eb84d4d0b8dc9f2a9aed1808f8b1cea948221a14a9958b6076f8addbb762d7b2874be910fc96c407da2ea6381a0eb5308822e8f9fefaf1e0b43d4dcf096896b18fa0b2b46596da190aed9d1e00c02fda6058e1e1228893727ae8af625da73737ab26cfafb025301384eaefe229a72ce1e67895036a7f70cb941c042eaf48ddf755b412b32ec1a2ab80b204f31bee121ab31ff557805b0044f8eef8565125f4672144259ee22fcdf0d9b15b7d00db221f26d2b74c130faf5b054cca57acd450108e287f8f09d87a5c5d93536a6b7873f4817bb3e972999bc69cc1491ee9e1ac973201d1657ec1eab7a777ebf362b7219f3fc0ac677b16230b63fd768bb8fb5dd0c1c1361590377d2618f1e4a97ef7422b1a75c59bb8cdf5399dbdd77926798509e22672fbbf38e1f7a6eacb22099ead5a26bfbf7e568c7b008296e7b7a44f3c6306f36e95792443b8be1dd5d44bb4ff28aa2138d3eb2b6f6f7582c4c95f07c852835d0b0de811ac0fedb4b238678998afee1581d6259fbbcb9ea063b18e613ad07eee0f8647496437b6760202db848980ba342d9310d7627d51fe5be443ab1ced2ebb289891923eae148a0fb63cc9ddede8c7646fef0b2fc0d64ef74ed2bd223097e75e574882542393d0444f8f0a1faa3078382456a3de73516dfa954c8d62ea1ef72b3efcae1d8673094da9c1a35b73c427f36116db01c061093ceef852d547e0dcf2970e8df346258adb459122ab4701cad889efdc75dceb8942989413755f77c0aa1f705f50e8d003048ee5f1d2ad69b6b555b82c3227158b8fc21dcdb2871bf13257626a2c15c9eeab165e1e4e1deff3c53f013b1e50d05f1c88e5d7211650997cc22504620c887656c389742ac45a47ed589b01306d5f5f8978872c725ceb3124605c0625afb1737973dc61686428d262770863658dccd3e0a3e306268a591d2236589db6783aab5302cef29ed03fc6b3afb9d2e19a04a26216505741fbbd9b08971c9ba5be4d5f122ee4bb3799fb42c6ca4bafdff70a10c73b9877e4304c400e350d2bb374253ec6e03a45fad30a5c29ff7e655364a88c445ccd703d8e7414b798cd3b2563ad8d36d5b0b4b4d0e489ee8c2ec3c6116f942096ddab55b4dbe6fd16cfcd7f13e56f6174e7a57452b640ed6041dd267f08ce581773d2251655cdbbad29a5a8ff29680eaf11519165eacb6bb62fc65530ba6eb817e3e6212981b3559f54c7a0f10a6cdf1c3126b0124a1f16670eeac23735e4e7b8b8673e5d5a04ff0c6ab4ed754a6784e787cb50d292a4bf78d0cc01d33de033cfaef87ffeaa83c439e94a5e8167cdb662d4a802a6a5eb358b0de52f6e88f7d4b8fb6edce761bec909973a42ac9e7670d72f6ecd19e6c8cc1a5c52da97b488f088ce916bde7d64d7b4924a185c4bf058d7a8c54f180f3e3152ada859950bb5c7589b61d5ebb7bf8e5c8f7ebf5bba6e55f902d605a56e6a17691f5859b3c9b8e349851cec7f646a95f6b2f3ae3ea2942b0f0d13273d125b3716246cf893f497b521b30f09ec0b01e2959ed9d2ac62ce3872d6bfa66cd3b505aa7107573d90cf0a0678bb17d9a5e6eb27ad75787b75a60f5b95e1ca5a8d548174bee8c962ffe39fafb0888f8e3438ee9a2631d25c696af582c07b1b6f62a5b3409c78c539f8543500817c58be8e044a0c494ff9ee2a23d1070ba6d8e50de31118720762afa57cdf22feb3fab2fd6889005aa980211475925c2bf3e1102cd5f479075edea239aa26a8201db52ade56537f64d1387f998d86e845d11261a1919717f87a54ccda6952989bfa83294eb3e40a9c605ea364ef2bf79e145642714f1c8881b8bb804aef706300997bf912a6b675959f3c8308df3a4a6f58611fddcdadec4688cc8930c89460fc5ebffdff17206cef0241cb925bcd752d992c3ea140f37524b481882bb5cc274c1ba44b7cc72ad4387a1ebc65f539e99aec2f51b39e8d26b4d30712e096f013286;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he738248ee7f7a34de2e2f7dff7a02e6e0427956eaed15c7219c09f560c5c2f2fa28a4b71eba4f3b918ae384ea870fec9bdcb8b5eeb1c05745cd6fd62a8801a37e8fd60b588f6c6813e8e4cf57b2753095a16bc7732469c5ce965e2cf1df7467f0f48cf4a940adcff044e64a58091e6f3ddc90c38db861d430457610bd04458d94295a5fd8ca1b2a6519dc00a4d279dfdda270382d00327689d795c081b8fac609b518ae49fc5dfabbde68e3937d628258b02b2ec8d23cc422c24de763efbeab0222d7e21314e44e4a1e74b9e5e04128bbcdba11a8d76f810aa3f6995ef0543c321ada3c943b7d9e989f4fa15049c57c2ea9a08fb45a3f128f15cb0236d6b7c98b3911c7ae03ed57ae097fa5b992531213496c10902b3823c5ee3cfd75b01364e4f8d67861cd1e11d3efb305b0932b513a45a2dc03ed171637e5de9952bc4b573734ad8ce90fee6aebfcca0d4490bd31a64ae77bc16b83be2157434b7452233ce0770a0555a3f3d7e4db547a5a5e3a3e0c58552205d5db2d54ca459b7856432c52bc69280ec9e3a6c1efe3dbea19d5e692e02dd422d628fe0a331d95ae6ac675f5b202d7ae76aadd4e9b27214dcf36af66bd4c274567f86c26a20d30168245f1c2c95587f848ed54e8fd160f3ddc47613bc31ac2badb8c2cfe2a95b6a81ed59336a16835ea7a3e5589a9e270e801d1ac29a0bd5bfcf3df947c0a8841436728fab81da297c9a075fe21c54c78b2cfb45739171bfb7c296aa59fcff9cdfc524ec86d81d4010aea24c87d5752effb04b107be39f2b329ccd18f8aadd7f48bf3396d001b03d12879f99a986e13b90c9e7e33cbb96eb9ba99ee7df4091288718e58a4e87181fd22a7415b616011c314b9b42424f69911c271464283554f861aaabc05d29689f23e875fb84297b49af81317b1bbd5b559d6adcf06d1fb43074587e3aa001a383d2463d5ce79cbe878a3edd4841f80cb3df4e6a1cf517502c18a48db4832237df7d3404320e55daccdb1ef0b8d6b544dd17d68dd50a605b4a479c16744b3a24b6bc7c9ae3fb309ba024a6d5ae8fcdb16063b590a49385bd315fa0106a6d88f29f7796230f5308a79743c9b29e8a2246f8ea8939b373bc7256e5b818464a5ce067d722858e7b23c1614eb423c1969375eb2d267d52cd2fd9fbee4980899ae2a42866a7c5e4baf7b164ede9917dccb5568f2987907f76e7bafac91949b92b2130baa4316db1be73cc380a89ef4d0588647fe6f9b6aca91d73f7e416c6d05883bc076b27dbdffd39a10e40d088c54201e24ab40d0be9f9eb44946f87b4edab43bdfb89482a8770ea9a6aa10cce7f39a03b70c247557652f39e33148b6262ffcaf5f2d7294e801d69e98ce4277ee73695bde3a635a4b1e2c6c92d65216d78984ce4f9876d9abc0e9ea8ceffbeb354f38971633ab0947df9f4ca38150b888e2018b3acb57eb608ec56b714ff6c952434f72579d1f0ae88f34da14a346e545e99132871523df4c2c0593bbbdeab873687eca671c3d37ab6e55d7f0e39b97a6146415a22ae7bd62fdbd76fc0a43cc387829a03474ac3d693feb1480c2beee80fceaf7869ced93fab1c2136505bf2d0a9f1825b1c507c19b91a14f0fc103c53b3994dbf540c9be242f91cad9ac4f021db2272ae84a0fed2771485c8119ebd53c0f6ae73e258cda4ba9d6232e51eddaf62f385b05a96b8593d5580563fc04e368fb07800a4babade2e33f6a2273eb50be8a00879007960d28e3c86db4986a74e3376cedc5a4a023befee19fe8da634e53d0c17ad1d0b3a3de38fdbb013dba5fdbdb5ce5597ea9cfc582a7d4a326b7b18340cd82d94d13506af8bd10a4b18d3de23fead32e41e5ecf682080a4e0c08b8cd441b26eb4a5568b7de784707526285943f3fe80fa0634ce27c162e0b5152fa579c5b2b6fc709b058973cb7af4b00d86f1f83a3c1e3fc21700774c4dca6837a1ea10976dfcfd5603303769340fd84a5ad160282df8b88c812cfba1be43490b7d645fa00f80d639a72aa64172411eaf2be31f4ef06fa53e4759656965740099fdedc035af2a22357c2a55aea4c2ab1a3584d92cd16bcec7dbefbab6d0341f2716526548c474993a5f63d5c2b2aae3a9fef7f60e03beefa93d3a2388f43012926317cbfef34171398189dfe7c08316b15f8b0b203d5e40db27b5899c14b91a984257a000f1a43d54a93c4d6de19d68491b74e0b3ba6724ac65f78cf9700f6adbec13382ecd0eca6e237e2e8133b69a99130f7e6bd677d503151aafac2c95d78a6ff5c360e2bbbf01918db5a0c488cbc8c3c5501c723e38a6fda344058fc2d82c5020ee434afd90fd04516482ade138f706c5255b6ec506c093cb46ab0853a48b48a5ff312c30316e67047edc24698d1154209e20bca6f7377ffc521e77411c2bf5420efb7b5c3bc64cca3715f88234bdeb27c00ebaca92b444cea436e8f97a2ed9116a8459ed0a881f9a7bf58d5cab490b05c787a23ddc457697f5499b559258a40a9368739307075e825e25ab4d8f39353f508c2d79c33130b951dd53fdd60713e109df35eb3115a86a7f5ffd75275dc088106c3851ecbac3c52cff0c5a476802af65457fcd2c0d8fb6074148225c03b62ab873698a2fa8eb5b7d81c0d1f5d9719f0064c74ba5523ad1f5938cc179993950161a52854ae52c3da9cb06f3bf1f692e8b76b08bba650ebe7835f30fa56880b6e81fe491b061c64a4021bb4e4bd3352a39bbf7b181c3a3ff8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7774367dcfb688e802f64ae9b4154f7052ced6c74b69c333617a530fd0f8148fdc8b32ab690a6f0fa510fc4bc87fb4cc1f1bdf799a3c8c3c210739120ee941cea16b82170103aab39df3a48b599c908bcfd71cb079a925d9f22bb5527dcb29ceaf8608d38e10dc3307fa3599c6e8f6156167be7cefa391a24775de04ee09288cc23eb40f048746c45cc71d223616e717dc5b72eadba8f2570fdaed6dda3f7136aac1e33cfe6cb5acd1052aa13e4202e4aeef41ef56d4d729e1780bedfa1d829e41ae95b0fdabd243524b75f7ec691cdabcf43b068a8077b5d802e26460555ab93c826d227277b3284ffbf525aef14758a9a03493863f59a2d232d284b2094dd36fa40a3ed93aa490ab26901ec18c3d1ab5a2cffab0579398e814e7302cbfd20b7d700f67ed04712ae5a73bdfe8419bc377c768b913f8b12066fb7c19ea4b38c78eb9f438f8b41786734c3918570423bcffe509c038fda28928943247c35899431c95d358abe49264742ee6f4e3e5c9df74932f5a335103c8ae2ee9f6d0024c814873015549edb28b699d608dbd127c200fb78ca243a70f2487215cc0f9b5463182c61ccace716d1f4232efa0f6ebed11bc613822687f18200beecb1e03849e0895a6c03f74b2a0080931548b62c8a7af5f8b766fbce4a18e5de2b51904b93e9583e40cf4cd7616947f5209b2799dda95c1b9c43596251cc44e0aa77032717f4b7c363fff2df9ac871a00534a87a3c8de6cbd4c301649d57dbce5f18610270b10e28ffcda4c2e04939b5dc30ac47720db3da233484493b719cf932f478b6b2cfa0bfa6cb9832f3b718906e3c94d6e4ab8fe2bc33f6a8c6348769be1c4926df892338f4538314b9a942251bf9b86871ff84bfcd61ac93e5f26a7be9560fa4a2929d25ef70c62e2fbab8c048ff79f56871434806c2c4fc2693a087cc4cfe38c8e71679b8d8e7648db8a203b9f1a21ddc45cb44fa4eef19224516530d2ca77b10acd18129e9de0953189c589ac4c8978c095ed096002d25aa81162d4a7fe034cbf2afcc990402647e67f944eb5fd0e459ffce430130c7e564a129368e068a673eadbf84bc655a5187e0183ce0ba5db0e01465f7090fbdb4f190a5799763f14c9f1a2b5a130f563f93f39ca484c6180a27dfed2f24b72795db3acf9470c46e68d138b1d51ceda820f48b72eaa9a4352f9a7302803c8935f510ffd8f58675c90a9ffe67a0ff517a5c26fa03a1595e11a5efb373b1964d72b34c443a236d870d825d43a0e11f56a1236af9e0fdfc98b4e922c5aeff9f8b014545d83244cf6c1d41586c97e27a767a494ab02d8d44408613d5a684333255f8c483a8c26123a88b4eb546db6a9c02117e44a527b53f22fd7f840cbc3e0c394b441a7179f0cc8476c7e8b6c6be39e7e59d50a3b80997331219bbd08d4c9bfb3a232869d41678d0f1fc9416bb2a7987726ee89f9d350c3a7b8b0771802ca2dec27ff895ed78ecbb9bc45de32a4d880afa5520dfb920c0ef57330b31ca4b440ff69f38dff372b18e1498b80350f255d9d8af037606decb922e5b31119ff7efc803c0a34f203f8a27ca38b7b26978c1001d42490499599a88fdc8a8a38836d9860e123b02428579e64090cc17c749847bd1bd139a6c7a9bb0b5b6333cf8b2170ad7563e5231f87635a90b16e050e1cb456c870d95247a01486963faeff8631f5e0c44d785fb31adf472c50b9d01acb3e61184eaabf1c3fd1bb7fec645ddf730cc7d4b3ac266e87d0db755506d45577ef5259be76294645f0607a58698159e1c70d868a0a2d5e2d8d81be16204b7d5d3a6a1da3fdc84f13545504a44ae36c1887975acaf3771b48ba05371ab18cf820712daa218b56572e7a1b709530d62bf8e68bf29f7789c4f58d3461b9d49eb924ccb89f7a40728ddc52928f800986d7cb652a486e57ca4f364cf3abaf0e7594ab01c9fb5ca54d0b13f6c002e82d8374987170bfb6e644e8f8a328bb6a6b18f9d4b560e83d3ae6c0eba71eb8b433dd90f90155865e57ad69736649797a32cf703711961d11b214692b47f246e8254dead906ac452d4ff69558df7cd5fdde3d513363195174331bb1375b6abd0e7a6d123e8e78206c66d444dcdaf36ca076145193b8436acf5810a4ef92b0ce0e355d058c95eb75f0c55b50a0b3d467886029b875469b2b0baff530c2f0777152abda1bbadefe42bbadc356e526ca87eda8e88ae785e9061446eb9b1a11a8dee38ccad4e246e106eb4af60e9beda0ddbb692bbf75bda83f6f6f1d333a1382d6b229046448ffac6bb0fa483393c55f11124998e0f5b3078706b5734db49c71ca767e18d9403023fcb2832525ee876a981a32a6e50dcb5858fd83f414a4815cc08d6eae18d5c36c30c429351c35fe4eb1b468e768c1f6e396bba1591b597d358683fbd55731d8a80b356160ac1020f71e9426d5d5a6e61354852b0a046b5ce609a7c86f1c04d3f5df7f0e00febb09d08a2c9551a67a3fad93df64d738771b69d425aa6fdf2f24e07f43bb1f1c140c92c14130390572964413f49001602bef5a8a25d61c08f9c292de11f059433f03b49be82add8af1f0cfdd3557648268a986135fad0aa37b6e0636b9d9c13c7c75f3fabf22076e65dd59c9ec0a35c190c5d17d6bcb57c2b4ec7047b47447e72c3b8f7672c22e5ee7b73e317e203bc163400536701c4f24123e54d03ea6eab56edf1288295d0668c5b79ad819f01cdef29f60217bd93f73131661a5e3f53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3b4c85c92a013def2a3cc498074eceab3b27f02c736d6b7590e5253083d800e41a8804e6f6a4e73b5c8e4f87b4e19d9c439c4fa3f4d47cb1201213afe9018b8492d0b9a4b9df28732f02c3020977250da0670d2c9cd2798cd0dd19e42683416457f021f7b07d56fc038efbcaaacb030139c3d72fd0bd68ecd72beeb241953ba010eac9bb2a6fdc024f3686ded99a3b104dd2417384d043200bb47faf16e99ba2b8b63843a2e937d312f9275acd48b8fde5d091ab6e8cf61b0f9b2c3d1126b1aaa37ae6f2f17e054b6220e7e30a1c7e5c9c2e1e410de36277774f09fcfab830d36b275900a9de1860ffe051864a7b0be55479b3904329cee6c66a5aec510df0e1a6e960bbddbc72707534a79e81f973680ac6c24b3ffc1adb6302efa0d40388f652cfacfb0a3c74cfccad133673b315891dec8821e7b21bb70793e2b21817cf6fc9b32996e52281fa7924c8f4850f48b8fd1641bcc2241823237df6ce5f062aea10214c9edf396c6648fa25c2d7b7097a83f99457a64e99ca006efcc0162720947bc507aecc42394b10bbbd8b989235edcfe5e2cf309465afe43e126fc05b4a683010e2a37958dddfde56a7a896e38da1989b5e75bdcfed6ec58103ae382d2529ee6fb61ae8ffc180c303b44a0d49ab6a2e5463b20b3d6178408349af3713ec1c2f82d47992e93cf3308a0ea6eda911b15f004ec29c3be4169c13e5cd619292e955f484e2e720abf31180744a1a2e9a424293fd91a4ba635fe545c2206bac81ba397107c9161a89aab316782c142ef63896ce34774b3ce04d064dc88b5680cad43bcf3ec020c41504f38346543e95ca6e13af7fdf76d467ea0fe934456c0814e59d6b213d833c5b88486736cbef821fb9ff4e7be39e806b19ded7a44c2ecbd52720d0e52c44d9c75e03c29a172d3fad238bc15b1a17e27e93c84aacb5a2e9f626c4976c5e2400981aae46dc6fca524193021f1d926fbd0abdbee998d1bb0245368571095f5f1d49227d5d725ffbd7e668d30fb47ee55dc0ef3a238de120b4096448d18ae1e3853ba4d778b64366532ef50e802d86ec921b59d79460b943b440dbddad5530c23d636aac80cf02fe1ab00f7c48ed668e571160b3efa2bed647bf53b5584025143b9431031d56a793a8ede5664bc447768ea77639f2001819a8510e066787db59e78bb2dbda9915218839ee347de3c98467bd41c86887a8d80beccac7ca210f1ed12af9d99f41fbec25562c6d9bea613e9bd5ca1cca00933233deecb22ea6594350af9e7b2caeb2576eb0289c64fd17d576cb28b3fb81ead7714150862b957b850545e52724ce3213eedd1042012d4c023d97ae01f3e6d179fc70952a64fe89960864a7d46260827302493bda1c4634882ae07262309e922856dd694b5986bc502baab230cfe3c1b2ea976c4218f56b0a18f2ae0d46b0b1f706781d1c317669483ab167bb976623b1c573b725c277e90e78a9391638f89e00271bd7f367338441599058a6c24ec452c6c75d86cb07a220b5c19fbc5a4fc7829827bbd99d6e2cda52f8e59e0fdd3288159b78b2b44ec3507dceda8de6f2f2d589e4b593f2887391d79b3f6c87086f07858f1b479b9d720da8048f9f358b9934ea172a08695c9215af79ad7b0745f90b112ac17f6c23c4ea924205d1db68726c92997ca94da5af2b28468e7668da316c4a0b2ddb2fa49257d0598c2f1530f5e35cfe4a87cedd675fd3de5d6494758bfd3e971b9820def66c17f716012c1aa2ef12f0b14d753bc4eb4d5e338fd6cbd12c93b987073e19ac5b0e9982edc986010e95c3ab4e607e48deb89265917b1f4235bacbb136b21e05c956bc54609d9651f1f35a73eb80115a0524d6da1b23cf26a6bf1d4d6c90475628ca1588fd44e8300bcbe159bece4a250072231171e954e3afff7d181e3e6bdbc7f69141ba9e894478b98295ee047a6aa404a842979c03f2d80a8d6c6967bba55d7a0a4eb8186c7ea5d8b2eb087eb9bb01b5400e11113363516b12366a94f6bfd2a2f548cda9d4b98ca3606f8cedb8cf06f0e887e18abaff96dceccf50a27be3dfba6e35320e0efcfe03c18207ff601ae0b1f9f34236ddf896b3234423c9b769712fe124005f4237f1e0920dd60fcc75ab26841dc81231a865c8b1376d9cb508e42b0aa41ebbe526aefedc33ff3cd447893045071e20f80120d7c24b89745bccb01d1383799d673a00a357b4d3550e455259afbf7ff6f735f6a6f3b88e4a8795905f75c1931437fbf13918302a222ae9a1de9b992ff4b3994ceba4c01c01e137507518cb05a135765fc7eeba1c3e087ce006e0979ae4a9c30a59d91d5bf8c73349d624385cd368d1d3c4aa6b8ed719ab128f89cb3f401d7603d2574d616b3d46cc3830f3ff2784594677d5b255d9ff6bf90e16934afdf38928a844959be56399b57f673a2e0c72f001be3e5fca88b815d643e8f7aa02d06b7f1cccef81c2628b01a5ef036dfd525e77ae6874ffcd02bae95c733ce41c8581c274c7a2d0095ed162302df1e222a69186f89f970f578da904708eca4854d61fd3028a070ad6093e2c4f616f08ad438c9c4084ec1efcb4accee3b241ec83ba4539189d8a349e78ed52b7d6f035a56fb33cffc438d6548eabbf4862466e8021c2d94739f40a61560b9e2ea363c6705a22bc73378c068ba84b9357c631071c2116df3a6bb7a3c6c0745a2b442fc176bf045389b3489b0c48b65edf4ba424af9788dc6f49b4d0fb1dc12a95aa06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6f64897aa45a1cae2b72c29dd871ec7dd44178fa92d9aa77c294f375cbc9296c1e89aa420fc84ee9ef9e888bf328c124ece00b8eedc3fdc13073e2d932c4b31e8104a164ca8c0248e668281721dedfa2ecc11825b838da8c26af0e06f3a379c1ea229902493dbe88bad43c7fdfcb4e723108821dd437c959799091ba906b00efab743efd11fcf0ab7825f272ce1be1cd5b07bdcc0eabdc5f695feefb2f520794210ceea4ad5041f9bfca6546fb6f10febd750bcbd66a5432482676fbd6db908db518e8addae662edbf8bd2477361d158adc0797ef788786f557f7fb4bd8307fbea4c90262e70cde2a17c749373938cc8cb9f61f05b869bcac55f6ed7fed9ac34ee5470b659e884149c5a0b84d3c1e4dd63ee6876d6196730bfff11e392359b81fb1387a0dc0557be27f963dae9f8ac8c6884f9234a265bd7059753b88541ac2c8ea640627573953fa511a9609b9e6d121d769591fd43fd5b4a410a646c2349db3fa4eb9718640ff0bb5305c86c2b47176c074203b2f8204a97192195909cb8ac9996e950d5edad4dab1b51c3e130e60e94c1c8ca823286f00a17ae7d7c94e201b892f6013c86503238f1990cbf10f4f2b6d16d490b1da95c8bed8e5d953021c56f57c73f744080b49ab0603cd883fb1aab110695b8a32abf32215a5236ce63ddae44b49621817574841b37dcb3eeaa68505f6d5951dda370522d2e80f1c5749222a84d05f4387343be78c3b6d655d513a3f7877308145a1dafcb72cb53ffd6c5fda18cb1d8f9310ab5f82848eb58e2abe0b2a1195c28753cee8eec08a417f5b32c2861aa50e1bc4fbef5263c94561a8764b6f9e3d28037057cbb9f98b61136e16528b83205f0b11a6e13f93b6d2d5507d728e32c4661466409216a76519133b669a366b6414928f1b9ec67f7a7cb0191ad003810f4878498aa3e023a8cba8d3d9c261cb3c99ca41d3555acb40cef715c0d8ca1d372423600d189fb5d5f388f7ed846e7c04fa253c277fee5a0701035f71b624e0caae48f95c8c2d232b8de1fba7ff002401c80833bf666e87a3946f7ebe9641c1358c1e463205445b4f92a55d84fdc04957b9ed94e3a06206b3adc7b8ed1d8e5fd43c8c957dab43e2722e0ac4a37c369101f1cb1dd61663eed9934780ea276b74ef574e4eb558d7f17743355891b25abbdeeb426a1c538223413250ec95091dbfb195ff251048818803c031fc74ba9c9e21e7f5b0a77a6174ca2705028524695fe7dd783ba27338713dbff96fce60b86cc07416272ac5ed62d94f37615116babbdba41d4e5d5152f34729f28af8490236d248c6a7fe521c5251eb21e95d322cf405df83448c4327ec7e3372da82971114b247de48cc734051853602f0efb59425ec5af860f2b142e35ea65e2dd49d119a399d7612db75182f75074851b5af69c0772fe5ac64dfda0c97e1580e601936c0cda76ffd0e9870193f2f1fae12298f07f59cbfc7605f38b743c974fe2963926524153478dd73c71f48071a773b27a25482e76b7ad5713d2ef0277e915275d2deac0183849100604971c7f1bde78aa6fd50fad2f89b0d802469f54be017acba308c2a825ef8b0c2fc36a41e08124573fd969443c0c048343c1cb19d0a2619fc43f788c628863bfabc5e929ee598897c05d82c4bf13a876ff776b5cd1f0854eee86788d3e0de0f0f5829f5798599f3cd955afde4ee2fa9a04db9c62d3b851b3871e89f746f961c64869de7194207497a7e9d9ecbdd8d78fa1c4adc5f5b7c22ad3feda1bb0ab698ab9813a6d9b0c4fae1527f866a4305acf91dea1461dd4a07bb3d9f343ab0924050ecc4a071b8c66d1cf9994dd610fd715dfb247fa13e25e83c7452fe8885d2b972d7d5a0b65e6fd14fccd2324d1b46d6db65056a361cc94b4f38a7d98f54fd531d232af04f0d740cb7eca0e861b01d8b606352b0c0d24669f6d249512526ed97fda96aac2a10c1abb8707113387756ff896475e0855c05baafd7e9c98f2ec88219284da13548cfd6a65d9331b5b1d47bfe19fc281dd6f7800ce419bc58ea94d3162f1c82d1d3782e9a9bf4cfe3258486d6b98afb19a6eec05a515a03202eb648678bc691227632fe82ca8a67ff839cecaf7dd52e4173dec7d62084f9985333fe21d954fa9e89fcfcc0c769e99f1cc25b6f2638d561b35c40d87a6e457fe29a87458e3e88d294a7551c79c4d17a495c0333db074b426589379a75ba925062dd39629b13fd1ba4dd0e70ed70c7cbd29cc48d51687d3c2bb1ea7fff074a2126ad11eb40df1da7dab2b24c093baa6abe4be99d7c4522768ac6dd189b8f1c7ab43efe5ebf3d171be41049c871984542c78aa4ea586c79d5639d64775cba4e26b6b4c12ea51c26a5ea5d858deb69d5c94ca04e403b8865117efc9c45dc04d3e0835e042f0be514927f922b4ce7109a484d12fad3252436179681e1aa36ebd0a4e0722be57fec257e5d42f59f3f2b97cde26e75ce2a900bf620e0464bf970790257ac8e02a719b921c77bf723ef1a9e807c5addb1cbd82e5061284917052a5b3009a5ff0b2d5f2fde64212c8aa04cd1e8a7334a366bda35f355c01fd576eb858ddd168f304fcc8490ca0fb89e891f89dd9b070c46b35ac804ba5d68c91e2fb120d56306fa64da2b1b2c0277986272a1b83cc482099f588ec304436d49fcf955e05aa819be2e49d4539429290f5d068c45fdf0de86ac36672ebae56c3ad0b86345bd561769cb91e9007cdf3f7952d7d69b585;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he4a63507bb269b72a17bfe392106cc8c31156d1885982ea541734a1dd8084be329c94e9dd636439cf47857010d7418908d496556e64aed1d5a10a153a2e2c97e40e1dea1fd2e01f695888cbae999b14a51cedabfff5c92b4ba5147113b9a9588b9841ad923a334a6a4fff2ea00413e2cabf8121e2d61209ff6f10da21d22cd714c20e55254d1a19479362497bc4ec0eadd3cc55802bc612825768fabda71c5b15f2645515efb362f823a179c2ace1557ee31951300dd06380a5533bcb53f7289558c295cf68c419d7156617960953b3f028f12bc5fad98f3829daf5ca4727612c4f73dfabccc2e34ddf87d8b36739dc32c942814bb2bfe9f59d94a93b0c15589e47993c7cb5efa5d86ab5131ba92d8eb51e7d08a4d6fd3799a7610b043b3cfe3b6fbe5ed53559deffa1a456a921c0e4564a71c73714abd80857ec620883b3672571a04f002b80f99f39aeaf68699067c153ebf64a0fd50ad636fb3cb73b8bc1034938eef6b20c6bee11608f585f499a62ea0dbb2ccfdbad32df8ca47f5c492dc18d3170bd33819f32e48e8815c71f4994ea3ef439f29693c99877ebb51b2cc602aa189d928c19ae1afca050bb329363baec2c2b09663c4dc429a7abe460caaf42ea5287e61336cd8e13d8143f8171af78ef6740ccf226ee51e7b8dabe613ed73fa28fa19a059796620aa2015192e09baad2ecb3e05979b5be5dab24d28ba8462bfb5a1baf9c309f76ec2b8d6f76d3d69e8285048a248deb9cc20ce3a5e500bb3d66ddc0a99868a61839b1f2b026a75219afe923e3a2342c6de34c3cfdf6f653f13ba98a9fad59ae1215bc41202cbdf413cb952b7c3ea9f744a3fbafc7d1779b42db90643b95c39649702ad34f20a203318fe4b10b6c49ca2ab7181a780ea4d592fdd797de445046ac38f1bd0398542ca021fa97b4c64c9e0d88ba6b67b9d199965650ff53cb3356b9fadcffe8e8e987ad7866fecee3ef6218ffb7027a0570bf026fd60df953ba1b6fd9a3df709526be90a842bb83c92633c38f99dd29e5a0cdfea824f2102aad868ab392035f1da3497d585a8f245c92ec7adc728965df89745efeeb1e6b2e91be5d1980df0fba634ac7f1b2f0cd7b31c6297009f7243bc669a3029d3a770528a5e674d85bde1590d895e9cca88f73acbf7ac127b866688b1da2625ddcd117f9a4e91888c6dbac65d2cc3ba1042c166c5cc3adec7f9b43db26ecce7152323f8b6026affd8065dee511b6c23e3155d752a9ea7e37f48a8314c67db85a008a438aa059e318d42ab7aab5c5bc0b898335540e0a61a697c22f3483b71d92f2ed4ec4c6f48ccac0936ff5400d5ae7fc84f28bd55d53e80820544d3fbb92bb257c807bd4490f131085151d67195288f0d6f5c4e907a8bf6e14e845ad76349634fdc0932511bb1afa24dbaac390865aac6f1b57737fce178bcd57c5017563b7b9cc3d6ccb85281ad50bdcda874f873dd01fa0359a3fdf050763a71549a8abca7293bd5025c64f38a493406b6782af203b8c0b59b999d37a5d982b84a125511dd941c5393f57b66cdd032d4861d852feef10922981c7967f8575cead3c933a14e192485e84a3109020566c6930e219b22f5570170c00711c747cbbfec92e9d4cfb2e1f9405ee1e52f392d382be7cebca4a87fad512a6c4af2bca81af5dc3b0d1af3dc307c52868e8ee7a5d9bfd67d930c91b5c203a1e51b43cddc2755354a8b9dbaf440be3e8cdbaee93c6b66e15b38b2f3a07d27547619fe4f82eca3e711dda342d0ae98dd41b74052d9eaeedf92e0219fdac7341c2e05728ec7d66fdc686586c649646218040334a9ed1cce55716355cb0cfb275b71b69f3409b0e343b10febe72dfbf1c8f727c37e75d1a30782a102705d7d368c0571a68f31dbae7b17156633fcbbae073d054914a522dab4fdd369053f70dcc899d3decc58ccfd1678d95c67d5d80b18f1635fde12ecbb559a56b74ae69ff0e1eb73e34384e37c2866c1778c738952dd7b08212d330ba3325e490af0ad8f5391cc2c89cee675f7fd2fd5afc6eede98999c7e7ab51fd6513a33d9951166fad6f144f7faa68356f16b8728367c155efa2d024dbed43c96f4768d0729bef848619f0052d3e6a823ddf7a555a0b5c6ce20f04ca29debbc5f0d5ff4f7c9d28c3d3aeeee653ca8c80992116d6358532925464e2fb0bf9591e56459144aa1fe3927fb6ce72a1eee02c7f280720691b26159a8bc69244f67e750ba41e5e9907fd14d2503ccab342dfa5e88fca68ae91d5d5a721516692dd5f55d788d4310ab23799f15c709b631928d7ded696f8cc7e6692f33519fcf8271d37cdd7d6c188921811af81b754af07527c45634332c482bd62afe96551f443b4c3e68207bc3f4f5c0782b0d6432f3fb9b0ec284f9060631e053e1aa7c74ca5a3b2ab3f416bcceb13ca03d797c33d79196c0a6aae0c3ea594ccd5fbdca67c0d2dc9259e1262ee48feead7580f5a7b363bb6786e196d4a8b56b24d91b0561af980cb535fd3a637f484f69fd6c297ffd3bc364e545eb04f82f918096e893b530e8473a0a0e3af44d9a539c4bb75afc98ead318ea2564fb3c78ba56926e35ec20f4f96b12412d89abcc143acebaaba504050c81dbe3efde143bfbb2d0d6490fa02b97cda5ec35ce5c1c129121e603aa42355eede37e3b68a828e9343b40d8ad7b6d5a4ebf1cb4005384d9e69bc8a97bb1b492508466583527f6284fa6490d3106fec7190a1f6fd8bdc0ad5a1c45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h456c598761cb8c3a430a803431392e7640c9056f6f02861a34dfb4f692852e4b3f78f8734c4c43f3ed5b2a29ccd4054a6d6aa66a9dc12e19e268556eecdc09c04f48661d3649ac5caebf5b0e9f77d786c8cd43174214f3e83e9f53e14c3cdfc9e515d53ac882247edfb588d157fbe494a9f1ba643ed7b5bf0557a3791185648ab9c67dbf41cbaf76502eb878fd3b901b1c631ed5218980cb44d5325087651fd6fd1016e855d741e17c3a2e7a64c10c608c5d60062275b097a658e31bbb15a1dcee4266e22f07ffbb9f81e7d3c6bfad4e3f19783a60aaf103d85815078903f32849c2070065a9b0fedc81a17cd5a306c028b0f9e792e6da9513693ea35ff5184da5fe42d000874b69ff2f6395a0fae0350fbb7c930d555143973c41904090556e1015f4ec6218d121004fe652818e8ab59e938da9c9a01b47133f0ac2c40f50339d534ae065ed4ec37fd6f961b3feae24668d2109b24f5a615e93f0be24ddba38cf817d63c0f92c6637e70fe2ad645c2bd8da176316af78864030645562a461ceee220b865ce294569644087da08f4fe123fc1236a81c842e3b3d594520c3986e9d62d8eb5eee68afac86094ec0d62d89b82dd1a434d5fa6e70595d26b0c72ff9a0d90d240a5923ddbae1dd826abb4ef22a295356f4326f1ba6e371f120fbc7966871c1751be74f501f93633715857641ff0c179827d77d9fe344889cb9794cf1c9ffeb11d270ab34758be3581500c4fb8f07fd47770a6d1c29252045f0f7a8e0351f4caa12f753d80755123aadb8d22a1412bc583256dca1f53aed0322ec9b9fc95cd0ec548f47f5a2adc6e9b44e7739857a5d5c0240541c8b3e0f8d3c4d943bfd57db09942b851390b29622891f026271ab261afb5d870317a1d39c412b96a886542ce5af36a4d88e0bd63ba3fff0ec26b817e2d347fbc5e92a04508474621952b3701f24ba09c8a468f35e1d1d3869c0c06eb77687c6966bf1991785188d64002fd4160812d28e97241e26faa3f0b9278c77044fd058faed3fb7c514d06f011806c476ec1c1a2212ed555105f03e48fd6366cf71800b2fefbd3c22d66a41b37d50c6f04ccfcdcb8392c1bca08abc3fcf54e5f17eed3d1924854fcaf8cc8f7b3ed34e3fbda489c764ab7c847a67914524092a4730179599468285399f7a82d3824709e38ef00f1388746fafd8332d0071dcc18c886ed40c20f55f94b68f6b298ad3c2eb67124005b7737fd16e0e0c33b9d0c711a255716c2f46e238065e0990ad2d07fab9e4dd157fb0c71de58077eaad5481384dea049ed3ff4a7e77bb86a1ad413161b4c2889338e8645c1fa7084601c1d0e1c2ebe8bcd480f5d8ff6e983d251b0f0292a47ab9f351d642e2f07dca700af7f5a281937ade76b3a3a57f766338ab0335b0cefc1233c8e780064b9724237808619536cd6c5ca448c83158cfd3d2af2c56f2484244ed50e364578205b3e79e942e80c62e849ce475fa83bf0faec6cb63b5de83ea54e00569515efe9fa2e34f7f93c3f9d0f1dec9f02bcd657fdc72df686c195b2928d6f8ee52b40362155f0f677ced455d755bf13d8a247bb1fbaf5abbeeeb1a9a05df2f4c337edbbd1446015e98d2243e0feeaa3224a84987ea85b3e84860e2ed8dde92db413d915764dccc6a10ad26107bbe8333a5aeabc65c929a2e0b6034618fc5c8f6e969dec062a7e8e69d8b027cc54c371e5816f904c8df1ac5ca0165959161bd08cad0867d13ed129d0a8d0481924c5ac82357829286dc546696e72a66de4b5e724e2797a20d8bd4121ad0bf3cebfc660fb3bb14eb820ef87ecc852ca4bb46cb95032697fe6a20ee623fcbfd002e9fdb6b75b3ed4eb8825762a5b8acc408f1beb0856f4a1df5d8063542d65cdcdf77417c46658d01b86611d9dde0fa593a564d7f95c762f8c276ffd5b90838fd7b4639e573fc9ae5ba0ae4bcde4c5863f44f905d99494b13a5be3b82826784c7b6cf7ab552ea4c2dda76af7625abd9934d5faa3f90434b7f5d9c7ba3ae0cb6a4e96a653aad19c0577c51adf915f68c08bf655020a2d091f5a31a6169d8972004251f0f5f682add6eaa42aca7b6db7a27f25b819e83859dcb2fb00f2ece1ae5df6f9850a2ab4e296cd86515c927deb3d574f142d6b3317cda8ba30a363a23f0d20c03384a55756563a73c7d45828502a073916a7026e372dcddfdae1cf39b131034ab3ce37fbf59083a3f9b06d0e002b43c6895c6dd5ee3578dde06a8f9b747635c4c0cb257589da50bd7d2be153f751c9d6a3a95c6e04c6b9eabfa8ebe5a4ca984a1f04e9acdc74adcd0cad14fe0efb7da9d245def4b1aeb95326b5ccbb62ad458f1f5a1176923b13c5741a3fe310f7db8ecad3c58d0db833cedd8ba3c109a7ab2dfa48e949c1174b27e122922e252291e0f0165d53982f27aac92f264537c76bb65d46ad4308920944f8b9c20fe0d2c45e05985032ab01955771d41b77cde1a851907e780830c5d74d6bb7fe6589e5c065f15e78e2c85dcd4190dcaa0f5e21abc7b8edf5bbe70d57f95393a303c5879fc0bced10e9f8ab22d5059505a8ea39dcfaf13132c8bdb1c0bd138515a806e2e2432cd7c4959a435c2b3c87754a5080a50ceacd69a4e9e7590dfeb307d6e6ad923850f5b5ae296bdc5870fa8fec70ea2c23c3fc83c2a8d202c5f23f85d00352c15d27caff740217a11e0d885ff5359f9afaefc80ccf714f5e17547c611822a21011d87d1a45c6bb1cd4d936167b9b2c041;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc5e2b7bad20149c11d63ae9ee18a4f13fba5412ab56c6f621fa0e33a4c231952b5ce485e514963b03be8505f744b1c249bfc182db0d216883b34154b0a02673497f9cef77a04ee5915de95e813fcba14a5b454237a3a9cc68eaff8780f278c6e9724dc748b6a1aa8cd084f066d1d779cb179439a22d227d0c49cc9df91ae2a981f8813e98b65404af0dc725b5f7b81dcc04dac3e8906aaf75100c90f2486f9d5c0209d2a3fe4f2b1e5ec17e7053dd98bfca60f3ae519ef8fa47959025d69a36e11c6b75d3d714a60fd8c46b156d0a1ba3b904a47299dd3b33798d810b9bf4a4dd21a669797700afa791536fdba3f0a4a590541628290eef7b43444f7d09c08e57b23e4ab14b61094b2d060d54d507c59f48a1c07e9e83d186bacf164c15d4e7758f4b5b7ed0c6a090287a57c212c8050b217adba8cdf5e808065a39ec615b02800cefc7f72a5c3ca697f04814279bba94989338909498264cddff51fb4de1f5b8d20a6569234a26d2d52e14229183fabafef2352f075caae0edcbd0d0d4d01b0f26e1e2ffbd80b1ba7681b28db6dba4acc8409f918b683990eb860d81053d3744677dc4553f6b38b42c8201ef0912a07d0792274c51455e6396afae63603f4a70293139796fa06fe6a623bac23b9f491c89ed07162adc1f1f845aa1fcfebdb097addfa2dd9cbebdb771d3fd17503a1e9acab6560781be0bfaafa6f130878b1ed3af6e062099aeea4e87791a15841c47f0301d8d28d44a12494cb26d685570ce121e731d51081783f96000f403574680a470c92e8d3dc049bfce4822f5be5786ed93ad0db74bebaf0fc7185fc2cacd95a8a6b28493e18f20a1ae4557553cdd34aef7224059bbbb0544c106dfbede35eb9446dc0246b1a1227726ab53ac4f774cf19b0e0ea3695994910907fe2e51a04f5f34a58cdf09a1bb2238e01ba0cca6713b467658fc73a484fe17533f489bfefc4e02a6a0f8d71619125b325d1b07ba5196b4c05114f298b8cc79cdd1bbcd8ad73b0d2c736fdbe3ba8c8c51ee394b0d626bd25250cb786ceae9a309ac0f42c4885fced2d8d148788811bce99bd71d80817f49a32293637055ee681bf40df394d5ef30c310349942e6d5ef420e33dd24b8feb2fe190f089e83495ffa89ec391acd5242e88f78369a75733e59c0573f6d9c6759bc9faebd9f393562ce950dd44d723ca12e77eb2b921a75705ac0025735d3957eed18074ef7fbcb8c47f07ec846b58ab48ccd282b3756f5e58856590d329068148113b4e6bc97d79684771b3dc5383b6fb820dc8379eb5bcf2a0a62f94a8c1d565c733c20b587fd0ebebbb75a3d0918a741cddc6535dd9a9be0eccd09b347562d3294e66fe9151270ee9e3d578ec304332c1115266dc81a075faeda67800a1db1cc82c5b4a3b3bc9fd9360e8089907fe4625292399c23ec093417fd4b1918769c6979f4058262ac81a893efa2d94193f5681fc6fd329ba8421b454f7568f7b00aa08c771278d7a11ff7f53ac059c2442b270682582b682afc2307cd78cf60ae6aa8b64c134a69460916103fabf04311cf9ee994a9abb012b27ec5d34d6a09d849b57dcfe6f38cb1d027136e32eba4152063d920b600eccd350aa160509e13a709e6ba52c0ed94c264de8bceb2df5e4aea2918f97f36783a16b20f0ba003a0ec0749eb1dd6192dbb15161b2291161f7201746d80c4c39ded121a59c33a7bfeb030523bd9ab893f4e125ef68c64a083194095388b147bac97a55073308d5fb65e755495fede6d1a59fbde509bf07e58e90605707230b47a59fb215c4d0e985ac3c398b4fbf992e5cda6b881e4d4f45f631e6f6cc7a4f00d259c281bf62e71b20bc384739976bcf994a3def9c9a737966f02d653cdab00382d72389997134f755640ad4ccf82b506085233af1fa19cefa093d615fd4f83d33644903b664d823b6b69ca8adc4b207db9fc93aca34b2adc1891f204c468353aeec896e2bd671a83bfcdfcb940567a81cab3d7edcdd5a514a495c6d6fa1617f4c5c16716d23a9f611a3d97b4430247d28f3d6b64370eb5e72aae39c983de8e405d8fa91a3e07e0eab50f84b09e05b4d3b4e53b83165a46ea913fbe380f648468e5b113d6461e2246e4779c8919b4a10591b68bed660877f23afc85f9b9e5de3131aa61a2136d64f922dd087c52eb80d4cb46de3927ac9216b68edd29679bf97ed2dc5abc1f74292f5a6980070eb0ac071c36c5c88065b31066990d90102828a1bafb55b16174a1570d8bf314bdca6ce07f153af60c88190aab5b40ae804180cbf9c8108914bce2d0f8f5292713e061386cac407919f074fbdf49335da8146874cc1b6efc4e2091e360cc2d6f1c7d1083bab66bf594eb264f272034982c784c9f4b8457e52c8489bfa818038cc1b31e4d9eeed32a4bd94f51b54fa65e3b482144282d69c89d9aa5215b25aa9e1d5e442bb4f3c9eba1a0561a79f95ee71e9ebdcdf6993f264053b967b591c41a57721c64f28452590c35a20ea8945d0cb2b408612f7da9b88a3e120a0cfee9193c8f0e89c85bd9092247e4600df20b2a15620f8917fcdc1849ed96fa5b48ec82d0e18fdc0f2f708d7a09931cba6a0d58a32592fe69ec8da26ccda9d504df133135e44a9e47a4620a20d29c201f4bca5e4cc7dbe8ed2cbb3b6ce01d121220f44aadf0811f6713a62c754154be007a0d511f6427ef85511e401c2b28a910233b865370374432a2c44d62b539b684a69baf173567591;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd43e7a5673ce8626bc260509b19a1cc0fb846775122c2a12af55dd664b40572c676615411e878d78fabac8d8eae38c143a40a20e4f9bea920445bbb5a6c6b7b7e5b8d445636c410557013aca1841d5ef78589e55151bec4ad159204a9448a74b42b8d4db85c653b054d7285f90232b013ce503ed7433afbe4386ce7491760b42b50bda6314a4f20188132d8006f3bf1453ba45c536605ccd1ccd8a58927954abf6e4024905d3784b00804455dbd31cff51b2f6196cae899ec5173aca7f66be5185a3136b49e9101d0dd982393ad63b3dabdc8876c6ded7e90812b79177b69e61ec96e48352f8ad4e5e287dbb668266c973e6c95e693eeb2b3bc2193c56c7cd286c5fd6f838f7f8788398280f2fd53011bfefc06216bf19a4819786d685388b00ded193f9b343feb6eed148f7259b803d918d6a28372705c1287d3f783817bfd6993fa65f2cb9da46ceb853565b42d178e3fc7cb19fea850b8f5eb3f3f4ea2d0b5e7e0b75e2c879c489f179b05470da690f1780cb10fac0269dc816e93c1ee53b1919e0720159112094f708f316b4099895154accaa1a5a60d1b804b0f871fe7b12e1a60704629e44c094b52189ee1de37107717dd9a56f2933b860308938451a1f43609bd635b00573750a819a20b2d3e5626246bfe5d8d0612cb9332a6b009ec9040ff17bbd41343a9b447673e3a3072d53eb68ddc537d50e87ef1d1ea48b10bbd31b4f4c2b534fdf678b7ab640393bd10e6273358d3223f0ad8fca512962674aadf3ed7e1762f9fc81ac5b3992983070cc6f4f02fa3936f1e1a2094f7ac88e7a90e939db03405a362db2ef7d5555184eee2b36f680907adf8e078d605ecca873aa9b7f7a5a861b44c8db601272f680ccef798d6bfb8094ffb7e79db44eb733ad0490b8f82c5e5d73283c0f4246eead9b15aa88d01e2d8352ebf9eb29fc842d5ef411b8f7c1ae74731038a7e2ff487a7e8d4e53609c3c0fb259b1ca970e28aeb4ff66271cfee78e07e93db213a1de7349baefe600f3dfbab8ae4a62c47284d9c60f993b7d29012f296b472828385d665158432ae07e9be8e7f2f5c6dca42951b8be076b7b1846394cd9653b3be18e586c9415c28f638ace2befbd132c2e69ea2a78b7f75ae751794affe54d00d4c3a7e7bb5404dbd84637987364ade7d28b96a64a14db57eace705313564b37e052c91fe57cd3ffef733d1eaebfe722e2c869c24bb56ce3e4415b94548e634dc85eae50e4db05594152ba3108fb254f7bb7a9590640fc433e2d277036290c9245d9653c6985c3463489bedd3364cf585a4814da077d42013f40ad501b79a729f254df2765b2addce0215974870ccb053c8639b3b44650d5ff9203a2e2ded80ae418b155235cb2589f9ab79a25b8b00a0653790f337e662c9a897c134d26cecaf2726c4042b340b32fdaabe1f643d05d657889f6874c658dcd81c4facd6550fbe25c57fbb4b3b1539f3ccd5d370cc48ba2843dabefbfbb8f2e5531e630891a35f1a439ee91871a194ec1f5b87676f0574c7432fce4a1bfe328739e2f05c359e59dff29d3d6f7e373876c452b862679a2c52876c1d0b27a3f129f7cbb8aa169ca6421eedff431b9bfb3a5282905a8cd87164ee8d38891ada7b778e41c32cd970b81c5c26622ad2d3e53a7a93ca6935291c61cd5e86c84c6f5658928a80a9bcd84c81b14763d336702bda33e969cda62ad0d03810a1c9f02b1cf946f59aa7d2e86e279126be46c138f347fcd51f9af166152e3f2552b52716daf4fe525924cb6a65358c9c884e734313dd444298900ca8fbc7cf5e4c63bcfacfd0d911b365684d5ee19b4f292201ad1382a6511c7b0fa54574a04f8f9ee67a79166d633138f3b36e0e84a3e1e9d063940cde0f1fefe81ee70f9a12f766570e665fa3f4028f6a5ebafdfc35fd8052c291919a720f32048b3124d08cfde86d6be646c0f2c1f289b0532404f1b601731d883dfd308ee7303487c87884c4c14a07883ef6b98450d6485c152d3797b0d74f6de83b6e45b9824fbbe8645ac33593947eb7f50a7f29f2b9ea56a539a5574ea55063b88f13fd4b18394c6d1f03a806dc96fa7352dfcf4d8fd072c8d6762f8d4d0cdc92a6f52a5371d005c84d870a4ed2f500455bf3fdcfefd9d91ffd69eafccf369f05eaa0cf96a7f0b3a525d465dca648a437c677aac800ddc0ce495e0d9a907ede21be0a87ebcfbc5e228ff352e1e61aa91845b6a6a61737a83c140150c1e83a487f03353b10984e8e3e169f8356513db695bf8116d6a34852ce8d69b33f0ce6915c825e8e4847e7531f7629f4d300f58116ff672ae85762e7c6f64dff401fd0d6730e4cf478325c7eab1dfb1f28983656a984715ae6469dc4d2cb80efdd9ee4ef8f1a44569978fbaa186a152563989eff3e3587f0ab2e3a3d96dcf65c95c6ad019581185af0ab4be56077fadcee5e33ad4d23dbaa484cdd111241d49ca37799cc4afc77955de2fb0bc32e7912610113c989ed1037ca1aab25e3abbbce69388cd24316d85351287394f50325882a5906108d6cc37aaf9e952c2d3b121522f52cdb7cd6e529d34b5989d0bb051e0470cf13c2e235dd5d52546e3e7df6355b46a832851a7d5f78b982c921d204ffdf2b48fbf9da7e10e12900ce62d5f49f53de95ea71d8e1e426734a36fce71c92a0a083a54e90a0081d0ea17b861b44c5479f4846958ec19ecf6ed9369d98551490c347bdaa2600c579b07fcb75b99313ecd28b39986;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf8a89a9690e71ff7d5c5f5c93d51fc6c3ac6a5924c3c459df73fc7eb76664425889c7b4ade86b364c269e60e7263698fe5c71bbdb5f9f8ab5d3f209250ca891cdf2912cda4eceade1511bfc5bb77bed6ab1c1d42ee2885de26b973dac79e9eaf4ef3ee22238051e091f1fd8c0f5ef810ff3a4d8bfe865e25686bf3645bc1f08940f7f83d6c93567267f09e149f59fa137cd08ec771fff9fb80796abf0c107a76decb53662f92388684967738138f1067cacc156e61df00e8c3ccceff34e744bafa76c47c4ca7f36b3ec73caf2c5311bb040cf0ebfa5b291cd533f6f46f8d8b538aa16f77c188d8c54aeb1645487c46e64ce08effaa0e6463352790c37bb56e5e91a749495879ceddda463e36908d839bca96e2a55b56139083c7afb26b542e3345228ab1ca5c9fd09867a2c551daa1db61693c6242c6429430ca898969c1d9e792b5f0d80eda1cda9a157a115f11bbd5bc60a2c1acd9add2a0786bd421dee3e3b6faf5af336033795a785991ae2b7c5857da0f8cbf5b9d085e69d4f667e18fb4595263370908ff6ae43261a85e0eca444d33f799d0af9f3bde9e3f0698e475c4f7351243787edc5b91585e6ce491dada01c30cecfa23c0fef7efe41c5269b5e083616a657beaaf7267d3bfe7d1f2025d4624a2de296d0d09791a4eff787ddb565a786856c86f7e6a7acadee9ee4408e64565cc38ac1cc3685d0ff746780ab86711e97fe55716a9e66fc6f8100a46c591a340991b93c19c8a8dc86a0ffaaa21e174bb87f83ecd462330fefe686410bb017ea6b365bc8cf9a512ce8ceee247ca49430fe2fbfdec348764e511c7a087d3aafbf7467ddf2acfc57855caaa7f2b0fb6e5e8d95725f25c2edb3e3529e720acaa558dfc1ac9bc376134f4635ce92a3e49a436528efd12a2f05c2da0277bebeacd807f8cde8e32138447414e2ac7b6a92aaa794f639e5253accd2d83b0d65f361113b4012ba531f2fed710c7415375dcd3f03f11a44d0e2b38e6d7413ed782a5ef9715c57e2165e8ee00103730a0383213b725fe45972a33ab1255cfe0d7eb4a94a452a8445c29313dd555847b2398489877de64a21b864c540cf9ee63a66680472d5cbe93f5cb6ea274ee32391fd467dfb87547f114c0c373455efa652ea1e3bcd716f694a5c7a5ce71f669c41d726fef742cff6109982ea96311c2d4978972a8f82b0815a5b460c415b9de23ca560384d2f7e1518d135d6314f49dbb1009d58a1227d2aab18b0448235e5f373ee6a54f08d9aa8ecb79f11583756646ea8f3f3c66e414807e6ebf17a93d875d1c221ddc9f64d8c6aa66f68c7e657f8d58c171d3847cef5ec5cbb41d7b5d2aef0f133c0eb8efd983f4310b660aa72d51d67916135d4a99b17e03d4a8856418152113625385374aacfd4b60570b1be89e95e00c138ecb5f19fe44e74325ca80ab7f8b9ac1e23234ca5e27a956d7598006ba94e4e77562f8cca2bf50ffc50090ee542d854989b1ddfc677ac8d12a040c05612a9d1244ee8b089360fce120962065c69b08bf6cf258a9778c34c20ac095d882e722047928487a05a4c84ec75f58ccfb2a6cd55736db356634b0a874464bd44eeace8e4aec1eea218696d8939c984ede5661a85258cb7dc6480fece81a6385083e9c92ccaa38094af59d63a7ab8b1b1da1191d1815fe29a5ddde65b2c28cae5c0237546ffc6eb47417395ed7b316d0c3c1e1dddd4d27dc04a91cfe98bb44d8dc455c1b39dd900320585cb9bf450567b1258b0e1b111ad5740a89f2509e10481cccf93ce14d6106f76cdd5dab992b8701e8cb2c5e3fc58896080fef4a1eab4aa63c7c843ee8bf2a1b1a75bb5b0dec9528ae6e4462cf80d3a2b20531b11761831d47c5881eb39e1fba06e2c232e1e242c3bce40ec2f22c82fdcb05c9c75911196c1a87eee443dd3536681fc7ee2f19c26e36783ba742cdb2345a29395e7ec477380d6c60bf536a77f9de0b1df2dbe21f6d0f00c53286ad123aa9f6626b5efa98032934bc2afa6429fe1c74e45f12a06f4e5f51836eafa982cc404f5bdaa3941ab2050dddc8d9de45a0721a074caf43890e275e07b671bf01d8bb8c3f40dba6040c1164f20b66b830717dc6edbee8a04ab39b930d19600a350e51f224032b4e6095ca3371ba3e6650ed6e8c7990981a553e1db5ecb4bd0436215914ca57edf1e3d30f056e509c6feb39e1b073e2ccd817ee5b38233268a91a5283b0b1c34a0cf4a1e3974ed9129b722cf40a2d3f5bddcc322e0ab80a2622728dce5442a080213453f9234145af779e206df3b0252654a87ce525012c91275600e69a596e2fbfd289b3cd1fcd2d9ffdfbd938ae3aff7676cbec9074b2e72d5b29e9b49893aa7a150086a518c7874504ecbd4a4d895a85f123d3f4309967785112d4774829c12604b0757be750b35a3c68138ba1e7ce6b733786f35d8f6b7ed53008f0811fcdfbefac7bfba421c760f5f334c75a9f4fe591e62c8a69d2bc007603c57a6973baf7bda92a65f6bc2d0c00125ea1a29006d1d163c5da8eacc9a91151080af25ce3c91bbad2c71f8ef9aae96adec7ce88bbfdcc618381a6fbd04c15d265507480d544fbe48ba0cccea7a9c252c842b5a66c63d7e4eb13b4bc1ce5ed893e51c6aeb8488664446ed886b35046920b4beb75a1cda97dffe4696a23c3ab7a7a166658bd5fb9786254746b4ea830f1d40c4b336866b8512d02c848ba430cab6c70805b7f69d064ccc95c5629962266129ec9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he42530e25486bf1801b5de21eb2e9a0aaf0802642165c069d9862b0b2eca01a2d01657b3efa7f81be57ef5a571145d60475bd4be145eb2532a3add3e68452089404f3c96a7f843ea8d2d505223bde1e68f1b17bd1e02ad0df5cfe5f392505520616f665658e8abdaec0e11114b8d62d1aa2b75453c48a838f6b1aac8bdc6f273fdff9617bd73a6e779d470c7bbdd36c85731ba4e5aef307c02ce79fb9226afe9b7027c768eaff401dd73ba091070cdffd0c12ca6fb2e6b254325c6b6c2001c36a6f96266987a1efba101e47314faf5ac3c45db350749a5b4ab45e263d79d95da3609d5fc5b62b527fa42d1068979c0d2841ceb09705a1cbf3ffb888c56a19a30a81903bd47afdc4ba04addcff74f973865ad565132154ce7a2eec522d3efbdcde187ec7bc42cc73a9ee9c5db0cc28ae0200983387ac18e9cf57bf5229748a67f932fb460ebed72c54c8b74303e4cbaa133b0dc242c805ac5edee5c59610474d3b8dbaf866a4657000e875e7764d64db4bf9579eaaa013278a9f55da272823aa72b61001a140d03d53fecbdb8a6ec2b42201f4c1802c636336844258598f83f8c712a019d665c14e7c336b98256256cba62b54aba92b6fc197a6bec2cb3bdf8d405ddc62f3ffc54f9f946d58ec4c6f9287f788edb33166cad72d546593f3938125b946e6c1622bee2daf7405b2ce1fa3479860d955de42848f013a28d85bcde3893da60b825a1b309c5cd1980658608971c829972d660403d93513816efa539d24f5f576f480435acca0f1721af91460ac2a7ea1a053c8ca6f780c4deeec25aa79228ae6d50e10398a5d92dd23209fc6713eb5fc9d432ec679e9f659d7c3fae2cc1d9a429f74161377cc4554b5e36ef97f7792561c3b5b93e58f7d5a829b47a0ff32e2fed21d1444162864f78467b620ffa23055cf3b9fa97f747930646a5b98e6c11c1b26e0a3ea4671518a920ad3fbd524708267bc1fc11ec5b316566699c298ea8ff734204f26e1b61fc10e8a24cd75231e5f7adf5f78f2c73c7f2161da6e789ffd9d3e9d1d79d3db9f8353c027be6bdbc7972ccc8819e2babfb7b83b3a18820866b9ebfd27c75507d81514ce5159e07ba43ef6a51c54ea8bbcdf3d3b4a94a2784055cfcf49a10276fca7e0c7d49b9a3e434253af987a274c66b9b29507a177d838e788025ae043228b15ebbe72e92de167b6ec203ef358ed62db9bbe43a3d63dd9ef4d92d9ae6ff7be11c6ca3fab1c9d881896560c50b9b7f21d30235ebbabdcf69dd04587755d5a2afebc1a7c1690551beec1e2f952caf882e28c5c87fb2c4fd6685b7c194bd4f65d4a5ad2dbde180f14e79e4ec9977741a346fde9dbbc6a320c24bbed2cad2de5d9831fb9a4b35274ac8a6e7dce7d43c4df42b96fb9939589dffadd72837731a82809c2311de8195febb45a839928a7e9db84eec96a2ca74d1a21a51e8852abe417a78e561aac787594b384b0eb8cc770be5be190d0feb2f31ac526757189fbaef405c086858f069feed28b1ea1daa02df75da5717f1cecc5e4e2b29288aaf100b00fa25f51f2aa7e0f7243e938e2459d400d02e571e509d9fe8938311ac289d0cbac155f651a02c81558c268eb092c30a2668f7a3dc04b413f0457b4ecea069847825fd9f0e6385afbf2a2813c6c045b79fc5cf1dbc5ce139b3b35a3e58c304a0b087cbe18f5768143eda84c8ff123a5e7c622d5eebebb1be059e0784557b8bffdd9ac6d532e874a7c3c47a35c115e9dfd2c815dcc327421008bd03e1342a443fc02f0836aea84a3d3b72a3de07e521749bd34766f8435ba77f57eb920a7b612c06263723c80cfb06a614b554ff5582631c19129cc291d9dabb83f771411d6d8bedb555d99f7dd90cb88637d36f47acaf57d701d20dd26592b90d8bd29de4b8fb6ace1b63f9791e4d471e52e2cb0242f36199e6e71e296eedf6738cbe696f5a9b5e6299d19c17d2619014974ffddd13465535b9ba2a50a0b26a7cd35d4640e2c21f463a04d107b3f59fdbbf69f0227cb7187754943fe7e369d86abd07e2eae676c36af504c83a9fd87c8b4cd8f06990d8108f6a27e722b18dacd9077efde5fe0587107435cc960dc02902fed4d47a30cbdf4d9414991729e8454476ccdcd41199b31b96a786c344224f5053a4e7db77397a9334fe78d1b30fc23619a608c46873d804dc88045b62dc3ec21a95d1ba2eff7d04e99d4bd675f9a8a331137e0d026429687c4199685361ca1493327c1263ddda645686db2cc20b24bd011167a5e51dcbde863e571e9e0a665c4168042c1138f93f320ff15bcd0abe736b38fb99bb96bdaecd9ed541e2c6f92e13a22b5ce5c3d29a28d420608a5f018caac5e6c2fdba60b40b4bb55d2ab3dfeaa41d6b2a66453f5381b2373defb0b2d71b12ffadb972c1cb503a1b2c0af7360dfd35a80620ea34e85f6cd0553ad8bbc4bbd62c720d31fa1d12452a7107d1b42e2397a4c50c3e5fdc8dd050c732bb44672521e050bd90d7e307529bce447371d5083d9d2ae97a5c7cc152b120a224a9ab0d3617545e108df07ab77c1e5aadbb441eb0b5bfbea01b065cccb73b93c28b9af4a06d7aa530a8cb605756e8142a450f8d73e6f071df91efc0c81b43728ba87efee7f861cb05ecdc0b1c027b43fe61411b2a26b9a5a7777b493d37dd10141c7eb15ff4964e8f4ad16fd502b37f2c6375c3d7958cf0373bde5893c4f8942cb70316fafb05c781b1dc47fd9c114c82a171802f6270;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd3fcc85fa532d6d8c9dd041aae81ad15c0efa911a73d0d92b27a2ce673bb43a5dc2de0211bfcd4d60183dfa042f86477890d0cddc763bb85ba5f9c5f08c12652b2c3c68febf2bf372b118fd8579305730ec1d6c159dd4da49e1ba4484efa1819dc807d54e36e757c7ac7b00e5c8b17ec970dfa7ce2442aaab760602507329820b4a8ad654648f4814ed10c21d1b43b8790a92a308b7cff5eb927dbc6a9026eb46aed5781bc750a468fc00a2052984e26cf52febe57f3d75b05cd86d2ca21e3d55a7bb34f49f6d1d9c22e35a0ef999f0dccc1f8fa4b50542f111333631d5200f8a1dc243173bd07e9ffeafcd95048999938e888b98b48cf0dbd4180afb78039b17ec2b6b88ffb343bcb8bb809746d1dfab63a36ae100cfa1c7e986486a85aeec27aa890430139d247d9367a125bc96eca4b0d525d1207a97f7e3d76bfbe25d517a8499fe39e4bb72e2614700f1cd82f74a0b4a39f82b0499b19ece0848de8707f9df59247de691dd16d108b77692ec509b2b420d620df6813583ebb53d98282f7d6e8bb45d27ec4d53020de0e43b828ad58e0436577aa872f06db5e7cd38db692c006598fd91dbbebd8468ede54384bcd1d059373d3491d18ea5a74adeaee85a48afb84107656d6499e62ef596f4a8f1e19c51bab274f598e8c4ea1a56b0d0c2387ccc0daa67cb9ba8347a16c6203334dbc56f2ca1ed953d5e770415d9cab14616eb9c33df77dd6fcc53f5e9f37c32abcf8b49633fdb527e592d42df268265d05e31c400cda4252a158e4c35983eaa8a111a71f423f72915b5e9ccaafdd75f89c8b939b8d3b9a2ff5cdf469e375f04387e6e8b3fbd40581c657b3ad9b9682d17cf25477b94d82e9e84599d8d38f88ad1fce33ccbbe8792320787a1228966c75ab6f3155aa1e4be5a7e1399114c77329be7f4b97ccbf49d213fbbe9f83b3b0d3fa83f18e59ec3b12e6a3196225a958673b7e86b9ad86c6c30fa96376180af728eb0101e1d97e3d170e0b594eab82ba6f5fdc6409ba92c3d0b950c98fa068c87a91bb70ee7699a69123e49a719ce00d8fa29b0f59576f8ed1e403d84dc9acb912a7449c07d2f565fc7fc505244c47434e7d8a68a22864db4d94b7329adf9e117c9cc08edfc3c42c1e7fd66d6d90aca8a76bb17710769acc3225ae4f199971dc595d93184bc571297432ff78539a089d0054948b3bd59181320747de643f5a5d08cfc53b555ba1fc2c0e75682ed0882f439a4082b0615de979fe08d695e92621c4b30b2b7109235c29e3f09938ee811c7c0b2b9563f2403f6ad7bc6a3d36fe114b212b9ff2c882f0ca978482056e5d58fa9d8030d0c310e703aa32fa35d4a448e2a17d0a9c1524a7f64a69f43727b79d8d5a027a18a1e7cacd5cf7aa4c3808d43372edcd7993ba2f1ccd1846cfc109365098fad9f1a056d5a1b9cbeb927e37f2a353ffc7187ae5dfda6b5e87010f737033c5db8401224f4dd807fe51db98fdbcece5d03a11a90230d2d2ee83e0b0e81280c54f3874b9afb53cafaa8ad6558cf5c324a58e83b4e5e342fdf619ee3ead3915b9f5ce9d87677e1ed77949769d0349d981221a579678e2343f1902a6e16b6d36387efd5acb650417b90f07859917c138b49b0f8742da8a78294e68ea42e32c5a6d4b943c964fbefcc85f3dcc3879b0dd39927331c9c2202bd4433a5a6a152510300f29d76bf2ce8ed10df57535a54f1cd84de3423075622fa6dc055d7749aaec68cf1c1c7b3d436de519f1bd8c9fa191b5bc5e979305fd966047c259786d8ea39b7abbc73d1c470f9a38ca36bf19454541863c8420a8cad567dcea20b661f227d084c681122049f4328bfe34d24b77870916b867fd123cd3d9ecd9d0da047ac4af0f80bec0e42b51dfc158499e7aeeb858c8e610520ac8c87f2be0b42e909eb70e6c8a852237f844c735b82004865ddebb6b7658dde453871d90cb1075dc75cd6a6e686b20dffefe64d895fba8aa78926af274449546bf3f68e26ae396b08c152879a3048b66c01fd3c5641dd082841d7701ce0d3238cc60f51c6120f905bdb7351d8f0961f49c9089cb933a7a17c6607b36d37f9d6a4b3b48231041906a055bbab4f866bac994a504415bed5039e9fa65cff73fccb4df8d7908ff1f6ab96d6f770ae65c5e9b8f4421101bfdd64a367b6baa2705bc9ae5f3cf776c899e0d804fff69dfe084e18581ebdb1c7700eed54dcfd1bb3b16c70d2cb5e17b3f5163cc832288fb6e4a22a9251aef37a8fd43d224e21781d0cc23e508453a4e55fc52b9366dd2003e39eb918039e29810857481e283416fc964e4bde6392d280849cc8ca89d0c0baa48182ce480b875bfa67188712e0d1877fa8a2a3a990a2824ae91ec6d40d959fd37705e1a7814ae8a56e788ddfb798c0d4161896961db548ca5b16f4f9852490ce0b56cc2d6ad28fc8562aeed73bdc6ad4f77895b35ebe8849af4486ff72d3cee0beac15ba34a20efe4236a1bec088aaadec26e4b106d925ff74df428b87e0ed8a02a40a7562e8a28fc61b0c08c24973527eb940b53c12be27ff05ca90a16be3db629146b2201da75d06db1d1a8e5c957c5e603adc973bb7ede09b189fcd3b02bf9d54c20e41ec8742cbf598a8d946808f305f5bd47244e246f5faf31da67a7f56f68599debdd802a2f72f4fa033ba3c62c9065ed866fc9693349ec7a99818801060dd767b97466f91f68150a9cf98da8de44306ac01c4cc7f251e8a480a19134a9216b3fd0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hab0b79d496a70620d5a63f2af90558054e114ac36e4d43c489df6611e8e7d98ff6d49590074248bfba0976a2d73f19c00d845505d5ecdb270495ddbd86bf8dfcb6b2e1490680acb964239ef565cb37224002c980c839d94e86468d571f20386abce15ca83050b7e33c25b0373c0458416c165496b2066114cfe5f21d25d420123ec4cbaa9ab18dc2ed3956fa5fda2ebc1ad018c5e1b05e0fedd90c552db50a80a71b43a0883f7839b590ac1dede9769a8d252249f40b9dcecc78ba01e28fd3bb152049a0c28880d41917fad664fe5ee7c4f3498e5ed344110622ec8487e7b1e8a0b6a8a404c57fa6fd9c76b8cc3d41d80f9cecf5e806267e19adf3580d6d335b1627a7fdba44a194370e87daac7278ce470ea610ee23838fc9b5158bf9d03397c146c69f9b5f353a9ffef1cf15f1b6e3604a9432278eca4dd871c35a47d82bf24a77cd61e5e97ccb14de4dfc990d93cf8c2d66b9e19ffb6e5786cde6f8ca925b362cccc87521a1913302ecd1e2ec42a4c41eb9a5f2ca89c63a4d193e6931bbb90e6263d687886abcb92fa87b2374f85c9df4e856c92c759fe627513efe4226171a69497d6301c69b673bc21d9c6ec93d9583f711b373eaf70ecc9662944d59291fe0bdae945251f40433d777226febf1e4ed3f7e87a3620be9e7eeeae17f2d4e89dc13c38d4cbdc12201ae104ed524f12cd97ffd56859bd9e18ce80f89fd9b5dceb08412a91a04b2f14f871a1554ee30831d40ec67c952ef27bd5c678e989ca5181076025ed099fd01c2ab029b7cba3d9d2a4086467063e29e1b249d61a46d2f77574d8461ba907d44dcea4ffa49e50273a31fb8c5882bb28992b4d7c10e9081455df96529627ff0d3b4252e16cf7ed2e7e1fe68c07f0ab82428952bc0d65f19d8f7c29fa2beeb765696cc0561b4c413f5a2884abac23e05ec3aed741bab79ffc3ec0a244bc7bac5fb97308374a13296bcb56d2b5d34b487803157cf3ccad2120ce53b6c13fa9368d005858526b00ba120db93bf1e45392f640236806752d23641e95c7c08d332a9d4937bd2922d987b86c92f112e6da94fcff001fba8d7ddadd0bafb51ea97e956d8c349d6cfe96d911b5bb6c73305ec7b5e516c3489acb59651f3e731c0c330eee5651d4528621604349425fcafe9b296a1559e18a90f672f14909f39bf9c5db057056ebc640c9bc86d9fa27bc1b4b2734a71c508b0b56e015c219e05468f6837ff392094edb86cf44bea001e0c6d6031a7e0f632ad02e6763578c986f56fd43dc03e6eede56893a0370a3013ee7bd6241a99c546a31094d672370a596934a5e63e4f5b8597a72938ccc4db5ef303b96673b1035e1f5df19aa8af0fd4acbb164d32e43acde88b9a51eacbcaef5b67edf74697b08258f45de60c4a294d69b4bd306b9dd414aabd32c5b5d04ad99648cfc8427fd36ec75cbfcbd8b0d5195693ddf63fecc9deb03736045c1e509d8b58279ad9e2858d2932463b7e1e253bb2faa5bdfa01bfc6888ffcc9db943d9ac0acff65b99dcd766b750c4c32ca763a79ddeb6834040bc19fd823cbecb3807fe9b4ce23aff8ffb6a3db8a8efbf7299b5f1e64dd17069c1d9fddb14427910b29079076b4db2fa28a88f4a1f68c8bbd8c10571b264ce41ffc52eab93e44c201c667e5ca6c351c28f5fcf8eb7160308fc03cc5641bdbf98441f7889c6d4f4a7d4a2751f8c6e474e232097fc98d998082744b36ad6f75f8bc564af88f416a036149431a214834a64c2dd64bc5092edf8bb5bb78c8379bb400d953413cb2a5151d4f6ae19d8445e68109eb9b630f157339448966e0ab9e083565c4468488b205ef437aa79b3ebb8af8465abdb0231c2c529fcd981fe4db300652b686836445b84844e487a0dfd9ad0553fefe1958db57a329a96226a927761c84302e2f2d088cfe60480901d82f41d49038f6aa73cc7f7eb302832571b0456797a4481eea2989f537a724f8c7f7ecac3a367b3274b3bbe735a90adc6129f46f535e4cfb3eb1777e060d27c4c10c40701ce853c10d5f5b87eacdb8d01486c64afee087ddc55392662f615de3b02210c394e45833a079d8fac574ccbb8f75f1251a6f53f544be8f463ad6d596dd8b9577c45d5f3ef46a3c3b2300bd41b03ded601b775a65647c4a9876b819e260d4a783d2c675ddf4db4b1226dd7ece0cbcb481a2ed53301c51365a73f2a8e9587ba5e122f02e6b392ada8efbd2479c86db7b4687f4122a36768b9169bb555d41b311a9b2600c20dba1bfe2f6554016224cb0f52be0cea86d637121051dd167fd85e9430b80c7c6f8d1848e5a34c43fb7f27bc7bdfebe68be418eff5d5b5732e5f0f823515f5a61a4b1737898d8962674a0f1604eb135339258fcfbe7a03b0e5745d7b4cfcb2e4103be38bb57b040ce1d8b8c2be6e750e36c9bbc5217cf5da8697c02f781b9ec9cebac842fd8e55c14660112fbbeda2458dd2998523c8fb9f37072ce8bca83cf8d329f9d85f4fdb79a361a09f09dea098f8bc9ac18152ab73971d8ac1df41046560d2555518e0c78cad01c3fa152f19a5b1705f53bb192b964b521d26d2385984e7fad66f9b4e9af58445413fb5320de8fb73ded54bdae4fdb66e8762fd8db0c4f2780664306feef9f0a4ccc3ab1a55573bb5ea23e2536931573aab3b600b34bea3cefd79473ad14028a9f0c216b35c6ddf4712cd964c91a87d7509dfa8b11e9826e9dd0716b0480b3f208fdfed76474f4dd67c5d7d1fc801b42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hfdddeee9b969069d30fcc5dce08ae3188006a209f5c4a0b0ff1f7b3cd2851d230709dfe0fdbf9ab1e7bf5de8b595ddecc3afcd4290345da77e2e61da1f53448d8c13f72b3096d81c361d00ba90a3a663ab5f691a81245c746aebf0b1571fc680124164b99c9d12da4c4843c711511cdaa3b311cf9c2fe1b73df18c791263c19f9e2e6fcf58b5e84175572d8026d4fa7a4af7fbf829912f60034fb69983df99ba1e940971d0c3860a0a4a21fd59d4c7da8a63de3d26e9ceb976904e1a685226c99a7b3fad80d88c8d625ca0581fbfc3ed5cbd0e42a4dcf494862f29f38e600490eb71fabf554a86803e4b8bdfc01f4ca8d79008f839b3c632540564d350285f46d1d85da037e7b40207037e301134a7eafd77bbee00946cccc91a7ad49d52d703e29877658642518e1af4c546c81fb4dddb636eb26b8c3cd3f488da797164c9490a55a08b69439c61eb23705794fc17220d606766c6d62885ec2c6e8c649325ad922c9e3d6ea7162adffdf44ad54021a5e2788c66dbce69014e9c75dfb278abb159ef8a29c843056de3ae8bb2932d92fe4d8bfbc4c632c950c258fca5796b0e61d702bded5ef777de4d36625639338302383ecc51e595f7cadfca99660b74f88e8a93d468065dc18bcafe170b2a0fe9c2d11d278348bfcd5363cc011a29c562b29d4f16fb08bc7244eb143b68b88c530cfbe5be8acb3ff2e38d1e4f763dca1f30920456e1a5e42d0d1796f7dbfd2199d6cf9c21852d4f488e040b25a0d3eae232f2ed935cbbd47e2a9a7aa5bc37784c8ca8d99d0ce8c8b5c02ec57629139d7e97c83284b8945682fb652ca15ee047c360ceca776ddae2a7732a074884fc004aa2a9773e02a78e80b6b06eeedb62bd9c4be6682cae54d6672156f4574f8c4bcfe2f3b99c741be560da6270b1fcc121b780e54b3e57ece98d9160a669230d19920d999e00e88a790130db11b37ca3d345d4cf5baf17bfaa73b492356ab030e1a14abe97227f244bd9543f28807727d29220d7da7d97148aaf79b838348fa0a297835777e8cc5a07f3ba0011f37e52687469e72d8e7396862ae117831c9084fc056b85bd4ce616ca604aec7ddb061e399a8a005c552c83cd2470eaea46f85da7ce42510e503615704b2b2796858103f67acc24a9841a7fdfe02bfb3160457d8ee444d1c7f29d33063b1f218c342734e7a144703ce61ca47309e47eb7cbdc6a762e06df2ce927d30fa46774281ac0963a44e5de52aaaebc9e1f8faf493406f96f98011fd42b18b7aa4399afbe4e8d9014cb5ae1bf78edc6c9ab59c8a856239beca8aab086fb70809de4782f03bac89898addf8133c44fc422240fa3a7f58c5156a2c169e23550b07ea6a8ce72ce7864197f79b4ea46a16086423d3929d7353368f00f7dd6bbac1de5c4ca2fbaa48456e7adc02116bb47ad3bb21ca42668ca9598083c60f25fbac83071c823e0eb5b7e3e0b65be0df7c0f942061d013778becd9c90e2f6dc0c0a807067a94787126b1a11b63046bbaf5e7028d3a40368f9ebb7806fffbc86f45743b2b9b04c8cc8650022ce5d1f25db1a0ff4ea6fe03a2e88bff19d6dca20b54c937dc78fec0b0eb54fb3b0eeb50d5bcd29bc0cd4b5c18de64fee3094655d4adcf08f5952b8d5b104f11a127b4edab0ddca962782ab8d49f5a52ce6174a79e220772afc8836339389621293c319567ede89aac2793974ad2132900a70b3ac7b55a511eac9e1bb2fe6101aeb2769165958dd8893aae17e8c7478aca3ba1d5d47932894a62c2cf27679115740add55de20f38a01f34a65dcb75de4f0df497150b1ebb15bdd7cf59ed385b70f7b185182965139eef4be9566df0819e16bb0483d65b0d982fa177dc6861d8afd885e12ef685c0b0cb95d6c2124e5dd11a0f20b41b6acb346cf17d6ba1c900f86a121f3af8b4783a88a5ffef091d4b40d27a406172997045ae66b781bd128bcd480162eb0de0b71ad2ab96dc0d57ccd503b736c462c42fa30c90f9bdeda311f35f12acd074f80ae987600eb2342e911d86b0e2b569e6f52d460e30752bc0a1b6b860e71af7459e0a774cccbaefb833286e182390f9c6d2637ed009df9be5603f59d1f67ecf41e650d9b4e52996c9ea29b2ead3177c081ff4777cb40d87aab2624395ec236c073a4403e03ed061f1a5767e811d195f1e2504dd55d3b5d67cb2bd84b7eb8fd8c92c7b8f446dd8e59359820cc4c2d696e3725dd8c6ed85f319cfd6d4a3138b22ab2f41a0d0c3135a1305d80e2b34ee3e5a7a531ded5db58aa2af05b19afcd9aeda799073ee87dd9d519f744d066702f8215b65d63e5c268011e14fbb49bc0d643717586f5cd202107203ddb4383c744ce80c17806634396fa8ec53e9fbaee1773f635418711ed2e39cb5a83afe086d7250ac5aa8ee37911b207e5fb87129c68315bd4738f3c8b1b9e924dbfc5ae0548d91773a5273ec10005014e98b5aff5e65877566a8f1773f620b4a8d8ec5104ea0ad584c2b47588983fc7ee4938924dde2c67e5655b786e918eba4c17c152f7a999142cd375dfd74f284e416f72cc4cadc856a437674d7772fc7058fa5e3ac8cee08eeb1cc7896fad048aa32c7ce9f58dadbcfae7752c03d1017a1c7da1353b753566e0e8589552e1de6a48d1ee806355027e7c2312d663b573968958bf99a903c68818a08ebe2f9873057f171a7bb56417d663fe32d8765a87544ec267e2c0026c025460ea7f3c103ca812a3e4f7894475ef69399a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha03a14a81ffa37cb4aebe0baadf746810fa49956fa947cb20a505729b303e0a3465f1df93e77d29798edb2f8aecf2243484be308fbb968b21aed42b640d53632676133bdc88311d2013490f675857b4374970cfa8550b32db2c56d2cdb1ffc565e46150da9edc5a6074ad0d8acb0eff1d806af3b4ab1daa49348fc55610fae50d6f5ab2a15277b0f1e8faa896666708cec1910d927429836d6cf138fd07bbedecc4193372375fb33e1923ca90748f23f1a924771805b2f5afe9a6e3a69d9a261c055b9db5ed8f9328b3bba470a013555e8ee993af994331489007d0abe55f0bd503e0346a8b9bf4901cece426aeace8634dfd831fd4e1fbd139e1af99ae4e100508a4054d0689058411b642a3719df3627ac27fe73bb4ee0f19e3586efb2444a2eb94b1fc44b3cb28b250a9242ddab12e1681199b1c09c166a89632985ed44ba79b0955be8aab32c2da17b0e8eb2268f41938cbac91afb327cf1184d14f1c6363087fa8fed8cf376b50b90c3b5b01796e7715b3220f3f3655b2419cc4eae1b2d12446cc2e74aa62eaad35c8e7c41ef8dc5ea7c00e0fd627659678b2ad87c5e6310f68a5a58d3b27932197434b5ff5485c548865135b9d9def874de35993f11b9f28e752d7fa652d59369fd1b7472ae438f84fc0a9b665d3c26327f2ff972e1b210558c9e78656814d78218313bcd8457af2495437631d378f17d5f562dd363e13fc97c66d41e7b222d447e98d98a7677f1fc58f52b2be420351d7177e93862aef4782fdbb0bb53e7742d2989d36ddcf32337a50a72f62e68578166614af3ca83deb839e682da93c7832f263d0b8c32b1ccb885e480bf2ac0d43fdd41ecbfb43171bc3b8739139b16be0b813290198fde411371e1f78179ad86d2838a9d10d5d48ca6a91fde872f9ed1df1ae80be29d8c8959c442e9a1f3376cd88eafb0f724d138ddeb9d65db003abdca2500d668d0b429d06f494eccde4219678dbc86502d760d91b6b88f2438c668b9d26365e745912550d5f58ff9088838b38ae88740264ed8e07ad89a16017b22e47da1bcad5834280c3a7b077f77ef01adbc317a61a686d1dc21536ff8416aebaa61305775f56f31ccb0c4a4b6bde4df525d3b2d33f6c72bf5ea0be164519a7f56f3a0004fcf420d3747a35f101a80b413041f3dadf76c776952cf1d6e17a7aca36c0e60a9318622175bd7b29ac089d800633a0eac123ffe88534c5c47a0db1b4e0057faa556f4827d161e865bccd5b099163a44b2b4c4918b1b32bf2f8bae0636bef933609343af7655833e44381a7a0d65703650f264e04a190f07e3ec1bc7f43a8707643c83f157c62c1278c4fe6febd91f08b6dd5779d65ee5fb39ea748f2df44ee109ecd2bf82d2ba7ac398075807d390ae7ed773534c5292d3276ac228ddb3b3bf357519c2c5627e6668039addc619799bca93ef3000a9cc7b7d4608373a2919f416cbe8d1f84f453eba9bd6815a60420ee74a669e1f980f5795d6350191a934879c27196744a496d15e8de909562b82d59da7292bef1b61848534234917cf9258f1a7e9a95cf595fc70344317ffad2ab9bb643b2cfc68dd64825970209a7138270d625d24afb38ee0e272c3606f209832f83c6a7cd9835219ef327029fec890c9d6c53f46e68ed27ee14c61293759a299f8f5751c4c6f68e24b95a6ed7301c5489735f2bad3d1782e0a0565576f8d04c66c04c4891915e3cc8839bdf160e5d43066604fe0b8f09b921af6228a98f446dd61ca596f9443465cb2ea6478b2b36ebc952ae36cbf6ca8957ebbc04360ccd27d752538f29c1ca547986e36fbd6d464e54abb1c8c8916b928cb3442b19e13a3eb098f3305867b80ceef51e48b982e33f7c34adff7d65003f046ef19089980bbedfc1ca8c18470a0b7ce5a2d338b89b19d0558912cb2c31109e57c771152e458793791baa5a28487980792bef8abd78e19d2aac9120ce83584fc89648cc2925bd96a46ca3c6c031b3edaf3bff1a01cdbe203c66a3d36fc58f70588c6412bd168dd41a450aeda6025554070788816a28756c4105c2e27fa353e832d80288a84acf686ae6e004b62cdb03fe7279c42fb35a757dd27e38dc58b2da17c2db8150e4b4bbedcccab1dd9fddfe3c30c9eda6fdeb52c0e682cd1e573f2bdbb09b1b8e25b28c0bcca1758e03b0fec6177ce7dff730bba152f4855083f1bf18c41c4c3a871bcc94170c34961824c5459f86e58e1414a14c6465c43c63102eb22138c19fb2ba04a95593af7b190bd9009df4a2c227b15ebe681582129469e604566659fe246850793ba5aae25305edd0c68b1773064bfd78d53147c327b15e44b8115bded1455eee81503bd3bbcf9763fb3b43ea76ea27a1efddcf6c306a31c87aa4eba9e64c40b23cba9ab33f4369480b9efa1b523723e2edf20ca148d28ea9edc86bf2f9612f92711e2c48ca37479db34532ba1905e1c1c05e892e5645c118b2cb15c4ef120f62d2160fb1b7e84be278cdf862a6be120af97b998a26dbfcb7385b80a852dafb7e79804d10aa5c373ea47f80d105389da0fea16f16ff60eb582a7fcb8e043037d5200b9781330632b5f82002d75fe7bcbbefd5d5828fe4d12883d2136b77d2ef0bf386a830f5d1b7f20bb22274062932122a75e6797bf561f87d65353f8b14b73df6780fa1d9517ca72da4f1981c9f3982cf2e85194bc04b1682511c48aff11bb4ff1320be8c88230edaa0ce83307b19bb78f7bd0e0a5610babc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h53fc8fdb4b16d2bd8373e1d0a5b9575767561c1025fa2fe593ba609807ffcc2ffb7aedf4f2c76e4d52a418d1c88b5f7d9126a68493b58d7b318c562905e821e8c51b05366f8f74b64962b1b70d4c6d8de21b8e415d18b08b72d545618b75e8dea024c3eedab7dc7042339bb7d2548f78874962c6d09cbc761bb90c141ca0076988dccbdad79a90b53c4297d105db4fe83cf923c136ccf7c99df542d1a8d2da1d4cfb33a325587298dab239f346c01eaaf0748f44cd3a3522d6743a48860084aee3ac802b07577f1b8154f2402d3e378e164e48d75198fb08f0100f963cc9ba3c6b8460f9035483d326cb7f44cc8bc40dffd53ad8be390ee76a8c47a6f8366f7f9c427b9c19d3b813708c7a5668565f62260cab4b57f15975ea161c31368e7253f1c65074613d52ae4f1ebd61cf547f4b5d8e342e53fd1fd35a8c3b796d9f755812b02c653376f43fac240c80b4448d27450bef97f8e02ea68756cc27ed859927c3d03454dd90deee54c02043108ee5acf8cf6ec359900ebf215e7c9d54092f7bb8eccb82a892fe351d5f89ec785c78292090a825eaabc795ac96b4931f002dbbca82d0052a63400ebbb6477372915fceb915d50c3ac90f20c39d66fd27ed3fcc262c6d88e5537246b73317f46afb65faade6430ba0823609ba2ee54c010b9b286cbe4c8e969f424517f331fb8a3e2f14943e56c2ce8fc6478902b9ee3b6071ab0229558e1f3b524714f60d0bca17f1eecfd7b03970fedfa18012b6ac3378a931624e2456442e8aadce78dd213ad0fdc3c6a64fbf0088468430b7bee17c8b96602756e377838cdf035fe32c2e7e3e5da68c782ea7ac6d33d3f711b6858bae6a4a8790d4d1fafcf3ea7078dc9fd2a2817353b6aab2f5c609764a2d5c99eecc20548d633e4bb1e74ef598812ae7fc760432ce3195247aa5444f68eaac058868c3238befe0fe005c749bc28469cc7434ec5d566560e4eb0d3889410e23d951745b96f2b47cfbec2585e1d74f33636b806f45c662577f32a401340897a58f8faf79d09f8ed59967a13a39dadd647fea186a33b213595ea0f05f2f115c0c26e684dfa978ef1327b06e4b230eec98c3b3f6cf9ad1808e09168f31168af6d283ae58897b87af67232f14d915ac797c82efa9ba484d9eb73488e7be8a5936a423a82acc5d75648b7dd0163448983212171aa5600a5ad111e19de78e52973fc47dbe98fde97107ce590433b0621a23cacd8b424c330fa4a7e6ab77dbb00c04003c78d0e81a861f7c02a25ecbfc9f2d8b45529d312c1618dcd7808f3beebce053b85313b0bed8dbb236593a5d1c756138fb5ee0f855c40c3fbde713d6dee9dea9d01c338f76aea08df1f66e9f9d7ffd02983325afdfe70887e500725904fb5ffb36dc5c8dc417ca9e765c2054d530ccf55398600142cab95fd79ffa02c1ac04c2c7c307117274616975adef3ecee6910ed7124e5cee9d1fd12146ddb9e5f79f155b197011a11982ee798b41c4e270755c15488630a42fcd22bb30157507ef67e54c4a10a3b091c67c4c13f371bd70eafafd79522a8fd2b3b75c562df86eedc47c728cb08311ffb5cec0fe2c71386ba749a5682a36684cac19eb5416e58ce128d5f1b4adb8d735cdc98c5f05c2de6e14fb5b674a18c9f3215f387458dd8e8d0d8b3c360b4780cbf4f964e7566c642deb610935fa8bc0c9b0ca39a76076a534f226ddd7ad161ac79ae08a15bfd78b68b5572f40dc1a685acaae5f520cee808d3a7d645ce88aef1ca70ddf7528bbdf159a29ce9d8e73c99e51023909b10cecd272cdb4244dff0fba1dc3648d9f94b3999dc331f976b734a45230c824b628e979c1b8e3a4f9f10a9e8c854c94c54e48c5841b93f9277f9c142a76882efccf1d7976265bcafef5457db6b4e517350b81d28a7fc11f73615cb869c36e3ddb30a65f1e6fb1dea0a961496324360a79827447eb00b3c737cbda271da363279c390d90d420908bc0b4b153d97990aedfd5e913e8f837a98551c55d2710630678c526f5bf31018e13f2b286bda696627d533424a458a20db2f38fb00939fd9e8e636c3c915ae9343e2617d9c7d05a5d80c621d1fc259d77748a359220e075ae08e878c19360644d5306ad5837dfeb9282925ee244a4f9880c4ed42df62a7cf73d0755c343f1125b69e0879926b80bb3898aac5a0b130734ac9fd6bfc8708d783e77cc4e3665930175ee40c7e95f97918d29f067a434d6c18d74257db97b829185c8b659277b4b76ecc915108b95a96bab295185b406496106fee532ae42465f6a4fed4d6412f70540d0098fbff3b9622be5ec51895b530d9b7aecc82fd9098b66231f3075e19c740465462dcae9a309924a47e8a734ed097ff2a934169534bea8e3777344157fd8d1717c0c7a216695517f74f9ab9b61ee7764a4724f6c7847774668bb89e5a3acdf59ea0cc1a72622d22baa45c41465452560be65f3c2c778283ea7dc78f92e8db283d54d583057b13707100f78a8e125470a86929d710b48ee72654873d5399bd248e0d2a5cfac372f6eae8726094fb8714be8ecf0d840edcd8fd4815997f06b508255db19bdd4ecb8981404b868dd86d29ac60cb9a13f66cf698e24fa76d2f1807ff465afeb9e24fc5543c0a9dae961456d2814f3a1946045cb84fcb2a72d34640678ea8c39a388c90fd52a3eeb356231b4832f65980be8c9c63471e8d9f87f5fde3385cbf4cac9ef1c845f05d5876e60a7bb76c7b841869d1713;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h668679fb89a48789dfbf0fa491419ce2e18ebbd297e240c4f64bd8ba97f1e5dc50ed18f566a9c2d8b13be1b4fb4143d9fd3242706bf2e3b48f9360c9d41d5cc4f0f449159f43045d369599db16ddd949560b9ccce4205d9967b8ce82068d79d75ae641deb46713fbdc38e4fe9011ceb8d2d21eb95c76f346b985c085b820ad3994f1ccd7ce99edfba7558ab9628bd64ec1b9ca7e251d15220d2758cb2fa16229646d6e7bf201e3a14a313bba0f9615582c58855f19eeefdaafc89e02f8572e5ab0f4b557649d88b776839af29c731769e77f41c662c1415f663c5fa2f54fa1e113ffc889b0ad0d4149334f4a186f3d4d8149d826fe8533daaa37a71a1eb1f725016250a13d851b51581a4e48a7b759d4263a8dd79cd6cb914e85282a08ea66f7f831bc4516d960197b3f97933192d3b20ae8a756e35e93522cfaa4acad924409edee723bd1ac1b038dd07a3e959f52111a74aed8f4256d7919994d24e0f699b2cdff73403391867e50a166335f1001648a0b81450adb5a349cc4d04c5954389d08e3453a0769d9378c76077cf3a6e7953d5df17c66a6391fe12992a74fef08530adb099fea6e290061a70971c40267ede91ca8b32b6700984c5ab8f0b7a0808f841541762973eb5230352fdc6373af702538fa76024a07c4adb1b42eadcaea3a0269823250eaacb152ffac16d6b0d87826cee82a6e8a9da195ce5655e98ff0e0ed284a03d774c58f59fdaec40f54b3fe0d100de77c0f4f3ff1220e9618475ff7d5507c23879bdc55b2990d8b517c234c804702399fb65e3411941fd2f57c7c8bf0a7a9b7d4fff39ae8f2b2a268f723b6e51dea59dfef173f4928620e66c3f41da9cd3a7436f5eaa99260ada52901998d575fa6b1a8ba8e0fe01f8bde981e9c4c876061c9d3e4059b5a095d9a29b62d3937b18b1f92e43d1daf135a88a0496b96b1ad4089e69f351601aa6e63aa2f5595ee19b00713343b4fd46c2c51e76305cf7cee4d6ea8c91285c8f6240c70cd557166a0a9c7f943baeaac492ccb64c95d8489606cd30dd90b51f1c176f13f598e4e923857e5260b52d3f1ec3ec5c6e4c45d8d09a52a9eb3b2358f77c13ba59e4dee513edfa1fee4a2bb3cfd218450f13a3d4d2892dcc00f54376a9bb3ab2c3c8253bcebdcd5532aba53a4d331fa027a312d1891c7242205f565161f9246e54c60dc5fc340d15b7c944f4819057bd9b677980b072d5342c10602803182031c11c7861f44d505452ff1ae0863b33ab34ed43e62cbb02a922159c776eb176113026bb8dd60b6eb62d45a61aa449658249565566d50a1f2421ec880f8c9bf7ae31bbc900165dcdb85aad1b26a41bb84592021e8ca61a2fd1921f0856bef8a61b78e9a58f48dd80de22e19bc8e40f1437e2ffc2a451a4e14a8678bb51b802aa7d3165ca2b03582a973848dfb296e41f9144501016d476bf9500d8c389730ba2116af2c02d296f1bebb14d85f69adf82f0c863ecf9ed3aa746dc3e8f6be69317e026a425151092c17a22aaee4966f40b4a30f59700d0c7c256bccc11fae4eba01efc7c726e5616d6087c53fc7e9422f3fe5055a7c9efd21198a1b899a9a3dc9399e0f287b3891859bb3636062e67d0abaedb3a66ce86fa17a9f260a88b2034176328a1a765d9c8b76790b88c29eac2a8abb96191cda6b18a766f76281368dfacc69350f5fccdcb2b7806d42c337b069abd99d6561ecc0f9a9f236da0f5120f68b41d1b438f65c93c8dd6ab97207c459362f40051b013fd1c94519e3932f700d8d14dc7fc3025e8378c064b5c5083ec6aa7e29a4a5cda86207a70915b6f531dd39c8b9626568bd66a2a63902b72ec5fe7b482cc6ff114642a308987d9173870abde0208104f02faa5a5a952587b6fdef5911ebe05d8fc0413d72f2d8a39bc0c23ed0f4adc5ac56beb50e6904fb22982d6e766a245e326a74931bf89cdff1a5213839580f881d2fad13fd74b5c4ac8702c2bbb02dc6dd8a71c831bec617308d45577b473fd42437d38f9f40ea2636b6ad84adf4e17ae4c04044d20eec57176a49a660ab854a2cea3c69e2aaae6d92aec85c2b1d405eea2439ab823e7879808ec9e04dc3c27157002db567b069d4e7bfdb9c9979c0207b74461d6d7d844fbe17a09f53e92e0b5785a8f35db80ef52b70fd5c7474b6ca8392c08965ee435d6e5ed114518c75fead64a9ea75a50ac1f09675ae864eee0ad1c4aa6212c0384c7cb3911069d947221d560edf3f3d528eed81a1d801ffcec8a6504bd77ebcf439e6181e3b6a42f03e8e584d2b9a890ec7c67daf413836b0bd28a129d2edc2083dc64d5e620ea3365b061c7203c87adfb402c768945239cb42bf76c027b9d72e0b51af0095d606fb5e4f489afef9cbf56df6b0ac8f0d5444b3b8d2f9e75a8d259b8b4a13aece6187cab80909597a14eaf9bf2535d5c3e868af94e6b501e51cd57b8db798b3577e8321aa692f8b48727d391e3886ca545ebe6424557e39fdcdf65586661b0c87b0e14d1259f88b5dd6da5ce0f02c6c57170c04151fabfe05e0faa406ba5c58fd3eed42566d85c146c9736cd50b3a8bf801688c636a69a9df3d70a02d9be3d04f5b72a5ac613eb6ff47cee8f4b18a8e856082e4c37d0833dc103e10aeba1ffb8cb12e3abd226a3343e7d6574d6052015bee831502ce9849d721777a90b609e2f9f4ebc732ca6fb9402cffce55452908b90907d053f6348f12a07185e54f3a44342f269c52329bf709bde6dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h60fa535bb532e30934100c7a184332a2bbc9efe0ac31a178b8905f47d55959635f71bd55c67ace96aefdef2f3be9870374dcaccf05dbf3b89f972c50e53fbdb8184e4ffa39f3c778d0ec48571ad6541a774f4a802fca1f5a285465aa4146d9b630fd47170d9c66b1ba17e9bb654495dbec342d4bfd396783f3e0d1a00e161026e1e7e23fb875975cca48a52f153e6f3e99b05c321fdd02a32c458f8ac255da467bad85006c5c77d53c507b07aea8a9f7e588ad04eed45104794c4e4a71d82d2ec215482585f2be1c88f04664f20f4d4d5cc5ee882d5fc3326bb6fa937d06572fb92d7d92dad49bb8f1c43f8e50ba3a4876302107208c42838bf6dcf0d6e5c7d0d8d14d364fdcae6ea1b4cb28c9c25b09cc8a142a2642b817869a4d4655a31d8ab20fa3aba628700d30e03b560bc8a00f82cce4dfdb5e404e3fa16de4352c25534d06034e5b10f2001e18af808bf92960e24cd80144fb8ae1a7c6e8a9e5ada222f2161bd2467acc325715877119b0f8407a6daf122ad54cb09b92ffbf229c8fb0cf38aa78cb6ca8ad11d70262ff92672967ed36ef12c81bd5711d89cb2f543131448fb7b24e993402773f0ed4ef90571174572abc11753f3ecbc8a116e9fd4773c29e9dc039c9d78fd252834392dba8f718668fbcbee1c4ad8dda0efd611d11b1a2989aad20f46e0449934f15a9b62924eda3e675076fe64723a440edc34dea8683e494340f7e0fbe5b84dccc42f800c833484f676b8c0f818f5c064af8afeead72c16a9e72b628d6af4e03a06a55809f10525a00588765a9b75db13298ea765b098ca50d4d76b9e5349fc93ec5d6a044c8fdbf4747b8f702b11c9f0ef9d31a0ff6e7bea01ba3b399bf268d83a5c6cdb705fba4668bb2507d3a73ef5e5606eaf88bf1c938ac58bd09db4571f8226571204c910332facd9e51d1202be0402478c7febc44e928b6e1ff33f9ede6e6cfcad1682ed1945449a5fa3b1b2d0cb161f70ae4c6c2e0d08e9463aa7a98f5ddfcfc64885f23ff970f66b0ed68248fc922fbaebc864b32419d32b93d45db18dafe6534c8621e9e3b4b8e08739ba7214c41a2dff679c533d297bc00802e2f2d593527f2aac24d7f5b44823d536e1933256495e878652a28c26ba479f7e22a19d130adb0b6e22253de3c298c99dd227f0f17c6818a6c1aad030cdb61247c4bea8d87493984100440171f92402d0192157777e3920efed6187c80891c51d83692994613517f5307e619fbdbe4004d7d8370742d13de0e31f48894c0ea631a5f56c577ed9e069851973731ed465e82cc5fda74ff1dfb5120109cab20934a2e8c064b6598772797067247e8b2d5bc85f7f807cdb891155ce159a1998586d48ae43ec846e6f473f474f0572a2dc4b556d27d51fe0eed72c7b90916c5950b7131dd4930557a67bd47954484cf8bd3a5c40aca17c846dcb414f25bae9ca53e1b2e1beacb9c8246a974795929203ca1f17fe08093f5ec0ccd181e14c899a3ab93b4f9e8cbe9fe6dd855501d0b18f82e9d9ff62d21bd4d1b4ae0fdd91d4abebae9ea074c2892f4ac840624209c3750700b1422d2785e7b5c92f924d6df07a007ed8c4385900673b1d78c1a4d00b169b65c4ca407d2e86bc0c3155e257e7c8db2a591ab511f49626efd4027872ce10daf864c8ffe4b271cd580e60f67fcd00286fd2cb2357fa493977fe462faeb93ee655ff8bee2527ea3d0e83e3da40048f3c488f2f872b59a136e9b30a646ac47e20c987d74ed98f4aac25dab3e7d64ac266743be44ba2ce2fad29713ce8a7e483acf0ba1e74273d17ae03927a6ad33c788c831f00da5ffd561e24d006c82aef12bb953f53812b3f772014f8973592af8dcd18193eac728ca21b4ab41e703883e2f4b8d692f8de57dac95d592b8e09b1739225728205fbe48ed0ed5c31dc4398a060dbc46ead10a4dd5b4adcff690c46e0193b00a1968dee57de70f5fb2edd9359f1a96afd60819ce5d420e74a899472219e3c8c67d2b67afeb3c24f072eafcdba43e20ec0db8477aa4e50c0272ff7bdcad1b7e91ed3b174edbbb928811360ade6efa02b5ad7bb7543ad6c14497c4dbc6c9aff686299022bc4883cc4fe692d0c98264c6b9c097709642d563a1e5bb9f5937460268ea0363710caba455ce57fa94a07892b982e088c4d1cdc962c7d8779295e8a65308020d32723fd3043b4453cc18b7284a925427ba14bf4cd3ca974a721998efd11353f59306065d2dd10badc7392036c6e022d03d10f52f5cebcae5c6e3b075c00e557b22d3e55702d7cd32dccc6f51e7d21bcc31c2e0523dafd6f76b85c357a9bac8fe702fe72e236771453c7767fe62df076dd4a6152fb388c0fabc7b463aded0d760addbb16dea187cd6bdb7c9d44ad849a55245e93efda092bf55cfbfb81d072ddf6855b548ec5eef13c0f868e0ca3cd0dc35b85933552e53c3545babcb2c127116a630a2e07d5c53f17ad678195bde6758c835fe653c0e9aae5538798ce1d0788b021022262d3d4ed0d4674b0956eed0c1a85e69541f3eb9c7b746e64bf09af81264c44e6e1c0b5710644798a5156564e24eb3b073156f6a5dfda6004378cbf7251c1be4d7070312ea51528daa534e1b88066f37da6f78449e5361839c5670ca205342ed4b97c35e297bd4e323df40d0ea0490186040a737b6b2fe8f71ec596a52bb7445b9aae3ca10ea20319d2188da2eaaf28a32436a5418ae6a71fc44af57e73bda6dbe6a2b0b0c899c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9b0a06770ff0d79b05281c4fe8f0c49b9ec341e88bf4e8869bbcd675b87c32e5bee3950f6e4cede1a7d91a54e652e94be22906173b15004cd0013d40519b06eea5c0012b67cd8314ee0e5b1a74bc2fdd89b56cb472e19e819384341e5aae2ad356429df30a1a567ad472e60049d5e7fec0e6f1b55157f6efce02f3d8d16535f556c63f32dba886f37d1fb8eb4846c2ff292f04643453850964a2aecb19bf0f17a9c10649a1b048862b1eb578ac742ab916f27894f5c48c4dad53021dcc39d410556216d7b86c9f3dac5b83cd83f07da4ff30584a63d168bec44d05e7cb1a0518058bda0e017aea4323770a36323c3f3785be73c64bdd0d23917da5761ec9e5ec9e35a643baacb53e681f06bf28893212d1345257b03f676ac5f45332476af274695eca6b4389ff7ee5d78fdbe1a07f06d1487a10dea563ffa6cbb678b08b781b20ed57d0069165d87f953217311d902d8c3d131cc47e8c0714fa571fef15d2d47d3ec6ad8d9d5ec2452f048b696fdccca5909ae0e6687848fd863660e0716870883a4ea72153ec487c50c5fc5a11fe8af28b375d6a3c45f722fa1406e1692e28630b37e62fb899b33c258368baaa68283afa106ae83f787da10ee536b734ed82edca18450e46446be2205f4cb668c7fc1b8e74a3b772e5c9607ec835b80b9a6c771f0672cda45f5b241508800a2f7aa5395b9cea2593527c41e0711fe65ac61a5f8d1c1027ccc0fce8cf6e50ffdcadae71404a62e8679bde94c75080123fe6377ee957fe529e7f0f8dd0964bf7853cc5f044d6427f951c4b831f8e6383c3f12bc1cdf738c00db3929b5e25d04b689768e8d8b9afaa619c0d87a4829521711ee625978f7b20a64e929452d4a562b2a196830bb592b71390da0927cf1676443a39f63b6136879e274ea3af0f3257e47a1068c2f549d950a401890a6d0b705d6995466fccbb7093953ab680c52c89e9e249cbd1ad6e49c9ff14c9e6273f1acee27fe7443294679b40eccf7a0d0fc5116a427be55136ff45ff5f9fa09f4bd2eb9a7c24510969d3aee3f3cc4824a4a886b09b85a2e0497c161f42b218530b8da594125dd78de14e105a0166607cc2141783cff1c5fa79c6d973ad6499b85131ea57480c483b8dbf5d1ad33f4723c85e61c97e05f9571d3fdcf3a355e6ba5d2545a4ed1b195fcd77a4044614dda3e932f578141e15e599c0d242d1bb13827f5b5af5a47f8940d398a442248815052f5b03111c8e5309461f449676a07193253fdc2ae03c47691809a4387cfc69eaca00d163e168f8e5f3d4c045273bcffc7bc1102e1467fc67a3e8120d7046a528e4eeac3c5945db4b570f0239dc036e883799c95075718a4b7b6c7b3d20d82c05b413f84fa347cf6a0bcd1368b91137688e3bd21e26fa3885d7743bb26a3749f57750336cba2d5b9c7bd6d30a7b2071597cfbd482ebe9a69c0ba21aae6fc2cbb403ed081c0fb247f8094a890c823ff723cd0719e7184a3fcb4f4cecdfdd5456b30aac6249b39acecc5b2ebfa632f79a66330ff91f9c4d2ed92d80de634e6b685dedd7b893110ea7b6e3bb98c4d7da7d696ae16625c380b84e14ec8788afda630d0e797c13046d22ae37f9e06dc39b73a038783c00b5b370f783994c82173dd50301e02351522cb1a341d63e708b41d6cc078ca90083b4f1af8eb937e757e196cd8a76412564aaa944f9598e932b1e75cf456b3b2038b5cc4d3514831c61336aeb2ba4a77ce2ebc98a7ce2651d82ef27c9f08962daf55061e27cba1a89c92331441189005143c7d197308500a4fc56a78c68b048fb0dc0ad1c372860254e1cfcdedb7db2a838bfb2eb7858e86789964b474a2ca1995f00a259753b485b48cb720835638b00fb60afe1d5ae1a1e8c3ba8def5bd586cd453b82acb2c58ed07d96382daccb1c6da22bd379c16fb2a4fb38390a17d3888d5c415ba41951a34dd20e05d78d9de69071de251ba9dda1c967dcc6d56c48745db992da1d87f83affa84fe04aad494d3f97caa5df1533c7007b4add4d1e2f282a7316a4e7586058f3141876e885319871e76bda4c3f4500d1f4212a6d0fb02f9aad2e0fe42705e7c6206d584e7a0ec08b0d6dfc3269b7e88c1c72c5de5b6428d47f24558ce4341c0a84515e3be7f72c8ad92d8b04dfde841511c1db933a878829d1ef11a34d847cb5d05e8070046905cd517569dabd9270b3d8620cad8eba664073751612066aa4d99d11761bb5c8137465e574521fc4b1406c028664dfba9333c6db3eed1af046fa3f6996574629d77ed1a097f2a44692e726849bb89e7f668b40a3e575fcdabd2f5260a0d911bf5caa07c2179e7eace7d7ccdbfd7d69383f02e41c521d9d34ab0f8d065607034afb3691616c3e2386285729b2927c9366e9b70062a60a315705025274b456e03a629c145a801917df69b3be839641538931fb9589f7095c9c538c4bc87d83cc1a8c21ae064000c2434cdb68be4800815fad87ab441b6a10330e01f2878d57045597305d68e36c7f0813263e3dbefb456773b808d14a83a59a958dc6dd1068ff133b8382a1a060e0ee1b6d122e285be987bb9446a7f9b0324b1a18132e2432ab9bf7e47eaeeb22c5e03ad27b09e13223fc6f6fe52352692a6c7d5c807c63450d380e87e434410a7f297a624adb4906ef562998360165a92486acc999e7df4824de1022983ad93c7a892557f32907f2f174f786ea56d6eedee4b2b43bf5d8c2a404e4591f2d3f52a39a84d1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hdb6ce5a7d7a1e22f204298a7efe2a4938b17cd73c482ccedb28015b26b0219bc78d04facfe0e3eecd6c3126365837447095c77095a28d70104ae18fe8e3535f1811baa3e75d3350d9af77ca31a1ee7afd8287b04cc29cf75f084caa958c2a69aa52b1a0fb08a41cdb1d485cb5ece7d410eac2378f7e9d4bff08ff2c774c260f84f26ae7887bdd1465f19466d817a3e28d372471402107e71e28346007478360bf1d9b34be0456f3e1e613d766f6250747ba860f69de653821c183d586d76d237e6ec906a07caac92d49d6ef501d0ff2c82cdc1760c2259af7f93a9ce698feadc6e6f00084493a6364632eb21696ddae324f04c06a6cce06f9e4debe788b4dd7bcde0a286754e2da6b88f7fd597a10a33ad1ea5d669ca35e744c60fa4b9f9bc8dd49195214b5542b179c5f6e9eea27b3b1605dfa9e19331af09d0d83566d2febae41b982939689368a33cf51d2372edc8b783631fc4b1ba8f9cfbb93aba70bf1e698d61c34af1d7def702ebc10b2f36c004888711f631d720787ed0d0d264edd12467617dbd09a9bdf6b84a076a76d2d739eeae5c3b75cc06acdedf58d58d4a361b3b342af8416d0842a4b36342131eccce94f39a141f4a3959bc5e50decd185e35458c6c6a3b8e0866a9c3a9ee5bfebaa211e5a6a06c1874c5d7e0f573434c898de9cb9b848af7f2f62b26c64d05335ef8e7dcfc93a811d41547030cb8c8b52eba0df052d4f6e18d5f3d199d01347b5c419c20a080430c16c2c0593a5c486814abe7664fac10d8516f8bee6a7ffdfb08a9c161ac80327b439d5d3f4c196b18fbb584f88959e967a95200d112b17222d2e85fd21f09e555757a203cef62a547a01f165cd4e3120a0ce191828df170dc3b46ec04e14ef85c6786c16794244413b94d62cdfdbd259a6e0fcf5a59b1b19df7a9464c2109eaa4a2e6733701bc3f1d125bdfacd220041744486a96f38464221fca9e6aaed8f0c38f9d28c6ac3ff8382dec17b14333c1d4867e3883f42019b4ce9fc754413af075a4ebe78e9c59f293f576d5f325c1fd376f1c7f3dcd52658ef05d3c82e4e9c1fa0e5b45ddaec8f20bd6184338ce2d0c9aa8cec70be1c90eb950bfcebcaf2c0b17d3205f60c1a1bc6bc3d1c57fc6a71583f69965f358628a69b3518259be87d93a3bc3ecef9212da1c4959374c30e9a176e9435cfd357e7f86c71f1ad1f5c0dd69ac533fd2d8f5474a61c29faa192e9abaeedea4d36d1250e7db5664b57f3dd36024ce55965ac7b2d66baeef798352cdf480891ba817af0b4d9c974cafc01ddfa09fb3217a314fcc68e573aedc38ef94fca5eda05170f65eff6aef0cbf2428bd4dbf626b5be4e2a39d337982d4a867590cbd19f9b7df553d59b861741fb994dd9ef8ff361bb17701ce6645d0a34d4bf877190dd8c8085e98a6bf63ed7e0054a77b3b420615c7e0f4c65b437485f28a80bba0b18c8beaceab288b278cad0c085a06fbc7e2e3572c5306d84787c0278326d0036b96729640f73eab59c57812fe7a0e58442663efbf29a7f1f20589bd341db681fd47c59129d11edbd8a1b4c496cc183ac245ae14cc230f5481679e54343b10eb33be8e64be840931b83729d4ecc172f9c129d65e66bd6ad840ec5c2af0e3887e7597832a45a3991929763463c225067adb451ab065aa040af41b79b9949625223cdbf352295f6617ff7bffe473f6128a15772293473a3fe82bd4f6457208c917d3142bbbaad1484397ac7ed6097e04988fd9e5450dc3392f54cd4aca0862f88958cbf0fb7f26f72dc234cda5773a552703e5051100efa8ae541ce260791909cdc57d2676908e66692f8dcba6b6f1b7f39cc3454a2216f8bb0ee40c259e6d7bcbd120d1deeae592d8ab2e320592dfd3629977adb2664acd18e6be5366eb420107cbd021f0aa6782480f12ccb962163794c9ad669c030d6f37a9eed4330768f5a3d3ce3f25fada9de648079fe5eb553ac8e207af31354821db4b7175bbd23aa8cb849ea99db3986ed750544a1fafeb5367366a9a57e7e6910350047ec0a825ee6004f6e88a2b1cef8b42fbbe17f87285cfc36c9a930872c3e506d803a1085ce8b6f2b19d0991191f7aabe436242859e2868a0d8b29c7a42bd7f8fed9677d00c755cfc54f259456b322420ab421e37c190cc920e74bd287cc8d527e38c4ecd40fa81f38c4f2174636adacdfeb549bdd5c6a7731d864e954dfcc4b85a69d8cd8288e1c5d95f138ff40f085dfc2d259d4686df8cfc710b6238c46d796361b0e88e25163da5a337a81a39db7aa02b21b00fcdda04618d13c369edff7fabc7100a9fda622b3836ae5139193a28a6d99569defcecc11a7c7bef72815075e60f945c45f62ea4822ca649d7e1707c4de57abdc1793fa5d1dc8ee5e29b492ce62679471d54ccd7031b1370270253d1df23cbb040101d8001523688aa4a56f02cbb51997376c9f023032298111f654c015bc07ab43e13a0ee4630f03ce12d315dde7a2d0fef16b773e597b45036618b76be8cbe154ffc088404aa5cdbc38ecfa8343f54518e314aa4e29f793670b09d9191d56fded93870c2f3871a6c6857caf8006968d3d70cdbd734c380f4264943eef352b3923b616df0286a56087fe7ced0a246231b12cc5d8040f86e56c9e335238ca3d2f5b5784207a07dbcbb2e29af45fee038023cf28778d3ad205bd358460eb596eff1a3504deead6b7a11aac642461e848b7e38a98c4cea03364c7c593866e718d7d86e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h849426b19ed2a1cba09d54f818839b5756174789640acd21c55dc7cd017baf1536489e5712702b98a82beea876f6de00f834ac0574a5e1dc11cf7efdaaf342063e6b0edc2eab219deb198238b54023b2daae3b59f14b2b3425611a3f790d3afbdb0eee6d6b944b314035c9f7c1e70e48f00efd14255fbc52ead1027db6e777affa502b6c2494c960a17f4be941bc548acf70d4ddca05975135d800b860445e087802af482b8b3c24664cc7468146c186089c53f89a91fe385635a8b25bc26c8b8a1f2618b2682f37bfe9be572820aa8a3b0b062b8ac3eb1668407dd925ba56f6a7d91962c4dbc15c6482bb5578d672ad25e48bbde952438cf925bacfede9a57e68fa3d167b32d8d9019f1dee528060925045d2c2ef0e149eea97ab606ce3d617e6db6a9615f5d84fa1bcf0f44375ffefa2d363e105dffe3ec44a0c09cfba9823422bfa248676b203fabf9727cf88486383250c0727e7bfa3a600db10c90cf32bcd56d2414844f567aded9817a21dba713d722f1297636dc0dfdf04f75af5ff5a7c7b0b12e46c2791ea12f3c15f59008fda12e976aed858e9c7bf8bdc1da3e90c5214c908629680131b34bc7e17e0cfd5b2ff059fee83f08f0e83a84b0f4426d9021b3b0e3a8491ddc07475556f2e022c07be54adb126f50f81f949edfa8eb61c553e87147a1dbda67a5382244ad799e41f886544bc0234bf990916f251508ea7d69bd2a1afa05294a1012fc2897cd5c0aef769d42eef700f1b84e0d1655fad031306a34d0f59df3c156a4f82ee58b28ff5e4ebaa95756f558c8d96139408c3ea8e21410fc6205f12328bcc1e8a0ecdf446a8aa925e74ec2c6dde24d51d76a8a3395e88c9298921b409075e5ad3c73e13a1f00f7dd2eef8c22a062b198a6df6c8907cbe4bbd01311c0fb1335f50ceb1b4b58b00b237080f0bb8de2700a30ae3400ed88d354aaeb140ccee76b58f6819afb4eb1c5dc1c8781eb9fe8f4d18121915a75d43c0240cd80fbf98cf2203ff3339d124b8e5d762b1aac7ebd0fe696d49a34132b96ba3b4975a4f3a6a06c3888a488ed4a3d72cbeea185e6382e9eeea4d508c50b9b62cdeb348e7d44e37c8644addb35810fde0e0b765d0a8fc124f1f2da8d1bbc1bf399643c0cc5adbb4ac813cf4504efade875ea528fae796c853fa3c1edd68062db31efa71c4b34d2804c2dd636edc0cfc2a12fea1a3480ef2609c8984cc4591609923e3d3ce3d38822a968c194f2d4d7ab1fd229dbd57a0f91c1351016360dc2d9a79b1887cfc40da7b1747c386607e44c04703434eb7b428424f47381ad88ef2623a93904a6c3ac07e1d4bffb26f3aff19f011de502b243903a966e6ecd1f80ed411b230acab8c54056e49d5f20dea993544a5d20f9944f7790398d6ea095e485a8f7a9f9482f185682ca4b7a2e01f768ea7eb4fa47b8b225bae2d8d6036ca64db4f8c145cf2242df39b08055a8da804365de15c0850d3bbbfb5c4a8e6b67f2d659ac892e74be5abb87d9ebd7914d938efa962cb01500fe738d38a336ff7baed327752d0a82c87bd15ec07e5d90d272f89b7cf6066bf9910a7dd230b8dc1c220d6121f7b5baef84fd1987b54ac1dcb5817672f84b8af63fa7a3955ad1e6e3122437ac0fae3893b79b067e32ae0ce07ffae0dbccae7dec4449263b124c4c1c2cb1edc54cfad61f7c8d5c7f62f5e80b9db4ec7101243e46767c325e90c12cf13f702a72e3024128018f6b337ddb49bb61caa73153fa3c15316ab466fec1e985254dff49303c604c2ea242a984bee4e003c64de5b33a04d1c4a5c3d83c1fd14dca9cd73b7605344853d087062b9aa96078f3c432210407cae3174dd9976a5354893a3c0bbb5973e5da6e25fb07e2e6a6159c35fcfbdcd9e97b8a97c798d05a646613595a9b0ae125b963fcf4127119e25616ce7664e51c1e412dea3181e3b34b14bcd3309fcca87dcad84fd903362e86252dc95b8110a106c0598070f108f11f60491bea1015555ad09a406822c5664f14980042f7ad967a644fac82663f12b2e9d82e91330fcbd63a684291118ad0c4bea47d44304454ece94bc3ad4e2b33138406fac60d98c019b8fefb672659d094b233d9c8e5e70e7114f20176491542e1a1e5577dcf5a1fa96b267b94871798e2b5fb83f8cf338a8fcb06e8c2e3de49072e4ab21706969ad4dc1298c3fa8080ce8d59667f21802f3031b335518d1a8bbc7555694fef537c30da8bbab2778d5b7b90cb4b4efd530ea4fbd8a3a5337b001a38652d98f54b4b34f9b700d85a8fdab976e7ef2c915fae7400d379b62971eda6ab9ec2120f8259d8b95e6ca47af6a506e26df9cadfb111f8f4838ac8a629322ec516b49f757611c1b32d68218852df6092a1f96b225d5bb74937b341f01608dec9df7d869f9adfa5fd45fc9124ea9d02ffa612c6d22ff34e8316b60eeeb1ccbf00593443b1bb453cf0e8c2d7d58f586adabfb34e7ebb7942157b04484a84dad4200df406361f41abaa14bbc7aedbd8595981fac643b1bc9585fa45558213cb7b8c131744c1e94a9ce9bb1c718edaedcb39c4258766898a85c8a2b978a2d1db03d17bc2bcdab017dbe014de9bff53a0ef88d4d3da286240958ad6eba16e4ae4d3930a877a67b9da394b20a8d337c7bb6d093a5f1d021dcb8197b4bc89e795b012f2367fe81e63764ab10a877b973de5791eea823d2336f9d34ac396fe164dc7e47f70674fc3c6f87c34287d134a3418a16309985e583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3fe681498a69f875d29acd749815cfecf728b4a4f3bdaacb78c9fc781bc89859f015997a0de95d6fff0bc4f4699086a4e2fffeeb23c7cd60d28d0c947a63aa27549a3492cb6e2591c19dbc5a10d6a42b2e5903127fe8c77f22bb533c25acf51a797beae328dd2cf48bc828357133e6d7a81f035b0588ae8f0dd30b922a35cf6aeb687f49a078fc52bf5de22334f7ad3b7387931c9ad28d3f50772df2fff595dd7c3f401e91b8c94b1ab6134d9b37fcd5fd13a8f1bf7524894f9a88736ca31bb357b1f9d5315bdf15886a95be587b7a63c429e91b278e888aa4892cfd9a4db65886804e7a5cc07704cc470b7a7da8db80bdd8b3bd4497c538575fbb3f6ebe8397f4d1bfc8ef0ec3b19da649bcfdaeb9372466a8b78b53add5f493c7e85b9e224124435271ade91c43c8706873db470c0438aba0a6a4bb35145d2a989163816c0bb8fe93207028e6bff00f9490f641edef7b7c4c87941a9486e974b896e5de2b7fb586d2d54413f714f5c67c2dcdfc986774942d0964b2ac566dbdddd16426f02c044c933f2b58d79e0fac2f21ecf8763c676b1c09bcfde2afeb39c03f262a2262d6fd35200a0a06ce11cfea1be99f01f74720242b0f0130351bf6314763877cbf28eaeff7304a23fc211c30aee4d042ac7ab4fffd08000e6db89f34ad7bc2a3cd0864ae749f285a16696099e06bf987f4e531551bf35ac6d74ff7228182ef78f6a7e5b26df05d9caaaaea2d97ccb8a0dc0d58f9111527db02b879180d0bb8df253935952daacb8353b5f9e76ad7476971c625d19380fe8c2f348d606c391be45db3ca4aadd514e252e5ec9f2f4941ac21d75d0bd1483a7b6a124a33cd0a17d08f90a587999d379c19f19c9a53cb04b3612770fd095d9ee122c552618789b7e49c2511f63e4a596b3515f50a4fc94bb31995217fb46bfd33393fe66c805b1ec0a630284537dabd7bcd7dd45d52b52257eb1f90b8dc747a1fa9b3f2eced140daf9577bec0f1291d29994cc19499aac96bb67a8bfde8080eac56438c0119d1815d07be571a59785f3d95b552b768f9f72c201045619fffcea58ea23c41dbc76ae0df6097039cd4dcb54d561b455c651c673d7ab677b16159dc30de76f70754c26377c4b2279d1f39b9bd33c039f2ac5cd4aad694508e5869e3983c84dfe8ad7d4b0f08bb4e565c60ec2a941760027344f297eb8f21fd621815bafc418efbf788e45bae020301ca3c077302dc24c75e6c5a25eb569140e881cd0808ab2007a198709562b206af6d9658617f8cf4b6fb896a73c700ecf5a51653d9619430642a3071951f41f19492643c0c71c3edffcdbcb9caa945a6c4a6c31dd7a5ffa1198e2b472b912788159287ccc756f6d4f2a3081e975aff672994ce60a1cc688b8bc924fdd3c363e6db0d82f0ebe5d587e79df6fab1c0219b8211501f45c5d706d466811c46943808196f1bdd0bc93b2d0b6df148931e97f7b7c8dfc5e69d9aa5ead9815b66f828ceb8a8abe62846a8d6e2ef48809a5e9cf91ac09da8d7fea429747581dee8ee20d1a831fb4d2aa9d8c50cf16984e0830e937e030f036a66a34f8d168c42db459dfc772a557724cf7424d8aa54e1553f994f85c77cdc6ce6de36a6071666585236471675232b515f932277ad4f040b24f7912413f2c405b0ed80568ee459a3b75be17126211dfababe7b15c242b0eae4e7aa4b34b4f922503f7c7f43128d9d497724edaf60549a40d39eb6c70b9ab450639d474737e18804e6811bdfc0e419ef0a7092fc25db74e13efef03c8b08968552d34cd396a49b87e18739f2d71be56636db78bf6d1f4c76ee6e46564f564449566db614f577e475675533aae329d641a468d94ae6800a78276e1335f2c9dae659fc145b322b01735bd835eeb9b5ba236c0909d8e96aa72edf31b9c71f649ea147a8e4b1b67e30af48c85076638553e378daea3e5debb1ec51beb7a33b3a8e234a364c88b922a02374bcc09dd31b98d80e8eeeefbcfe50c6bb909f3a2edef849639961fa8b6986af83e2d95e4a90db399ae8c13c56e1d70ef16b154ffa011d74995301ddde0cb51b0544ff7e5731809323da29f39dd3b47d13a531e205da0ca9ff941adf5aaca19a7c6ddb296e733fd63ee3dcb9764f692b3ae542a978a86ecf83321cbf7999e4d8104809077696de256ffdab9fdd8764191911e08e226596d35ce2c32ce187465d4f84e0bad1433a1786ea69deb4fa9bf1e5e63d6816e1893a48d21ff01239fc1b00fd7a094a8d9f275983e7d90da14f716217ef62caaf877de2a1c50e9690c963761c32591120c3844b2004eb4719f9e920effc555a1d462b28d92c3db14f4d6da66d35fd27e899d7b551c19c15c0d78cd3dc1e633ebffab2faed3339142766446fba28c95ec5e9ba8a6f4ee99f1bc50f68ec86956e37bc2ba804bf7390a1dddc7d333b533a078c9ef2d616bdbd94d93b20245a899c54c2fcdf34e0bd685bf9014251d7bd221701f8dbb72d9d2ca3ce3f97dad5725b15287bfe77e60cdb5791f60a71abf6082cef57af5ba6cf6407c9323e69bf8ab6f44808b21c7709c6039420252350edb52dd5eb73ff2accb95960ef3de2b3c7549d92704c081fbab73e14351b9dc0a889320501ffc0e005af83ca1bf4e17ad0c4f7ba8a85846fcc7540036daabbfd5ec43b5f6a73402ed061bf0e9733b95feb9c893d12ac373c3a3801d9d833678b5fb1295c344ee8143c261ca180a0b483c91b52ce9cd3b13509d33e6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h244d8fc9c31451132ebc55f9c18ba1c7d740799b2e4dbee3ce3817f5aa9396f816c702eb0aa9a241f792d6adae7e902172cb25e3bd67d5a233504b695759cbce515f006b485d1b574bf6253977d1e24d73d03c3edee9fd71f4c45f99e9c77716c7d129e04ea0605e4537ad6c681abb02af89f5ec56df995c803a7ce46f708ab279f6a3061fe97ba08a91159fef0cc8de9157ea89e15e0d79e0653a368359388b551002fa8783a7efce33cbb869113c692414da0ba226f87983399d5e2f937113b4e1cdc9ee6506f995dc4ab40f3d6eb73978388caa7076f170bc3753e5fc525a5e8ee988615e901df3667d6a02024cae31f7e501ca41ad1d03068929a909d9a35ecee5b0dd60281114e8f174760e18c747d1c6917bb22e7abe7a255c3f52a021961deacdac127b0df0ba46904e8887739429132dc9c0f0e724f37592f9579e4c83c33e04422d684d909af6d9df645d592cda0f2d6e2627d493190e3f0cfcd4b0460da947fe64a0c7ef67e2e827d28972065f6e160f5a20cf752fe5fdb5dea2a43aabf6132d45a892868beb5923b38c986fa80aa5e1d72206a5469d0fcbea55d29d0debf3caf9fa3191d6d2f50fa97eeb91997289004a4226118827662981412662cd05e91505661530c6a977c0847493ac7db86046bb87cbc152beac75f6c1932cd913d00335958b4bf225f712b6a832dbde43561a68652732cf6e53eb1e09276ae0d375e3555c916c3a046a10599fda0c67b7f18515f20052169774c718578bcc2a1e83f888008a058769aa179ca50ccc713aa5566a91cd092a9ff13983d32211f2bb1589c3519479dee4e572356805cc0a293b90d8160e214795a028894454391bbcf0889e1aa156662e1cb9406937ad988f1e78374ef30c8dcfe198325842b34a90973ac35166ae4040f373cca8f1d2e18a413ef1168b3226dc08d4993c8bc322886b134d54b9892bfaddfab5bebdaa21b34d0bb2c20c7cc90a5115f386961c50ccd0ec5b4a318bfbc714ac5f4b467685eabeb04e270db09592bea900578b695fa32d12fbbdec5eeb53f83dffedf254d357b43466e37d74542b16189427955cad9d78b10db00b07e87d8059f7565f571a8476d91a65a4141145509719b78eb4afa473278b2e69c193d33f72a06e294cce7c2d33f5f7b10435a5654e9d3e5d130d7047a7d4d8e440da32eafef4f7ec97fbb9c70172f456fdd21643cd811cbdf7aed87cf5d262b2733662d7cda25cb177dd77e4df0ab7f1af3b7dc6213d93c89733944c924f790cc3f0309240a1b6e6384cf42650fd759c62d3df2069db4ee90e7e95fbf897299c16d9da96b87744df51f25359213492cb3fb47e0e358234f158b841a66efb64b2ee8693a3d9f5d5358778fc8fd268f01541e723d60b717097cfad5334199d514b8fc53301c8b65d68c5f7035a9203daac1e994d3265710a5ac1546d7c6e1f8f3afcd6aebafbf5a947a54053e8dd710e494be7b7bd4ba913a21da8203e6ab69140daf7e43212151d32c02f22ee3ff79df2cf037451d18558079d6cd9916aee7f7357d9bdd8972a3b62d6ffd673592e0b891839f83473ca5eaee5ad112043a6ac0d7838ca303c1b01b5fe9b3157909d4f28782c0420b75aa8bfd11bcd5ed6cba2a03e3dc3008a1283ae9b51445dd2d9be0c132288dcbb82c183b0dc64e939128f8a6bdc652b3e490d3763a3750fcd4356cb98996f957778c22c9391ce0943d7e86e6551c1ce773c4383edf1040f1baa1ca3239816ff11a72e2ee158f88f8c294f0c8001125b562d38d0abdad9d83a782dfea3e2abcbba939d0f4e10bfcbf32015c6dc1db8009bd5b2579e5295d0f2bf83b27b6f33cd3d2d8ea7fa3810ac6fc2c638a85ca52211cd7b0f9a5b98636bc8a931a34532b9952df5f2297c1868c9e0cf66a807776dcedfed49d7c23c78b7c3a90af6c2b60a1bede18c5081968b79572f81df6a1d5ee275663b6fc2ea8a86893532796d8922e9d626d043901573f3b2222c5ce63f788f0de507c658bbbe8ab4ffee898d730a778f0bb2a5cdb249a55a5df738189ec5ae6d621805d356e538846e0491567fe540dca7b8844879a23c943ff11e82c52fc111097f1c243dffbf173761c5e4b0bf288c1ccf4852e7f67289296446853feb09783fced1d0d9dfd6f780ad60318635df3dad2cf50370cac5f6c52adcab4f3e2608f3ccfb30177bf7150ffc922e232292de0cb603403025cc21a9d978dd95482fcdc429074f9ad3b1eedca9279820fa2ecf943b057ac2a0d37dcfadf1a896a4fa4a7b34e88c23427b3062e43cfb07b970961bbc74d68238c52a048563972c382bce297a1a2a21c4dcfa51c7d98458c7546fea7d98a41a0efcfbb18ad064b551fe9b0701d27ce6e3d734e18a8fa14433e3f9e4a7a19830a0c8dfb766a3a6500e994f520176e43f840827e7acd9bdba17d03a365ba09a17909604842f995617fdeac0a47d8d3b18e1c50a5c634ca431e5c619417cba0729f9c3b5b9e7c51b5875d0246164f1d245605e752b9a3e381565a67872f5df7352ee1da85c740f312d6ab8d30f84db39492125066c95a12464632181d4697e852f30e149c21185a5e24e20c32ca922be0eb75fef963cf1be6c5f33807f0a673117aa9f63b48f7748c81492c803b883ffa4e400558080f62f440a840ee0956fc049ec8f036b7383aa6eae09ae3c3870a08ff8aead12d9129f2271397ad6724cd1f3a94a89fda699e8595709ab55cc65579837b8db166f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc6a8c9169c44c5575b2368185dd953e4c4bbf0c4102c9640d9eabaa5bef82aa559216c6aaf4bc9052ebbe71fb2ef1a76fb8d638544aa926b7700f59a19f66538e45701d660e52e690d6999f2ea665c7d4e98bbfdf8d0d2f2fdf5a174f3f39ebc8389875f475f2eb6747b28caffdfc665a615bf9f8d1d5a91c58e82532ac18867d65df99982f39537a304f7c92486144c5da852aaed542f59074e4d570b954cb494c237b3851fbafeae7dfc0c3f9c358018a3dea34d2b444cfba6caf9cd50f5ef5b17ab3e347166161031ca2043c78cd2abf03300025bf356123bfc45e46ea27ba07b2e6a7cddf09577b3199b46c87b0563d9c0306247aeef4e03d9675b8efea740c776ab69a9a698d143d6499a870c4e7fe6cdaf2ff39f4888ca517cdc0a2ac7279604cfc7a609387cc0f8c55e82932efa5ff18f7ecba00f052b702c43773d859f5a4225917b3906ab87e40710fa2eff662da3107552f2ee32c76f4d4f1915c65bc6e8a2e1a01699276a9fc4bceca29a93ec0f0f4dc2db44680533dcc2a95ced3658232338f720ce998545c27e13c506f45765af9f5341ccd9be1376d9b93b35002e25f5298ac0ceb74a62c5d74f8babafc699817b242be5abefad2b6db18abe959a852a97f344c363795927fd7d764f349f465484f5c8faef145f1df17066b7cce77e6c756d595f2ba982e2714760546833310dddca5b76c970ec9a587a2bf7add163f6f58e3660f540a4703fa4777af1e3bafe797994539a5fd4ca2186266be21f18e057603bf6fbace7fde5ee7e96d9f219355a4f08d2ec1c0c497abfdb6fd4beec263f820fbfde9898d3d993ae0e7243031d22b70d7414f9cda2ac8fcf6499b581394211a0f8d9df1561f87e9093d68f7d2bce75d5a614bf0f51920de9106beb832d2fad34bc0eeb5820c514485dc2be9840793dafe6632e335cac775937157b482c69433ffc655e354f9f154cbddfa201fb5f1f002260274a48da4b55b87fd18d65a5539296d92027c3766ce861d7daff2dbccf2453b9fa6cf3e2947c3ee258cb24eeb3f17d67b576c393c7b95557367bfbfd183287d40814ed803a8f1ca53640cdfbd83a77b0ee0f4318d847e487c022284e9867dcb3fa4027bb5a00369d7bfd8b043619d85d21f1ffa21e6c50228305992439b78747bbf8eeae730b076c89d18849a88bd0d219b40cbb1dfee8b69af4c1147e67da5af782857e138615fab457f4f22937ce94a7ff31f26b70b2b56b726cf0038ccca845b71513abcb1786b25b56a17405331672e948c7b627d4b832b19436cf3850370fa657aecaace53a2563d4e5e375596a92cf2ae4ca4e8dc86be015d138ed19dc1fb01521b0ac3273c058a4b71a05c9ce5636c28d13376165738af0336b2151123282d4a03786ecdb7216868db15d2af90203da0260c4b27a2025004b67c6be1ff8f313f98810116007524d450563e5653d8727c89ab5db778d6f09ad9687b189942fdcab0ca212304f2a93b3a77aec746dd6ae082ef3e3594b540da9e46fb256feffbceb2352a505963e0d51b6d4c99f0263e08d8c210d679f0199bcc3ae404a623676857d1b40dbd8189103e817eaa5f242b3525f5492120626a604803e21b4240688652a830f673e4a44c9818ae2ada4eb0fea5499351d366d4a75e93e97b7c6b392e3d75f04136ff3e5d46f26bfec7ddf10e8d22c16eb49f40670b8da1049354942f8c469d6ece7899cd208553d162ae5b8d9f902b6e5b32919550ef8ea3aa7476d9b4c82d789a289997ae458a5e7b65dc0c957b572083d66a839832a3582c1d71c28d188229acae37dbe6972311ad82fe0149c44365ce168581573651eb80a58b0a6e2d376dec57fe87043291d45ce4d7f384b1db10af17e50c31da0e01245c0524f73fd6293e1035029198bebe0783f6522ffbc6f06d291a9df49c73431669c063dfd868ffda000cee446c44014e20c4548fa8f55267a33f6f5ccbea29b10c3379fdd5ddb560682da4b9ea52910b08451c8d05fac32cf689d5f25deee20eeeaefc0ddb2ad2a55198a8c37d6b5762b1450d40b94c30d6755d00afa6e68790e34cde9604f955ff4482f1af315f0c6533811ba4a185729dbd18c278d0474a3c3fb0494884b9741ea3e0dea34cbde5a09d8dc083f8ded89c5afcc18a4227ed873cc57436124cbadc45eaeca873578c9497b5e7bda58a2d7c9ff7466bbb2c03a5ebd3b87723a4344b70c622f08175156a7cd460e48e4392ec1568b03449b2410b3543966979fcbdaad2772fc4ed70d9c1a638e2c62f7c8bb058d56f55d7a8265f57a395415197de212a6d0f899985c0317c8a279850a69769d28edd3f3d862dd7f5ba974423d28b1213191d028e84eb50616ef6a286dcc302453b61981e5888f02ba8ea237ab1fbd996bb9bde8c291755750559ee842df39d138c218242b5529b8a208b2b5bab76e07fe5322ca9115d7aaa2739e14ea01e2bb3e16e2ce350a7c30ff60d7777b641c89fd53709ef3eb556cadf016feec88204d706745b4565ecfd5e66449446c8d5c8d678dbe72f835d8216d0538dd6847342e1459860d427c6a11d327620a62b6fea43f3b90c3a608e79581fc648bd9504dad39de5a6e9af354ee242bcd246beed9edf98c0de4fb95002a935d78da93dd17187f7f1acbc58d6ca99102d76bebe399f59432149e1fc09581db14ca396502f74e8d724d784ae6271430e2b8d63f8a8c9310e395d4868a4992d08a90e6c80493c188214f50ab52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6eb712ffad171cd776a33f508eac19e19586b2b726fdda6f456c59110618623428b5e96c1f939007e35646bc1783e64112a4a72a7ab1ec822f4d3a561020361013016e87d4ee1779ed6aa00c13006ffcf26e1a7db188e3714173a0f9c0b4bc63060e7daada68933f8e91a13d3fd10d2ed385f8590b0072a70e8e8fbb7c4c04ee866857fdd20120fed8c0d6c0fd63257e3de17bdd47efde0f32f0a35194ba52a046ab93d174028b0109bf8b5e48bdcd089c472f04df5138610a59bb259f5e34f32e5cf78f7d09c9c5db5a2d5edc4181913a8f4ec02f882fb5a80d259949e13e66c887ae828320e76a826cdbb2578ebc30cf5bcfa887b426e5eef04e73fd3f90c6d496042a24ebbf8c71b4c19a94de556e8c671b2507791d73bd025f9639550c999292a0e298366ec6531df06eb62c87b021378c45e4d8d5ae93a7665c2e42f6d41c0b4d4723ae15c1780ad35d01f71b8473b7bdf22047695c746c978415fd5e85c034d0e1c9ccf650bb8fbb5d04ae8e117c42bb38737022e2e20d26629f6f231b5922c15b8945528171232080cb28fa44a3253a3bbebc5ea9497e91dd0f08de0185cfc0e08bedfe4371d8df93c8a6bb9a182e3446938bd518564d3cf85e454bfdbd37cc7efef6a4fd7909ecc26c811f4917c1c2a37ed7befe071881751cc2c28be355d1ad4014696534e7893f4a3cff7a8bed914d14ac7fb43750c371fc911bbdedc7e0297256b4f3c0040c18ac24260b1c8e4429b69b2cfd1906a8d080805e9d6ad011eb73d44627e4715ff59736e624064575ed358e3144748b1fbc22c6a02aceb3e5735fc9b4388bcea5f90e11231ebc15a7154472fd74b35353a7ea7e0c486c1c82a8527c6bbc65953bf795e586d74436d4d1b70e85ee4f835dab164a3fe072ce1664129c7678c73d161752b8aaab3254c177eae2cad46dad3c49b3caa404a05a95dd67c7c4e85ef08bce502f560f0a4ca5706b116880dea62324beca59d29048b48fb437065f0d015b053c21384418a04efb6941fa3001fba0c17b5ab4ab4d7907e6f637cf2f778843615087512c1488b622683b067e61f28e213514cfb277b4dc4ad4caa23add846fb2beded8ff1cc8e1641350c0fc376ce9823fb0b6391f945a14ce2aae18ca8417279061d6ffb829bd5d1f4918135e92e8b957d70721461d7455198ac892c4ca7fd972bac46270a4d99432f0012b401efb953bc1bb82765fccd45b51ea1722c9e62adf0ad03a90bd4c33384125b5ab6044a3f99907bbd0b0276d8a3eb0fd8c8945e120fe7dd758ec3f3ec795ef5ffa75ab28337a29a56ddfa28e572317a52e502f8ff740d25535107a016f2d4f58093fe01249267f4c914e00d10ba1276a6f113f7678fef2d2b2cbcbce46df8ba31e3bcfbdda8b9400ded6277bfa7cc3cc5773eed2d83cd30d6be95534019d9efa9eda88a99d8e73254996f296796117021c30782de70bb59c0919edeef3e1ce04f960188b2073963957c108b623fceb3b6ed8406407d09bce7feef1d2164fc4a747c7c8abaf7c526779bccc6abb82621ca8681fb3a33cc18eff51cd32ad441b874baed6f1f35c936654b1b29273685a77de85ddff76bed5cc06731177d608565e278ef45963879173f1ac1dde63bb4f0d9bbf735f81bce94ac0c04ae5577136b0882c65f979b0cc8c77f00b1c5bf207e39f1f64cfa49c60b48cbc4bb957d6c4d0475caf72c599a01d07c1180396ef745bda52961196572f3c8f2e3f0a1970f746f8588bfb8cd56031f1406132526d1186cc2807078583c071ea35b1995dae14f61b7e7bf054c59ad53560241e051daf6cb0ff1e94b73f393202a12b61993cc489fe2f545386f1fb89294f623e0695052e1cbd9d43c8ad31db5eb3fed32d26bfc7b429d2a20f06915a64dc3ec8d4f04b7ba24b6e873dd53da215e2e5d2797e9692d05e8fa294e39faf1685771925623f94a350c696745295031520393333c48a8a95fcd6348cdcc43d90f83dcb782b4f7acb8e931bba50468c829bd7cb4c25878ab02cf4b47de6c89ce48e9f14820c0e9a239afb2df306a563e219fe4f796852a31db1dc3242d2203e2dd47ea3124b2dfb01b8c57388930f41d6a60ca2e9ccd95ea4bf88f78458449ce920a9e06ffce44595506fe13f73ff766de6989be83e612e0fd7998b5266c58696449043720df0706c8a1ba1a91343c51f1a95cbfb6acac5cc865bfc2468c3dbc5cbaf81fe7cd4fa0c4e2c9f213fb0df25b6a96b0b19e22dfdebd71a8c9fe4f7d693ac3d6b56dbbad2dac49ddf807b8cf5c7e564dec4a1ebef7ba6c151c7e731498a8021b99a1c0f03c0bb4f8152d282db7922694fa30c40955af1da9bea724a1ccd6eab8b84762c4a3949d7294f8ed1577279123ef07869be84ccb1330cb8aacf30c37ed989f5d3be5999d53d54a9702baf1eef45ec4b8042820c2f2af5f4a422acd6995adc9445d9a8490f45b602ecf5902c3548b3f07092aa1f5a311bcccfdb8dfb952dc2cedb7f3c1eab0b3f39a8f4d83edb193340e3ffdb5f8b7b94182721b0ae9aea9a10b7d9a3ea78f5cfc27d1836d7ea8b62b476fc7bca56f2786bd62d90037c99018732ce6ca80f84d416ec5f4c1851ecdadaaf145b35f867a42a9876135f55a2535e33b6c2afe69cfbfc0e3140f0f224f50a69043b52929726492bb34f44650e7fd300e76f25b002d6aa1d259b239991c43af957db1397e9d164306cb4dcce6d6c84927ed003fdc01e2f93c314e65f44274ed6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc541effa5d2da3b6f6b310316770a513b72f4520a6f5c686e4756a239f1983c91593ad70e9d77f366a3e10b4642b5a1bf1f8b0907ed940ea56ede648535d198c838144bd037587377b3bbce75fc5cf4441ef00de11c67e3f4e35712793862db5f65e249a90a9338d6cae1abb13a0463cbcec35e1d7829ceb4ae3a0e48a9ac9d3949f4ecd2018f7b7c85c67412c6bb39810ed1e371042cc658bf7055ece01eab0a7f796d5c0063ad4e71601e30410345f29cc5647251952108fc16332646a70d2105020680a4a53eda1af8f4aa454b9acd07604502a864685e6ca668082dd00aac36dc755016ed917d9a76cc6ad11d36bace3b7573a2810a77fc84889c0a8f748fbacaab83b6959edbceb7bcb643fc0e0ad5a29ff2dc2cef09ef0bc095edb6fdb1d726cf02fb6c39d666e5c60487968badbcb254ce411f45b37d5425516ade948f22e647b9213ff3e22fa052962be3ef77d48ea9b03021124cc8b38dba306d8ee947681a60a410daaf088b1bae3256d0709987b084b23d19adf157fcaa2baeb563d9b6b0921984aef0a046867f59d609e664499378b5d3374c95c8b594590a1c5f86b94611092cf007131292adacb534b4b8d47b47d120c58a721693beb9d7969d3ef7db7d0136d837e0a00c4b06616a8c102c344eae170f17cc2fb80e53980752f84824128aac1ce13fa6cd06ed1240d6eccb5822dbad5c1f2972c5b0cf52686f4b0a4bf7c6e0ef9073152dea1abd46211f33576f34e9fe218819b3eb74b61b6e9c6e2d30881c4eb21455001cdf92f73719d9396a42e70dc4076b1e7de65697b778606bb858099cde673e4f9331f638eeeb6bf548627824d1d60f8f595ccdf0b75aae3b3b3bf96e3a82badff2029c87fa38c5a72a39e3cc98aa22bf3056d15e61140954235f62c573323e86c5e6ea94d112a83c227af857e0116977aa0463f6946eab6328199bd33af76f5c0c9c9920a413c8c971b7593b794437be82714a0b205a808b2479f5b9df0e40856cef6d9d50147ce106ad4345c827cf72da51b6ec502b6f6b5f188d4dbf10b04287af8b5e5fd36bb368487f79244d12843badd2584b03983f01e7950b310110164d8af190eaac5954c490c5f3abeb521ea2c51bd256322a41eb744c2333c976257759b19f072a69efb1ddd518c00e0e9bdf0973a3387fe54eacd8d2facd87fc77192315540918dce533eeeffa2c154a1fe37e92158ef1c35e1b2971f067ef139145cbcbbfd2cb424f5f36378418e76463ddd3c0fae6e73f94b0acf7fbd73fc70c92918c93575c337af0e390c5a6136beb111785605e080a4386d51c35f8408190dd203a7d6eec888128c77ebb3f838241337118e6f3cb6d31719f233b8ce62f4be130ba249194920a927706c0172e958dd28f81fb7c011db88dc44480a2327c7a8626f59b682d4973ef64929b6b2161a40fcd630e6cfb6b0a0cc0fa2d2dcac293c913654032d880505f31a3d9815b1a8739df2bac39460217a35ee03dbeac7a5ee0f5171fb9b813944388c7118ed335e0391dfba9fcb260b5cc76a97331a6b4dbb924e3d8946a04e58ad3df165e2042e5282577656522ad560258bdc1f2d12038a2982d1f959af6deac75968d7aeb171c2f8db288338b13b0ee13111d22167dc223d7597414f3e234744c355b89847e4299cade85ba46695a4ac9f47c4f14be92cf8a6449d321fe740dfdd4603e7e4257e82dc4788b846b7684b2574c8feeccfa9608f2ba07a351073a27f03b9c3466e76261a85526d8e2ad211c63fda1b8c4476816906d9c48c8a87093f690304cd8a4a92be43253c08894e8f4330b009e57318a68a3a23cd6c4bf6cd9b6df7f28930b868859c45d5d93a3a326dd21d9b1611c503457932ec3a6a1821c2763143bde0133416bb1439ebeff51ec09831f1664975ee14842dadf25263d8f9bfc52c102c07a107a33a41f157fc8f732b0c444882ed53bd4595e133065b0ee804d4c49d117da6a3eaf8402f9dbed1f4a6aeb37b2dd0b2ae21b89efd0f8750aeceb64a0efb2d653e07649b98ea94c786c0417bc2cd30ee138c73b1e04d7aeac816af1ba1395c791508bef83a35dbe47221a75c56a64532912bc6d21c5b70d5def9bf4005c9cfc094625f34ae6505d7a7758ce26a1498505b845bc90cbb7065e52479d8a4da02fc384a6d613ece401b1f9f03f476de38dbc6fb99d929ef267e5f6a7c06c121e158b32580ce99afe46aa6e9b2c4c8511b1c1b2a7defe593d14ab99cf3dbbe4db5e30ec528695b35346798e4acc62e98a89d6752603de3aa4d9de94af151bc134b436cb91bbf492ec1d85692c5f9c8b7eed8e1b87def852fc9e60754cd22113520dba512d1899ef6e495f7220a1185026f1f73aba874a50a7f4b2ca2317049379d12cf4d212b752b30feccd3aa51a340bca18701330cef137604259cbffc1eb034b41de84cdeccfb1b6b9661b7dfdd37cc4f58771d46ceaa489d44df2ff00c4c1e1925494d7612697f4951e6c4ce24e919eab099a2704a75d3ab021d35ec369b6885aefeacf10194a6badf325c6965e313e50d5b55d7678775f7e773b0261c2c210e55e75729ffb14cb7097e34801c611c48f433331759e4ee40f7ddfea4122452b035632187099dc381580436377edecf774b439ddc6fadcf6c7823688c09585b6b50ddaf09f23894735ae343c086bc1181a5dc5170e1b78a661dfe8f8725a8358df473bda3376dd65053dc606090dadbd853eb76e96d278ee99c2c88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd9f48e120085b3ee81b3adf936dc7495ac6f07812e59b2fe3f761c6f7565cd34ab6c98403820230ad84c96ea24dec60b58254894fdce7fc64dbbf62629bd69cfc08ee8fff5cdd5dd3cbdb0fee32fac9a423db72b533128f7d0f4cc4ad4cad508224226e4895a4df3eb6a574a2b69b2c758e9f06660d0e6e0a1b490a68e23077f4ef8ba04126eb835bf4907e093e2ca2389c762127be03cc84431861b20f69f3498c75c1e3ac9ab3dfc30b05dc38dbdc69136432e00e02929ea6a80b67d4e04449b0b79e0d36e101c72ca2af66a5ff7e304448f13ea708910438d933cb6cd1d9ceb30c5edc507c20e81c3e5ee177e9da9bc1cb31d72ce5860d54ae229e971d59ec6a919ed75e114b9f8935b831f4c7ea43e4b05eb07e35ed6af039af9ec4410e5103893ccaa3d4ebca1c65273915c19185e67dd31fe0e30f77def4e2cfea5d829fbb09c33926b01518d7b123f6882e51b7110f64ed2032504886f7d9d80bf2ee04d5e2e018b08189a7841843a8767eb30ff2ffbb9cac71f3592af43da0ab3a53b44693d688806bcffa54319877c8550b8d8015dd37dd9eb8431beea209ade33ebc95cadce796b31e70c6bcb239998b52434e60aa2fed6752b68c502d5c35f234749e850d50b729e2c1d026a4e39fa156513a52df9ab1a1d5e3cf633ba6167fd37868c82438cadada92a165f8d9d7cfddb8e3c567478701eb23359884f29530d44b59858da698a1c77c3796130cada55efd980cbcf99dc5862b33002c9cfce6436df90403dfc3c41effa358553f7d777eca855cbc15d8ae1e5dbaef644627f64370c95e775c8f81e0eb8c7e96a6bca5a5579098cc793ef8af75a1c7c494969233c95d2b7845d83ee27e4a55e4a4b7abd6eb88114dfcf802f5e859e6f080caf35fca4d1a3a18d8e8c9f647f874639fe276a943cf06aeddc9da976b0379090040c730b6a6732c3e6f75194d072a84c58a741c553230529155c803666034ab0c6d59b6212d98be5f56aeb5a1544fcdeba0a5b1bbbd3981a9c8da61aee9dbe08db30528a1f3b987b7d437a21fa1d14597464e7c00dce8f1308194ce90196525fc5a55fd1eb0f2aea8bfcc1e9e11f12e52cad66cb9b481643e6501544a9f371ae2600797cc88ac6cb9e0817be1e0527a6c459b80afefb7b880a0f37a79df6b94eacc2d3c08a005d55ccf301dcca56c1d0ff747d2da29485108c7f274c18d7916abed564d38e1b2d01c8a441d61c6defd47919da16f4e195f9ae85ec60ec669a1e01502c19c0c0cb856b4ed4ac5ce1b50293e6362e0c8b610faf85177f8ccbb2f9080ee2855047502e6b7d58ca1a0ebca9d8a619be4cad38fcf870cd3ab5bfa58b6987fc0aa1121844d746fb58def637b5f9c28ecdda5c5a05cfdc310cd964fe78a4368a77795664addbb1fd286ca355b7d129dbf05c4425ee7ce56c75f3196cea4ccee7a193a62564f1f93e41c695b6ec26afdd7f65b535a564b12fccb11fc35c93293763ed925597bd4d7c328677831a31440b1a6994d2e5038078e1e3fb564776720b62c65ed85290ef3e59326de933c9d308a730a9d12f1308e6a21ce3d51d4f1556c4075fb3e24945e50644f1c2a833508cb323f5d2f715bab0578d880025d1fd8b6b398c40e2aabbea2de214085bc2b60da00c74ec4d8aece11b3c5a1c72c1a815ed4db9204b67ee98d884b4fde73b486e6e7d1864eb4c29e8cfae3307f3b854c98cb0b2e35264de6b63bc6011256f2448ff5b28fd8ea9645a65d54c1595e05c1191d375ecbe8785eea0c47bb0a1610c569ab7ae47ccb3006ecce1f29aa7e9a2e798e114d5e47b9af2b2cc4aa234bb495a23eb8cd38aeef98a2a4fa52d4b1862902d37247f3372bf9870931bfb25efc02bf7d585061f73930ec29d53c44ba84b2d31e221d6193a6d5ec667ff2b6a37af2a832a4acdcbe9f009d928ad702ca3eb0ddcdbf995d42ffffcefdb0feb9a91b3343fca48b40f806fd75ec29b302f256e0019320bd625374c4234694a451920c680c23b6da9b26113b8dedbc7c24b11b71556fcf2d1c46219ffc5bf4b6b0d2bbbe334d3d4d0651f051a0a87aaefb79009db179a4c35b92be9feca5665afdb96674e6529695f5f1ce56777acf05c978f16d72eea3cbbd23f122fc119ada20aad3e6f5f3090d586eb88c01424246513381cbb5c856867f58e21492443041d089d36db2dfa42e7f4059dcc72af508a2c9d84c6daf49f5955c7460806dc7463704a944c02744c7c87215f29837721631796c0b23f604fbb67ce41635ac6dbe15b11886291077fdcfa2a81bde315a4b50ff99bedb02003290632e036cb8843f0e52022bd18f7730b211aa446955d84f9df71cb119aacc046f90d506f13ffc6cf0167dd017addd81243a912b9b92d1b7c9325d6e10725c1d9b54a7207000dee181db37fcb2fd64b40ae5f52902f1c61d2be436d2927f8f18b7002fc0cfc12ade7cb41f466ed22118b50a231e0a7f784dd9da1da5d28400a11e5d43de1bee0fc30f75297c82d200c255cadb7ded16863507e5cc80b935e314580ba46a78a3ab16c410061713ddd46c65189d1ae0d35939621fa46838dcb24f840d677453d9f84fd7fbaeb8c72940a7d75a7452f88a251f867c2d8a4368ec5f23ff29246f368b878be083b3c664e61a0720bb718268ee180680f7f526b20b3085d0ae946470d6b3ce2952004b0594f5a0e1d73b010cce42dfadc1340c8dd91f3a3ca159f5bf2775c299fb1ef1ebeedf06e56094a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8cb52c028c3ca612f24cc5ed06025093944b6d034f14cd5dd732cc11784f048e109504787f519d4fadeac5498329f46fecf8fe179eaa904107a8099e56ebc1b86a5ccf88e35a1d5ff5c25f17fec2dedd81c0d897c20ad761294a3d6fcda3eff902bf42acad7e9e0656f3a44721ae73d7c35073f128f81e6174d5d7c1989377b4c9f9569aa5fb2af01323f49fdccd2ef343ceb32b22d7fa3d2dd2d8a6f09a4d2727946ae277977d2dfd0570d83a09defc6b31c201410bf1ff76675e4a88a82e7b18f91fcafadd0e7cd43976044b8d5637d74eacd2eee5fce016fb9990e5117512dd2d2d1edd188226b29c841a9fe0619b3f2da354ac7323d7c6063935a14c5be187aa0b254929ac999c621ade8db2d6b415a6fa01ce26fc8d3d6e8e23785664184cd4c01808e903666802fc41aeb61e82cf9c6ab910b734eedec1946285ba319afcaa42b5a8ed53197bb873219dc64bb74ccb35e28d636843fbd5d9ef317dc86c2a490ab8608294103d023a79c9170f5cb48133e490ebc863d373a6f1977393c614fb4c005bed631b563319c7fe4ddd5d867ef00ca9e7e7749ccdc6a82194425ec6e6e2cdd08ed6b3f34e65c89f9c611c2c75e11f85c35efc6dd0fcc2881ae128d839e3351cf2eb59d41dc5a3f341d4424c16c097af6ee10773c73f8f96b15e1783d325fa3a37836b0bce353b7836d7f6c9260d8da7cdbf504cd15cfb8099b9bb9153d1abf1d8242109a78b887b5c179eabca11cfe6e75f32877912211d78db5d07801514da8f01f01237c57d51c98f82ca510040360cca08237129ce94bab9e327fd5caebaa7bbe23a86a7e636dfb85dfde666a8022ccb4c613b75ef7a8b9ec882c524dd80e29aadadb328e293e2becbe3e08d091cc663cf444934b16383aa4a5e4875fb6b140b63725584cf6d3c45d1c1a96557f5288aa4a127281b3717aa9ddd1becf73bd48e0b5226a9f15d8cdb7f68d2beb687c8271b927232430654072b0f97c6d2e1d641d6bc9521d06155254052697eb2ac9bc7701df0c73617537eb40fa2266cecdd752e5eadfbfe55318034f11aeb2df8e9f913689af8deaa9bd7dd6253a4511a15983159378724e69c45f6e7f8c5aa05e5ec416019c6b867f87b4c622c7098732466466152ce44423de5fe0ca6115ce850b056e00577aa51d395f42c4cb2baad8c2eb8dbb8ee363a9daa956684d81e9dff4a0488e2b47450134b6e3c22a357ba3f568c2a18b445175d3941a16110fe442a54adee04bec6c9fec7532b57ff24002981b035fc1ba623a73d5e643613409b1bd08c74577229862f5362bc4392d8fbe2728b0bf40fd1aad0d3cf04e7bb3377c73c3b9062bfbdbfd1bea748f76ac3a58e902e22867754a66519730ea501b82cb9870e7d47a6add37ded4df0d4f3cd460fbe0641107c8cfb3deb4ab9da37c0123721a8a70e5e388a2aaec7901ea2ce901507404cfcda0cf14921aaee07d608d9edf93bc709bd0ae7e10382350995c7b1cc47a81913ee4aab8ede278cfe2b3b1cee25e235ec4d3b8f99b622f685b6a01a61c0b6df9d8621fea5781d536f7f346d818d994a724e755b9a4d75aae66925bb7df53405a2e0f1c442ab78afd50c70799e7436ccd869bfba46c9a35382d617f32854d527cdf2fdc68be800dd059524758c51e583b5fc31648a0041ede084a65f5e47f2247c4b622d0e53acd0e2f6d38cc889a1e60f25d14cbaac01ba4b2086d85da64922534f8ab496ba4d8b522e3755dafedf42941dca113da64e8485a2020c24d6ba42b1bf26e42bb334f7c665a1e28151350f2a5bf7a3187432ecdaa9c490b38ea47f04d78d5aada43fee2c0f8a4f10f00f4ec5c709eb242c09f0a9d304150640892fbd999882626a3b0bde2945e8e992a337c8968551fed5e0c4b4ed544216c65b4fef021ed8c5143c94977b7e4f324b6e0c3919953de253e35f3db45f89d73ee88b411c843e744c6c8c4afe9c1e01a986336d907ebfc31791639e5d31edc8c2aa99cd297fa618b0c6e13a8f5cd810aad49be534bac92663a764bb39f0ac735cf0da478441bd7a13b001693f2fe78102f482c550175152a231292064971faf13cbcde725a369e2dc7cf79bc6f49f9112810094a63171d099e653986535abd3a6c49dbfab2f92e56a5e51e0e61e29b9ed045545f6d2a42e33ddfed3f356c4bcc54571d8f2a4cef0f18b63c948d07b03159a5783c790bdf0938ee40238acb799edcc76b6b260b7485e049918b555101e5bccc7db79afdf02f97eecdcaefa3c10cf16fe275f90d16e146196bce2632958977e877063835e534e2e7f5a72c26d630192c4457798c733b9a5b8836493b4a11674751f84c73b23718de568c612e30dc8b96fb098ba647a7ed6f93c04c94490f24bc9e4b9907d87f49d7a4b1c187091401c39ccc5b87b9815bbf1dbff0cb79dd947b87d811514a69c7b032e17f4ea7d6ad16a95a1b2c8663dd85df0e8cfa390f881c58db26b6f350079852487e8499cc93e70cab5ccc27ed8874bb63d74ca9e0966c429ecd591367e17d56e4dcbf3d49d17d0f7afa0cb61b7ffa1b1e1a0aaa03a00515d43cde3e2e7cdf59d0859eed7a8e3bf1d9fb1e2c13bf9a7de69a8f09b9db087681413b2446cfb9ebbadb85b1c5d42a71de27967618858b4d4683173ba631780ff4edccfa74ad2a24999e3c057a437a0aba3f8ff9d463e9fd2433d1dd6ab0e9a22dc05209620915fd560474242e301e6fac393a35bce1f805f694c84808eb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2e595fed250dcc5e154f15233773003ce2c5298d568000f7b815a46a7adfcd32b7f2548b516c9b054122b0504548e646348a4d652475f3a80e6544c3a291fc2c7d1fb62795100acbc09a555ff2195da6a4a0e0c36e0eea41620c1370fa735cb7f5aba2b16102af258646721e1fc59311e44833ec54705cde22d3b00af5562b3606016ed43153acc13129b16f97935b2cb2c9d55af853149e7c8b49df886d5e797239db603de7b8ec51793207b3aed6fd2697b18c0621b4892e81c8b2f0f8d8a5593232d78f0f48738c74eb0cafd8435265bfde2881497d0f323ff188dc63326f2c2373b0fc6556e44b19a6c453e6155401c63fcdda4969e8b096f2b46c9dfdbe5726677692f089f8352a686f1858a1dafa49c65635e77041e5662716f59e75d598765e24b41d38d991ba9f1b0f03b6f24c60ed2cd9523fc45d8bc77665a4a5d52fda2956265436d80dd10e9b084b9cdc620257dfe3f0ad98085223fdfb800b57879dd78087e7cc770d2a57c84110c67569eb7ec2190b3709fbe4c30c7421fac970c1cedcdb0e5c4edf88915d6adb3ba2b8bede1283fc916ddc122f7a7c7e5b5aea2d1eccbe42a5f41221067e87e8680612da4f37d139f74dc21b58792800f2a71c5d899872fd2b902de6519ef9e2a8163bddc4a0ab226860a84a276fd2ec140b7411e39fc08a0049138078abd0fe46d3320a49f33cc015ce09e558ef2ccc7f078b68fab82f9d5ad35e61e68206a4c165e4be1e1747b428deaef783fba961abd368204119e691f1bc680b4c223089f9a8fd03f75db52ae10bfcb0755224ed309042a708628b4b5668ee6392a4468a5624d745d90dd848e819b61df1037bd2f0a137b28b8185c307936a71c3bdf6c0d63e23703ae41c9d50105391b418496d77d58b181e37526fc0b6a2cac34e56c801e473beab5af107dd56faeb09e0440b690bb33abb32ce15c8a67a4e5b6f60a58a670d33efdf8451b10f5829d4542796212d7393710a8f1a33b47279aa0b065b47923d58c8593dd29119c96f19309f4c2e80560cec803cfbef70cf58db025c00d0c6f673cf26094031a75642d235e60119b68034d73f5c4edcf8e13bab685fd6cf2923c27d6ae2298639dfdf293452661c2e57bfc797e9285b96db49bf05b2d3c37b4e9a32afd03676dcbc910f1896cb744b47d556032438583ef251abaf3f6ea867f23e8b1e36fe8ee625dd71fbf3d65593af84879f80b5032b1790e59c6e0fc587f5839f30a769019c5b914e9aa24d958fa3218cad5b71d6590b2d82cd273f91951316aaa381cb871cd3028a7499d5bfbfe29b09988fdbf95f000f60e8250a90c19ffa5099e81ccc0dc73e503f39477607a2da78a6a5c8cfe16aae1b02b254c73163a8e4ad28917c8bd0709bb6d79e05b3344241662c1def1203ec08a1645b904f9d04e0e50bff49c7e37841cd4128507e5ed99a06e5c5c6fe4d578c22dc34112ecb47547aa5c42524a1f3c0bb342456d57cc50e3cbf2fe222e528a426d553758b0286bf9c986760b263d78dc5afef91ce4e372f95c60fb35ebe203c2d636fb26538ccafffb44a848541866193c92580192c119e01e0db53df6c6cf12fa17ed04155e85289c50747bfeb9ff8b954b50b7e02ebe3689f939d07a38c3bb6ef32e3d61e3c8dae92c44390bffb58498cd4716ed7f104616b6c23f926db27b76f6442349965ac2421d72aaf5fd66c52537696bff64c585fb6f1d05e3fbaea3cbc9d86013f9f3e04bf104ff5bb338c81e4f50ccd15646a365d7f3beec7f7afb09041f4a87c99647871746d7cf377bd1e4bf0029b69ca4cadb9d51a86636480a58cffb70623bdf0350432e2f33b58ecae0b266aa44be2a903ae3336564831140d8ee3fd49f158fdd1f646c609f9fee9887e90d69c6089092ed171be14afbce5d69c6abee2b8b957d241ab9679ddf063f93f11fc9c57d39090157564b5765162b03eb14ac82cfbad385c82f21bc93f80569ffe5e89dd9521acefcc0dfdbeeef6881486f180a55de06da2321e1ecd32541b58894c66ef11533b5bf4bcd087e5c9cdf6551f79703b2dcca5154dee76c078ab61cd3623dd5b566d3ce70f91066851b31f97724b198926439dfd744f66adac2cc49c157a454d04cac4d13cfbd38a11711f2e605e9afc120030644189ecae0ec22828c5f214d26dfe0499608d3accd54afaecb5aca26b1e97b1edd7f625f187a4f1ce59fa15af595294957e70a5746fcab79c7a6b6e16d2a7aee5d048090ecda107cc38adfdf4537580bb5eecb71170dfc55bd05bbbb0e147f774415b71bc8abf64291ce1abd8f4d1e3df880b18d8956452fd7d9312f1f00a89129d376230aaff88f060b23a0d0240918de6f381bca9c9ba5a366ec1b0278d6373330bac4538122618c0f2d7bef3f828639da8152993ebeb9c4c88a1502955181fa5f60dfdcedbf919af4837f004edc1c16d9b40ba3bb9b5194a9c2b99ce4c84c689a828e71e31b9e1a5cfcaa5dc028ab65ec9acda1547ca1984797d9c206cc11039aee5fab7672a0cfc487dea8cc7e3bb493d79d9e4f6ff49dd0cc11952656d4b2633aec1ddeed8d45e3d932028163a551e21d366ceb6779608045b423a7ff68ab1add1dc6db9869cb7caa3f858c7cff9345e5ea412ba1965bc31a71e91e72b336d39d138ea3b2c9f3d6a245d51ba39413ecb50ba534c00fab2f92f27d44321a54a231360d19da88b603acfadf9a21324cce81f4b5a2b7493b51e81e27285e70a796c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd9601d42e2c4e3c6e7cd8579f7d77424bcc6ca3a73e5d6e2ca5fcfbd589bb779a4ff961fe9f8b05e89f353ee31ca555710b82305234d44867ada034441311fb56fb3f122a57f35983e026b92360ac584d335cb735f5802bb53afe467d2ce103cf962dd9fb5ba223c4bae73519668229fb221c31a4525cf2221fa080d2cacae7096d2590c4e5f2be5c3eb0ba18331f76ab0024f0f4271db69a256468c91aa402c68f1970879a689fb038c4e74a35455a7b7f1029a245f79f5baf5094a8b9508ff3190393b4939581b3e53974131bf1e8c07fdb5c505011a313e741185a9cc9148ee118b83baa6dff7e120cf15efc70d18616c3e05b228b32685d050cf579b67d39b2512280d979c568a3b9e8890f965a7bc347d4f471f6886f7847c4013e8f6b05395a4d8be229362fe5e7f53d83771c78c824ea595cb826b982c297e0cd55b25688ba6f063bd93320b09793bc98b773d42ebd69384afb2185b68c358074f6f53dbb4c94e29460a3a41328b8b857da35fc7619f8bd9ba6543b240a4ea7b7638de36766cab611b907a2fb969d803e834b9428452218ec7b4ac88872d780f8307044560659f0feb585a80c693c179bf3efbc3f5b503d444dca40afca8f7a54c8f5c087918f36a3fb569f666a3dc9a4c553be51b0c56b8975d825825423d0dc0fd3f415557a76bffb3e8a9df7c550b196b14f5bf184d0eb06fad3ea0ad1b17e11505b840c1edbc0b4b241e3233e40425793161ed78de852accc55b7b5def8baf3f7d8ebb2378efb52b3aaa5799ebc6d4108560398a3629cb05332a230b0760214387873042ff4f5113f9a2076ec2f6f9f4727628b87ce860400c7e5cd09957493516ed1ed1a2db218930fc56797f2dbe636f553dbe0f0f4ee5dc378e058dc7c4c8207f01fbd9cbcc848524e5ceb8d94fa214b9a901cc390909c648a8922332866ae45d5b49a66597270ad3038860cd60c82736247cb0416222fe4abf4fdc78be07e4fd7f1c85e2d8a160ba99d86d1ee5f5a263d7e148dc3b8ff373325af56cfb34131c29480c5b5120a87d014e9e262a2288d35e69b6b463454eb3433f498eeb658759fddab4af096168ba4670a8870ad813045c53c830c8e4acb6e5c2ca6f5b9b1fa2dc641d1fad669a0fd4a5675d221dfa45586fea98d99552490d02d71c023dce5d4165a87924c63433e1f52f6b205a71d014db735babfa0ac486d87351df06ac878106883bb63a0dd905813c2dae1bd08969d435cb6392d0130ef70695354d9ac1323a80ad347f0382261220d87e54cdb925c07bc5582eccb84c28ce90e0007d32d290cfd6c7256d218f7d2920d9fefa31b110910665e995caf1fc93168234ac3594dbbca5dffbc781e0b8a2c14475a05fe155c7508f21a8cfbe3ae7e71e062c9ac420ce91edecc08819d5ce535f2061de24fb8d56dba9bbddd6fa92f27bc596fcd4a15c11d41e62922b1d950c4d9c1c9137896e846145bd3902014107da453955253271533f8e7993db64d473db5eb532ef8f900a22475c58771c248e340eac1c9ad4fb91073b8ac2f2bf86e6f410a3aa2a5431f26f306dc969e79327006827195b8c559d53c697d2891202517793432953c63ff3544b9ba33492038d695b4960e5814566d5f7affa4f453da846ebcc62b117388ad00f99b94bc9ec0e76f452a4b0654564c1c58f9fa6f4568d1a4d00dc22ef7ab40aca9bad1552510a19708bf208ae77a9766d27d7ed00d800b9220acea6687791f533b814a07b3cbe8e2ca280583686966094ece94ecf5db682ec38ea780ebe47c54bb5279b86023696380c962929d9c45ecb37e65176bbaefe9f96346c6033eb46f0521a30eb876fb81b1d66b9f536762b8b6253ffb9b0ec06b6873bc4f791c131cb28a401c00f2742c3cd897d797d72095cd60d0ea8669f8f06b59f838a056ade945fae403d9d320fe608dafeac843c40d624ff49ec87b7b8158d62460f818b1c13d710c4837bb07367e2b8d2a4167b8a59f2a4d4612674331b37f49132ffbc12d993cbee2a254b1940bd65768a0e67ab010abe701719dab1793f5437d1f4c166c3b5862b2d2c9e46944f1e2919c0539b8459059f97c00d9e1edf8b86cf781a0e38daedb98b2d1c3f0889f299150493661f78f14da77edca758a57bbdb1ef7c1af0cfb446f8d5da19f0962924b796aa1901bac9ead646874bcd0c0030e26b168da02b97c6c40092b3263deb1e98ae9fb0d3f6fe42d52dd4542803f532501bd68d5a2381d293515a0ba78a3c71f4ab6808725ee9f0c54f6e11a36086c1227e3c46d2f505c937351153c08fcd81db4dddde342655520b8a09a6a6897a487b1e179c050770e9d16445c684fd97af6182934c8f3f5cf35c771ac2cb4644eea1fca0d900061be50c103036aa988cf20727cd503f551ab27bb0739999ca2b3fbe9a0b24ef07451efe40b923910a4267917dcb53dc0bf6beaacdf69e01a441be00e6e1da37338a699991a61fc13bf6911a50d03af559faff4d5f736ba0966a8ee18d580b746f6a757836bcb1715efc11758c39cd6e949afd2703085a742c656ae40bcdebf8c9a56de3ffcb5fe1cd1da2a267ec686b8a7400ba6df3b37cca0e04bb09a5bb5c70bd6cdf898ffa521a9318fc1b00ee5517ca46f1ba4f89defeafd42e6214c1cbe3e76e0aa0206588f0040ca3098b49696e1d0c2354bed0f867bed91f186869dc6ee0c9f986d68843e0f7363d46bbafc5294eb34d69a78d35d6e399fa1b6d73d181;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hde7e2c2683eacc168db57c00e9259d67ab6fa06c39ad83671a471aabff32d9965e2afb0e703c9ea93ebaee81a502d390ddb0bc77ca0dc9b44cabce58359eab50ded09d86d50cba0ba17a2e8593513c7a754343959ecd3278000e07f4d797de780b2f424681924a263d860dd0c20efbdd98902a9596649964c3e181ed7f4721099ab84c71e726f74f17b3ff0ba1dd7119acfb7bfe31e969b9f4f8d13b907c9649e0c399706e4ab8f7edd3984a585810aa565cdec8285ee41de2b4db05566acc516f3d9845e984d01ee464c0c1a8497d67cfc25389e71328ec0fe8f7ed2b737422eb5326ccb3a5de119ae267e713fa05913332b42591387997cd8340326c19b0df0adaf7e7382a5120a2386052e4e03df986c16b693a72819a382b5f536e1b4a495fbbc8157b3bca8064e0842af4f937b9dd366c132e4cd136a0126da4ecbe95ccc24b1e1a734f3feb7e027b5da9b5daf909f3b498bb591ae5da1779ac234d8ff726806429095e5656763e54dc20d9e3996c787b63469e6ff37cac4fa87e17b2e3c19b4c74e4ebccf1c080ba3986a41b20d9c5706d0f3908ed46eac5ba148f1451ac5ad0b7dee6d09e9925c4aede3cb9c75227d2e1d04bd217e21513c65f9a686d40419c9f673efc57b8b0d02fad326ab4b321f07da0d9c4952b8a23839c9a254b8d514cb3874fdfcce6a230a223c99d32bd7c85f3f9cbacfdcd1d46db5e5752b80418e84eb6bc066001c809612af584a16cce1217c276e29126c8b6b613819eaad040c8f040bb9e9f0d8d71ba242cf4f93a719125c2de58b51a291b67be19146d06117e7fe4cf8b9ed42b7885a4567dc380141675ead04771b11b8e48e9bad1aa8459a351d48c0074328d803c5a8d9397c7fe8d0458e099c69e7f621378becc968e4a7ca6923b4860a6fddfb8f79f5cd465978b931f951b0f68807c00c05e9bebb05f91ef9ffce2d45a27510639b586c57f157017d054701e3a907ba7583b6b13d198078b9486984648646339f2b95413bbe5b03094d4d55fefd22593a87a2b5b44c0248a44f17df4129f1e008bc3e1c23ffc2df48c17ea6622b7767cb50b1b732e2e383d547625a53ca020de5a14fe9e19bd738d0c717767ba089cbbca5cb1803d6dfe1549ca4c2977d3f24314cc0fe650e88cee2ee86b11e9d0fda3d09c6236b566d2693726c972ae47b350e5b2bc4d0ae57dd909fae5452a4cab8aa548f04c8c29dfea82b2350e7a0fdec5225b807cb9fad36e1929c4ef547dcf70866b7274bfc9d4b1df38733c25439a0eff4144cba95d5b10d0e43a228ddc0d88de57783eec4594b4beb7f29093c6fbe55f69734e048d2ad34ce6b4be5aeaacc5ee6e4ab2732adff794fede4a1c030055165b16dfca8a1e166b1ef2e0a58bd085c7683ff6d78b72ee6c95d42c446bd22f911467cdcf8eca53647b6d6677582d6bfd37cdaf06468ae75e1a139e8d12cab7532c3825143e6d7ee3a8345ddf95bbbdf772ec891da1527869692426ab5611ef3a884a8fceee7cfcb5cf65e89f46fca098285ccbe853c069b43614b02613fbd0e8e58af9a9be9367c91ec3b92a09ddbfb270cf5cfaf58e3ec97ade8c6f8beb421cffed82244b763fbed0b8fec97eced111f65572af84f2be0c082e60aea3851cf44913df3e674902ea8605b41f872af942dd9d797aa8c457710f351932e17190223f52089c86a2114c4f272a045d278c7fd4bbd9c21b2453ce38834ef022da0fa683cc9c41b3c46dce2224e26f8eefea4e26679a39d73f0b72097b095137e78b5eaa4e4545957ec32b8552a69902c806160b4b2f78d3de649230b76822768699bc9bf48043355868e09f581b87c1d11f65a519024530ef695b66d947b44765e57a8c9a2e1d85251e6f145486bd3d0af638924493c4ec0d3b1cd7bdbb6160f5af9176962d789e1322a72b8964c960c47bb69f43592990ccc8ffba29bcc9158cac9496e8ffe56d3ac64160e01dae03c54e9f1533381b55fa01b00e3e5ff8dc9df4828616754ffcd8ebb26258531dd018890541a121575d457861f2db6d7a81fa3ab598ed288d4da78e9c1a5ec26811b6f959056f2c0f8105503d127d448be0702027d94685a021efcd1fc02466c09f37b720c035fc8fb4e146f7d2f31d5edfb1f34b0c013ae890fcfe4ed69e34caac577801995e571d042220391fd594f3cb1125061840c6b204a3f04ffbc1e69856b4cc6eef2cbd280421673c8a45c122ccee409156cd971d0c681c4e89a67cf1e82cc0b5a91ad7491059a49340be909e73ee0853800845570c78572aad95c570e3a5006a4e4303b92d6203c18c90f60b915135428a97f1ec6c22c339630fe10204b1e788d07eaba96686bb53cd7c675cb33da4157ce4a54a6c041edc3b6ad69cc4e869e065694b67451c51546b3264a5cd3f635f8103bf28dbe14719e7d51cbac6e14fd23df6a02c8ac1b42de1e6e93cd679e83378477ace31d6adffce3bd87934bf9d74d5f894e370836f24d96e437f01cbe847a2a0994fe361d2d4b420ebe301cabe834bdba68ffd9fd140e226f1c03423577486db0bb757dd577558930a4bf05fa78bdaad8dc0d63ed8db3ab7e271a97fae5584f02806b7190f42c00d3728180c4e504fd8268677ad76d6d1b263128293cab71c12abf5ef939e6d016d8a91a3e1e767e17785cd16298f4429f30fbe58c6b20cc19a5ae901f89e55bc7c0d38e15b16e3605cd2abb23919b3b8e5a2a6ca5e58c9e6053248be68ba2eac9a46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd52f880ecd595a02838bb8c00381bf2dc08234ac33be26baab97fe32617f7a4641bb488c0b8212218555b646517fc4d7e3f65a1994b844e3c62c8f7e56bd6341fd2c192414f1fc9e0e5ea07e7a3da9521e9d3137f0ed2d6cbbe806dc60880dd22b2ee6cca0a66f38dc1ace9e6c9432ddd9b5eb7f3435d4fac327d53f81d029867e964c545c3dbb665becf589e04d9eeb9f6eb54482e7668ee57e7a74196fb28641380059a86793d6e03b1b2a603b51efd47e1aa87743f29a5cd641d9918b561bb2facfa195177b881f8250bccbc112312f36f6e2874447402e3abc54d349892012db99a10ea5438a7692c1c8c033a6dbb850122521ad22666c91314bd206ef0587a62a22a7263abca99862a1f02f5d0836976a7d9e5927c459f4cf48014ff354b1f3bb8f976ed12654e4f0b246daf6db8bfa3ee707495f896f20fb4ef54a8436d84af6c003e4b5e869f9f4be3027564e677c20093c5f46b9f822b3ede1149fcefb9ac1bbf7c22465b24c3b66a07889d056466e063a06fc79595bbe2a12e69594365f97db37679349a53abdb12784c5bc29248e6d4b347860462d4a83aab6ed66220a9c6dc5656fcea1c4505c8a07d17603ab208b86b8c735a949ec98e2e537f68b623227e3a47debc861e482e8a6177480f84158d7af4fc1e3871f3915603808275753a98c38ae1605cc043f737eb59be9745fb5257d60b5cb99668249471ae01aec183b722c2881465c95f5a68f97404f171e0ff3fd21cbd3ab3e565a7e4dbbd6dfc63f34cd7129e4e24e7fd7d967bb34751fac9dda8189c104cb5acfca99dcd0468b27777803fe01ec1680808388c5d7fc304a0cb12a5af08d1144f437010fa55342e223b654af44eb03c2d58681a18688b41737fb0ea1f9fb46ff09ae46db07d826c70218e9cb671928b0071325042f7fc10ffa5e3ae6949b15d7db4c0ac98018ee4edf124da67fa0228b9c7b416cba8a8dab4375420f932518332f0651240ae8e007b0b331ea84c751ac0fde25748015719023a7118235e2db3ae15208afe34ffff04efadb68a248a856abf0fbe0ff666fa745cebcfe0b6d2e6434732ad2ab5c83bf36eec346d21e50da63b358a32fdab69061cccf41a51aa0abca03ad63944b8ee3ee1e530de96f6ebc51c60534e63aaeee1794846082a249f2cb9e69d453d06e4c6177b5a04132eb31998104833b802904f363d1ca4d3639e7d4f42c81321e045f9fa933770bc3b0af2d0d38718888f02adba197ff892f03acf5e72ad5cbd54422d3732c073f6d1d436f9defef9a5e63be095c54f49d2446a01b3554e777113854c977e0ae3b8e76f3f3bceaf9d4f0b03ef9899b2b2ebe3fd2034290dddaa2a6821a5188a6fd2d4f44201a56c5ebc450aeb02110d64a5632c6887cab7f304ceeaea0612925c966c470f8c8dc751d86fc7cd0d5c6ae48087c8c6607d43ea9bb95c54c3891187b311af841590d4129d701adaea29b41619472781a8c54b233067acdbf07fccff57bf9fd20e565a061f5f4669b4e018b4fe15ee66a8c3cbf4167aab460a22ae401a32dd19abef7bfe3bb34b697241b35f8749c24b38adf0decd98255a178f513d3beab7fc6837871fb05a906c39c0e444b9851165bd3c2525d7ccd0e268db70f8d3cc1cafe8932130b9fe4c560db7162128f4f6c7ad558deca0c63d1c27e09411e18c64ab4eb0d89871f3798c2abeb140ae68b4cdbf0c263965e6dc1fa7f2b733db5975af509c90cf8eec14a500e74c09bd17db3d28ed32b3f8456185dc7066e1ca7283b99a4a9076152b461d789029ed8e0dda3d4d9459a4f1ac3e0b9b2f10ae6c8f328694cc687571a0673c246a37afa7a61ebd3a45307df3b7b5363d43be5f2e3106beb09934dcb0b0cc29841e4808630d7bc98b47f4e7709b22619b262d5edd07b87c868f97e7160146d0b7165f1eed741cf06c3ca6da62f76951f6558a8d3bed7b76989d7ffd0b8986809be6fe57c5ce7b34df537958a7baa5212055b3909e8f6c23a74aa4e85a71d77ec25d304d46fc6658f33f0ba556d3bfc6646f1ff1181b82db93361921983787d47f858932d124810adbc5f5a0df1f2f1145ce37de9b730d4c7c36cb03779f7f0fd889fe0f0a4ea84204360216835e8b7c1eb239bd5b85e5b7d317b125a09852b3159bf97e72c5d480efd572422d2c90c129aa538d30985ed1fd9158c9fa89d9cf2d6ff79df674a868c9a55e6eea65eaf23fcdafce39e5d55334a1c1d9246423adffdb5441723f5c3a189fcdcfbb876edbdd05d4b16093cc00125c0a3313059c65a867b777ecc588ccf30dd35a71496021173ee772f891bbbd989a8a71cb1c011407af9408e560925a7c2fb77e7c9b777bf54d165f4d991bfb6335eb8a49516c0e703b22b63dd7181a3980019a1051658cbd24255466970cac745d95177365dd00d9f7b23f8c4249aa60b3fa3c68d9553b064c21361514c283fe6a515e244f0642749e9e8b1587be6c3910a7f87b7a38db427b252a9ea81412262f5bdd4335fdfeca39e221ff76395920ecb23388beef66d2fe73234e2124e2c3a34cfa5251ec0345205a5f77af254d14f027b31d8ba6fe5e1bd8743da3f4f21cda0571b4fd7194c38eb021a7308c184aca91b78d50ef827c57e9411c514b802c755281d0d3da8cb577ff40efffe24f31c1d5d23609dcb3c01ac0362210ed532eee8b69cc2347087d4c88392bede52cbde13bdc76ad764bf3b6310d5de0a9d0cb1371818bf7cc7959a00ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h54316f230448d32f9655cc0d5619c7ad110ecd9d2a67dd874bd4a3afedae4f6c55f1a6c6aff48ca5d2da11a9a6fbe7395036f3432f220316291f5da53b0078a402022688c7fc0f03c999f950b502c53721dab42c9a8a8c1300b47d7e9b1ef21245e4528d8d10f06361f33fc45e798f1a4315c52d3a6a1099aea8dff8092d06041648de35d3956c0e96b0166b5ef04401d46160b2f7befd232e5be362b4f06e404ed10140df69e61dec35a227fb2ac9efd19ff97363f7cf630f88e4195e03d8c1529f0c1c04c072e290d0c26ffae1e0bc9a4da91e6e51b525c48141e303a68cd14b8559e1f1a69f08cf8edeac6b52fbf6272ffed1089760744d12e73405d6e2986d4a1663663e284ffe539ec5436cdab929d7fd6dbbe1765d64b9fca1c92db7394faabbe2625f7dd5763bffdb25013322573df142cc1557fdca7ddd6b9a5bab3847c4794248bc946b173d1f3a43fe8abfee095fb211c2672b14ffed41c1d565ac0a33e1e0de6c7f86f3a718577656907ad61afed9603cc3f69a6acc364fc69e65aac1811474d93a9367de5621b871449c29adc0f5b8a571376ffb20fd0094204d8f7e135b9d15851aeef2a807cb5403538faac7285c5b432a1e403ce8d430f2ecfcf0e67befc3b2905fc2580dd19a301658914b6e3a772731aad8d9f6d3b8f35c3bb66ad092b1510cc0722554eef1003e5901b1dacc585bdd74c84ffb5207dd6c7d342dac5d4f1398eafb65848305b952b73f4ff32c3d630a67a074cd19317d2aa7dcdeafdb40f3dd3f66a6f31669d0c32a265c31dcec2b0a5ff092844d93ae2417314b69c3b64f3ea5c55d098eb8edb182b7d1fe66bc0b4b944813e18d21a8c3692b2f9ec907a8439be50619a29689c713d1418b00186b935bc2d82a2c65df4b5ad0e509b8539d4926876ee6fd438703ead8baeb2ee334e67e55fb6393cf375265157dabc7b2a58b5c9568fd42e3f18503d356dc08c28b44cbb64646fa0297eadf0a6a6a2f9a8f8c6d7edd240f858969e31ce78f270b24356de0c1d7c631e159d3d3ed9ec30a8f53e03032beb5507456be2d6b3c611a16073c754423ffb8587389b40bc13babee7309fe0909ebe8450aab915e4424066404530ce23f7982e592cc34cb9f4f8672a181a976c61cb56cda3c3077ac69013a42fc3e6c0be53cd7e8ceb18bcc95d09ac814f120f4e2bf464681133c3278fca5257e31fa24d578ecccbb088796bc5f99e1b12126e497ab3eb646b8d9afd7d331a3c5cf4f342abb2224b80954fc86cc38ebe3171bd7cc76ac73c53a4a38b17e5d534c901b7401f9ec4eca69b84a893b6ebd8636caae5ea7423ed521afaf08e8b0a239532d2d4b671612b5b6400160b1ccc641b868b252475ac98d1f7bddc6f976472d2bc9210b9ed5fdfe207fd7180bc98f4bc391e688a028c374ac92072689f4258006c5c895e2a06a65bad57d5a4f38b7eb6e96659684610454979015e91e48986883c9279ec9db7ebe0b192905819562ebfb2135961b4ca9af8af021cfdb3ea541f99ebc6e1211da3fa3eb741b460ec9932022dca12ada833d365a0d91f5e7a0543a60abdb2a5c638633200db266a820b2d767df71bc7bca79a48e1d45afa239268a7a903dd83b355398a6dc9a7304b3ad8a6f68b9bfdde3de574bdbc40706c676113c97c8d79862a8caf5e819144bb05fdee13b6da9226c8b7cb2fab7b6bf2537e831848124a4ebccde4a32841808caac1c07bed21432cd7da3f064ef7aa5f9d1392b2d2d633216e7c6a50bc1b41d31ed3a981a94b98d39ab04c5e2d07536e4cf68a4779809ca376963da19940f18a53ff01701db3e613fd1c7c7353830de01f637462847051e8592ff386aed77136295f37b0a28d0f4c7a841f8334e92d8fe735e07ce2bc9602d8cd014f31941d1b308120eed88a6c12a3ec250eda740d4cbaa7664e9ad09d48b4e8e5ed0053a75aa76d0143001e858eb242615238de2c99183f91c59eb39e4a885cb47cfa8519c5aa1db0e9e1af711839d4b4c3ac3870b986f2a5ba528b52babfc8beed131f00d31bf782abb81d9429d9bbc3922dcca651229db284b5873c14c6a024b8170eeea2f39451ccf610155b6f0cb3547a48801d4c7e022891c7e14e9471736998d4531dec6b539c99e411de89f2e0986c813fae5853c27a362a5f5aa8f4f2292b710e9fc57e1235c2d330cdcc6ae697d0e38be55ccf0ae7035bbd874a8eaa33248ffe48e76c9d04d285fe22358da5b1af0c776a2814e7542c42cf8c21f4f42860fc9df2a4d83b1b24b0726024ef95dddc7bb69efcfe68f322111fd52c22b2f3cf84d62213269b33ff2940814e96872be9ba842167e01de6512c43630d7fe0bddb38bc3fd4a198e05055c886c2a1720387160b3691180ddc68581edfd7a2a35279efaad949f70e6086abe63f594a8558b1879da87dd57f7107057f824c5aa27c2c3a3f725c967bcb56229f8f13d5b26b2a8c3c3d770064efbd1ecac433131fa5b5ac491c36993f75d74d293b92b9713f5a107ac8b6ed6284cbff418d368fd00394637bbe226be4032d00b5f23018a2d06472c65752d888db15be026b464204f41dda605e6bd44b5ec7241a68e3b870a08de86573dc3ef3191dc359746b5cd4e51aea428af8087cb17ce1200ae01b429b75d391b41e9320442a467997491bf54f77eca7c648a25571d46490b7a18e5399c6a4032f8d9b93809308c494b6f1cf64929a212a4909f9a2eb6c78074a9f4e29ecb4dd5a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he1a0740a7b3b847268bb550905eca6226bd418020750c3a802d5cf7fde92a88fb8a3238309f797c182c4eb70c5d3c8626e181c473ef2f81ed8ca90cde996ce178d0211147cdb165375598d6571aaa9fd05925b5e8786fa70b1599b98a5a92ba0e50be6bb3b253a47f7093bf1de27d092f23dc6eef29bfd4e446048aa50bd81654c8262785a4968ba97319e1964471e3c35d69ace2ca99473369aacfc45dc604cdccc482a58a71e84ab993cfd3571b17c941816626bb9637ffd06a6687f04efec4e8ca068188fca0265219622285dd646951ef5d69077034dc677002458ecd34a545c412ce097085160e0e492c811106d4a598b92cff800a07aaaf2ab8b073cb21098a64b6edc2d204628198fae16c72269a0ea5e90d6b218ab0157620b497d98203cd011d8133c280fad0786b0db84912c11d1c0f0fcadd52dd23714a87ff63d73c139992441e07ba8521b9627344f6fe1cf02a1f7bdb133bf52f40addb11ed528aff3a6506027baed8f1ae04b77dd9196bec16613b5da8110e69adfa3f3abf8684a23e22ad57954176513365eee764474bbcef6e3852512e1332cfefdcf8b2e673356dafa97a11c9f873dc3f5dda0ee229ff420e46c93994c7b22429325568b18a5ca74402bad4742ef1ec8833330663acfadab2aaa015711a225a0c2e88761da058ed824684439167ee6e3f47c80deedf9b245563a98689757ece0d7bacb2dd1bdcbd66385d44c102b8b6f513e3f07133939306a42ce84dcd06a06c9316b2cf5fbc0b5da9d86385e7bda3c58fed36c43a558976c01a6a5e00e19e43fbe918627b9f6b7091913ff9df674fbe086f8dc5e9db92f20423e00683388edf0ef3c9f0492ae3d80210c20e4582648bcb2c4709e53c7541c3c936d0488bc9d9f290ee3a5371d6a83626136274584c71df5dd370c90b4b3659db766e66e897a23c68d4855749a4613b5470a760bc9cdef2811ddd4c31a39716011d75b7c260e219eb94463d6d16dd2ea36158962188600d07ade35d0c4cc6a4d9508b34d37e27ba0034f9b2dcc5a4b00438856cef48439b29895db1d3d2f44e60943c59d824a392158104a09c50a36a74d33594f11b0306872168156176862b36b527d9f1496f547373f12d8aaa98786262491bcd0d7ef0025aa5e9d14b9909316cc45c3bb3c034e9b0db2c819a730cd722330ce1736bdbfa495f2998679cf6dd6e1c925f0a70ade8fc3c6d179178fe88c4fe036d19e48bb6009dcb4c471c6e7a0ff20cb5232b1fa7868bbaf819018c1426c753212e91ccb6e77bc7102c7ca75f35638bc4821b47ade5cf7fff92f5a2d5e9af397218656ff666d6dd39f0c218641c132e4bcba5c768b54431b315141a95b92d0f622bb62debaa47b9bf8fba736b64706411205c6d1e221306a0974a248f02fcc1025bad73b25315c2a21addd38e878365a146792a0852a9eb9146ddf97fdf96a8b8f32ca495d7ff6c4a8472a6889dd0b90bb5ef555c3e1f08ebf8d64cb97c292141095d14aefee001fa7f3c0c08c66469d452e62ff861212ce2787f61cd7ac15ae1e894fcbabe2fed410f3749912adc53cca284f73a39a0c54bbe737a3b200ab11fffc8001c502bb4d7cfcc734002cd9d5d4c77d2dee006f2cd5d786032061c149c7a4370ba857977da12ec2603c9b81a2a923cbdd08e2cbcc4d78ca6e7f87cb30b42f0733b3743fa6f56d702cbf6090c36ad6146f30f422a7182b6bda4138c7763753fb9f28b83a593593f2b82a2607402083a2867544f0758824f5dcf75b061b7b04585f576e250026ecb0bae46fa21a274b99a8af667fa51b8d1b1187e908dd6e5771189b5c13b907ce17cabdcfd3fe94d8a24e000cb7832506dd00b21294ccf1fa31d505ab8e2971141b62e5bc7fa2d07a4119314aad6decbc5189cef4e9954939b046602f08d904ab10e1f7923641ec4d4a93870942d3b8daedd0a6e3488cc4819cdfcc1bcd6daf3d3c1f07308e3241d1e0f10da7832944cebc3cc992ef72b4769ed7b21ad39a21fb8b927bf6b11e849b50206328ff906a93a1f35e54b1cfe75e7efdb3ff706191499e87c49e7083cbe57e540881a792d74cec79740defeb4650e6470b16b95369ea20cc365a118afa35862d4a85237928655f50414e08d455cad0ad44f162d60b7014d3b6205a79254a9e127f91e0192a9443ca152c47082f99b67d88da5bbbfce3f54dc55ccb4122ff609a7919c143b378c106ee2eaee80c12217c22f91c88798d66f1f1404e16b9387155d79f1e012c5a4dadf72969c623571be6f020f3e27f9f750eb8a1379510a5f21f86bd904e3a5ca762c7348bbcd65f1ab085f283222d27791a856e899b64b59f9ae19304b52fe3b021640a0f77a2cbf4bc874ed498a8f907574cbae6e61a7a4db90eb0df7af175170754d6d593a0c161cc087099c9e287249591e1c0041c2db03833292137e052bdf244cf892fcf33fd8e01710f7e9e7c0ac893e5b814cef66a168c0e9cb56746f209f96d0840c7aef398ff7c148f2aa11f03530624a3b0c3a9034a5e6f360b4a44d1df3a99e6b59295d85d6cc62db8ffd2b133eceefdb4b8200f22ea0a5b7fedded751173bd5f5aea06b527412df187113a10b2837df7ec79fc77f72f40b76a11843601ffe096e823a2f7444363dad479f4c62d58fd911c663fac77ef37d982f5f2c4d36bd8d57701ad9b1bea223a7cf8d6702ca99f393483167aae099a2cb6da44f8cf3abc6c1c7cf7375edfd426961bee4541d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h83d5ddb48417db92b66032f70012b8482cca187cb5e4be15088345b426ec7709bb41a6f909a9c78e7ddf466c4b3e390c4fc5ad4c92b16db764295a3e8f2471c95a1604ff0f407e1cff094892d641a0edf0a21193e67bbc456dcf2543b4f171af6a450703c541e630278b39a85fb3f7f7c681b9f189650b184dd947e447136dc307f055a51dcbcf6c4c37f538d190850472b9e2655e49df0690a208ec02553ca93789c419815feffbd3564f98623e71904da8d82b0d7b613297d7443465ff9324105b0d7bca613eb3e174f0fe60329be27a455fdc10034904eb820fcbb8855c52a3470b1b379af47f0384e4ee0c871730596beb336b63a09f8be8e1afd06300f0617cc3bc5ac1fa06d57a67d92bd0355f51024a4eb619ad34c7a2e6da879b35b004b7457897e8422268c9cef44c64220b93344dff87725be9f60cade1cb251f36a258fb23e6211168f208ead56db296ee3cabe68b1ddf493edd734d5b34f00485abb83a874278ac437e9dad6cf4e5aca1fb6e3f367c9a6344c53882d1bc8e340b75465d882547bb599c36dd18096b7f5fe5051c980e0b12136e9f18f8732c91dfe34c40a8f025bb18ad29bb03e59519823f7159684932b317a4108ecb79712269869661f03d8ea7e8d50eff15bb27e7336927909e1fdc0b0f3466082c8b3ab54a29c6fea3e67fa5c21ea3cfc9a92e60a4ee9f65adb70e749e983bd9156a847bffb07e1d374558127ce5b4b420f5a883636b99d9100beebeda2ee0db2697bc89d4cfc0d48a5fcbddb03cf89d0ba8e8959487768f7fa4c50568c2e0314459c591dfe077a5ad7aa9539b80e0eef3d600e72f28b2ee3e164c16bffab0180edb30114bc1d4a5a34b6d9ba7e0f899dedfdcb1e9121548f3b4b064d10765fce2fb84940a3f0102e3c6a7667e1596035ca194aa3420438590f7471ca79caa9115cf51efa66478e22ac28b3881dee30593992a621d22440e358ae04c8d35833aac6467cd496efe3ddc46f94d83cd5e6d377bb18342b60d5797daae789931406ace759561e86e240355223869e578257871ea05712bffb9e3205d620bf79bc88baeea6bcb6b5b75c65ae7500604314b5c395e9b2bfba91ca1a17a69e3102f7a90fe6831ab76ca628a88804376bab5f4fdc792bcf15aff6e783e2f11a87e9fc1096cc0d790376b81d9b6a40334ecc0e8aec9ee49aa900706ffcbe5a2f71580fafe670e6adab41ca3df61b3b8a64a4ed19da67827726fb76d6051c4c5e502bb768f7d5c70e4dabf1f19c46dbb864087afde1d5fdb4004da10970d3359115a6e5c556457cb7d04328bd7fb2b81a879cfe0c4f192169abbbe14536f78d094564d8346abbffe06ca84c53295a8e569b6a4ea2cacbe5268925cf2f6b138e34c5aa0135adf5b83d9a81c30da98e4325419e7dbb8ad0ce89ad5332dbd5b29569699cb6122484e6f82b9ecaaeb3413e9ec42a846d9d7ee38648958498cdd5136a00b8deb3b95d17c3a102ce64ebb05a3718d70ede60c43a1a4ff12d383ab465064d62120e243ee1909c249327dbe2ef9a7ca94385090c6508ca332bbbbd6cc2a76712585c6e4a3ea2b862e1e2d2ed911935e56e887201976fbc8afc9a35e717290159d6d71d563b800b392b6ee1b9acb843766eb066ab0587ce3d30e53a2e5cb7ea6911454dc260b626a82c958e52cb9a683d6466e938b8a13a82069cfa857c085f376efb64124747dcf558adecbb42555ad5ff38678e42ddfdf40ee15fd2b02138fab3c8e8df1ba6a15605028ca8b19e86a0b56d9709d65c221e5c7e045431e669444aadabb370701963babd795a28d10b9e54b5680461e15408e8d3f5c704c0650a7ce947a30589310c02373676f04b0de027cd4f68694d08aabd519bfdca0792af1fbfb74ede07ee679283222c3a1b10851e444f1a0c2e277332cc6fac3cbd6e382251ca5844e53d3452bc27fc62a7981ef1a25b7cee126958404625f2533f53436a4ad8250550037758826647d4aa9004494231a77e5391e50ebc56a5fb03a19cdd1afb5cce96e13009ca0f81357375c0940cd4d735265086ab3f331a755c218759d62055fdf3864a1dfec78f6ddc8bce452fea673f30735eef260f72af74ec677f5cdf46610c7efd64dca29e3c3cf2ecfa839061565eda7107ff652bdf4d067eecdc9de5933fa4098d7071d6eb5202f11af7618cf18ff61c3cd623e69added2f4267db9e64f8f43ec4f0a4008bd8197acd4fd5b0dec1957cccb66003e5388c9fa6ccf187c148212b9a37f355e487f0f124e7ba7e2b8e45bb2c7e187201c85bdbaa542f747b2e93a2904e9deb5f0902c0132d2bca42f5ba34e63dcadfc32010a52fbca6ce52cc8bd30d5230c36fceb037263708ef4f87414a51de52bba595415de9d1f64e9e26fdbf96a110015e9c9c3a70820d8198de98f45837bebd26cdbcf8e02040f2c824398b9724aff366d1c626d8e61213610486adbee37b757935398e71ac1b2bc5517249e0f140b705826777ddd0144c97132adc4ae15b3b2ca99e3841acc15d0c7f79f535c736720c363bdb70bc4671d31c01e27c7b06148d29a5c9a24016a41d8bfbdd43b5842c54231192dd61226616a70cb3657deb4cb700d23af5ce3344ae65748927b8cb0ac7931836a6553aee46abfee5cd360e7e94b4963b498eca584fcfe0bec6f9300beb3c7731923a38d2895358c4565c91b7b40d38b6e2ef94ba5cc95b637b161e62cc8d479b73608bfb92c66df3fdd44040ad42c5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3251bf93a040f5640e2de8a406a0d6acdf8b186a7b64857f8cfa8c694b766d06a779d2ddde712f9359e7b5663ef2d2377c66b5a9e021ba8854088aefd1a8d2d18c9fa27b66d7d6771cf9d4e277cdfe11aad96f6625ff62e1e8a2270e3f8fe099bc36fa4e9f6a5b670c51f2d41c2668fe834b58069d852ebb6f84cb0aab1ea61ca0157576a09b7ec521ff525d903fd176a4359f0433e80e11952dc245542a70156955dec9f48fffe1b6b10f760b6345e570f7e687225e194796cfeaf05bbef24cd7ed8f65a6be0faa657f001f5a72358c3ed71826ad7a8b16b72209af2fe4ae26caeeb03f5c734de0c942636225dd76582c607fcb7544643364312253a9a1f4bed978009513f4ea3f1b37d5dc42d2cacf12b734fe681003eb2a76d05a0b6b0d2a1e54df0441cbc53f1490aa62d1867c090473ff646f85d765fd451ba1b24b0349e054d008d4d7643e88424db4982e7ec16adcbda9d0d11a7632a4770c55a39a35906843a2d9aebeb7b65c3fa5c084eaab5721daba0ca73b75c0ea97c0a8fcd3e1e0671891e02cf3ee240d4dbf02d2900dd6e79489e138d8ba177e5fc475039b3deb081d4d5eb8d5babbd74214087446d9caa394462ba9b40d6d5a76a8235a4e39fb4c412a59ded463484415fb85a475c25610e47ad6c719eece130a8c3a1c0b595c468cbc3864e2425c2c20053cbe3533e344a17a8543b79af9b1b73cb7440787758130d25831d011fa61e371af50859532e06096f3efeb5aba38aeb66c896ec678239a1ea45ef994d9d8200182971fa062a33709d876cb0c2d5248ae2a1264059525fe64d533b6deafe2185dc932b509f192c5807ebd8370e6bd1b57844ade83d7292c1528e48141d5b9cd7512d8e995f583169bb98ee66edbb0cf079271617725116462a0ed3faffa22ec4e0f1039d3e66b3a1088688af6417fc6a7c3a3438dff605170d2639f380fe5824114fbbf8ae2ee71d9f3cadfaee53c3e3825174ca29bc56feef68752011d712089310d9ace55aecc9a160e7a6b7309ace3e42643a9f11ab7fdc0791c23a8e7409ebba598a4c55a8a2054fb2dfb56c3c5e9523d2c093b8ecce1bfaa4300c79d8f61708eb9d07dded31997e41e53701586eb1138fed90a90f264808006bbe3c15218e47330b55a3b43101821f8c291e57afeb2f5340be6e5a5d320b3fff0d466b1314025b062f23015709377bfef2c8742821181142756068319d54472127e34afc115de023996a188024ca5c6aa1440324ca6ddb40b3bc9bc9099301be97526988eaaf3bfc82ce9f7ffaa67f54a8151f0bf271dc9e9421bfd1cd689d8faa6f4d6b1b3d81aef3c59e9fa5cb71db2cdf652470caeae8986c9e4eb840ba499d814033ece765f501f841e1a0c1df945105761ea015be25b8b17f9d0c1fa6e64264220a86ce7dd6aacd1a0c222ac646d4967f16d90a8db67037af64115e135cd437510609c13f04ae2d47b86535bf97707bbba76f670ec157c536a0b914ebee14eb2ef0789f317d9811d218b0a01fc35e3a4b9eaf45d196f3ca6d66af1dfdd1de88fe058c3e53d64d9f12b2d99e500e8397ffba19f7a8468883a30e19749fa45cab353055aedcb418d79557faa38542ce08296b303a4627c2d109237f5daa65c69966b91bed4c1384b1963d032c7dbdd66b856d73df30282bcc53ba50dd1bd6b4f4ac519548e73522de872ef28be70f8dc7ae2019cc919d43c32cb6795a7820d5a52c8c61638c6fa895029ef1456a7aa5f4cbdefed8f1debcb9b47f9022fa338165c3b66ad7eb11b6a711f6433a3218583d17e1159e2246d40e7972d63518441de5e560505b559385d769262a5ec10c87f84a6659e6b8b3e68bac31a729125b3d63654c02f7d6b6b0b1800628dd71bd54747af3adb29965f78d3cd3166af476231191bba5e2573a47990a9e5dc70c79c2159992d0c49753f76599e6e150c18e970366c18982dc1c615ee1bc36c536601df22195f7e34387841190da43fb116de94bd93cb0ef9accf460dbf6f734ad715b6e2ebd83951561e494ad4360a21cb65294c39245dd3243479f490c9ce0423b75ec784b332a9b61aae5373687d9b580c0f797023193ecd8dec13f781c734214c7e7dc14dc846790367f5c6800ccdffa5ca598244784ec6ad25667989baac6d4c82b0d1345fa1aca3edfe0ff0a1338b94472d8e2d936b59cfcc695ab362df9653e8d2cb78bf2b40e6d84ba8241cbc0ca3fac38ebe0bd82666d957c890746e184662cf6efce101d475adbbfec089758062db483f972e043c7b3283619b8cb7acf6334487af95bc2fe34e69798aed6df6f0f612995428c354293efd7a37f8f259682e460e43ea9366233f28f1c3214fbb6bdb8e1f055bb77490075809a69f7b9933f9e1c2cf3f99abfcc13396479e67179c41ccdef56d688277374024a9dfd40b24028e0715a7f0bd438c79f64bb28a707c92da851d1a586776bd2e891f0d6d4e275521fd575834628afcb908f3656e7d16a3bb8597d0f1a91dacd5bfe4909f88989aaa3670af3c36dcd281573469ce14c87abf03643034002c82a6e0d378ede38d104857b96ba4cfb5c17be43d69cdd134a3ac9a94af015de787bb078c4e0eb3866085b80de4bad84d2658502319ee02984ac56e3e2afe884357dd089609026bef9f1e420d9949d5cae047835c1ec3802addb3275d5fa00b76b50190c7ee432cec4c72d5724359c4f75e9a126d95ff3341462b6d523df0422632f0ac98b5a56c1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5ae982219ac71f8ef82348036b827869d652ca3319ef3da6dba290346c8fc15174ef20d6dbd00e62ad08dfec8e833048b1198cb85a134dd16351ac434148ac9847869cc5ae4bd44b335f14d5af2bd3ed3a4845dd1cfd56698916521ca139f6c3e849f53c461b81e327cd665d3b6899eee711d0a6e672fb363f4fc0bbceae64cf38a7158f31d6c3c245b54e0bf28f2dd612afb4a9f8b088341b1db7664fc6ee741f9c39a81309c177f6882661d13d2bcc78e75d9a6f76fcad3a2f9c62ccb1bb803381c97744489cd81cb7262102ef20e056f1f52da67822ead52503d014f478363580885aa59d9cccf1916049ac1eed9d5e3a7379f28d00ba43ba49334963ea41d95e862f404b440d8627482e538d106ab837d25f8933bb4af112d34bef082b22e7a7eed8595ec9d46df52132fb345edfe0eb175680a46edd21d1c759aa13a8d513e87a1e260cb3c141c152a2357c7ef5d6b890c6504dbfd198370f8e3558ad638f44453a635733efec96765691147639422df2e915ced0faf8292b2393789954e9b48e5cf1784de97bf2ac8cbe30d98a830071c82f32a72c11a0987791bd432c73caf9604093ccbfd8868104354444bb8825a7ddc3f2b565fc212f871b2402d551a5cb9b7f1703e8a8642f7e903d1732a07004dcbf40f4c8a75372723ff92aaa9440cc48cd202fdcab9de1e24afcc31f47371c88357a35c3315398a5e18349b0f8eaf3cb8c88c38cb0d8be3c30de792b8ac4cf9408cdf534cc2143910208292b905b6783bb976c845b5c8f6ba5432c5c265b9ff1a6772d350b783e95840dfd592540271cfcb386d883ffe35cf37322aed6caf7544b648bea724f5346cba84cabac2ee66210d68beb3cb6589109bfa7d843c68261644f2e7faee2a2dca9d477019bffa88fa6be97bd372c7a6ebbd779a72e17c6bbaf621fd6026862203df4cb63fc6351ec114a30e69c278742804a896d3203dcbf7f0596868f75e6a51d46b85de16b3e7e329d61026b71099f1f5b353e914a992517bc7319ee732aa9aec8ed13a2449639428aa4be41a7c816942505e9515aad6a1469954e25822319c287ce5b542531ff769276f07784717a6e4114df8e0d4cd29d1639b6f63ba19dfbb19597f3e17140398397a3a5b1a999853b10ede5ee6c8c441b39ac994c826aafc746caf5e18ed640b1126d3f115614c94f87ceff26ef816b5e3708d1e24747b83bbc71c67a75ac8b05191986d30a3f9b29dfe1937908aa648e1a1b2898d1fad7283a97c3e193820203e8f09b57db2fbb455880e73cc607dae739a6f86bd419be42f1a8f8cc14727ab367a0afcfb47e6afa56abf564b0d8bce47cdaf27a5faf4ed6b37dfc10e031bcb0f1ed34366aebad12bd6daab4a54bfe42884d7f8b993ab10e9da982aab98c249894288cea13cec2c7efcbe90038c4085f12889915b6fa61369ec8eafaf9bb4c60463745440946d6a1c0388f427a70fb5a609661d82daa505f8f5418883c7d48d30b5ccdc530ee1340c7ee71192d2d2a70dcd7fddbb74abae42e394b9dfcdd1c2544f8cc4022f0e58992acbee6621727b5230f82495cec44eb37d3fbab5fa7283b05e5601b12d950bdb598e6af499828ac27e83430f4b1eab8c0463f8bfd4da8ca9f055bb9c4b65e42434dc2c6c15e911d5cc063d39d677f4a3ef7045caf9ba63659a34116e0e43794b99156b6a78b122b33b35155b4e8e8c812ac112354c9bcf212daae2be6c8b8dea25fbaa1d33513881f29575d80cb16e173d23374ecde2921ee615f1c0e1d43f12bd148b978eb28211ebe5fe636d3c9e59706d9dadd96ee42725a412f0c393517d4ce3cda0a5e1fba02789f2e22779cbe50c8c9844a413be4a914d57a758c67cff3878c2358c408df61e9a65ab5c56ba42e1e58ac2d231374068cbb8cecbd0f76e5947b38f0bed3bfc592db01bc7eb068e462a46ab0614b8d837400308590512c9c4b73e5cf949f400369fcce204dfe9b2078944ab90b95a5a435435027e21d8d93d9f642c78bf69d001a29d11516e7e544baf2298931e18988220a8353e6a6d0deb4205ed97c6c6ea5c14a67b3031f0a8d20dd2325b0a0ee0bea0fdfdb398dd3703b2d478289362e160b5be562ed79e6c6e2ad08eff41d647d61139eafd2c7fd92f33446abcaec7ee01a29385592028a0698de1ebe4eee2c5b3e1eafa0c8511c034f871cd257aefa08fba230e5a0f6fd1c5a1ee5a740eae244c8659fcea60b2973341a0316efc684eef53100f76b7b4ccbd35320c86f5fd813fc121deb67c7f5b8d19c2bca05c3a754efa4ee1fd44c5fa875333a18869d4e9d513865e8b8ce3256b5fbab86d245b0c16e87f19cba6b0621c06bbd3f9f3fe0d40bc3a3bd73664745c357a0e53ee4b0625e37f30fbdf5bb32e2cf4b776801c598d715bc788f5c8599fb62ba31807fce6db62857e9f5008ce4760f443f056aba4a3aa0c42cc7a5b10c9fbc37a3cf120af5f69360e6b4d1b81c5e73d448ddb775a59993e6b01ffece2b5b19b35fb9504bb8b4aeb40a57c3f4fae0c0e72db3bae6195d5393e6467ce269414f23a87352d3db81c1af1280c707be0923e6cb4c5ea5f567eec01b874b43b86d726a843912f2216aa2e7c586e1c4206b4be8ea57e849c760bc67924f6417c8b1095210ea4260e39ecfe19aa0d342f98a997c2f8db8ddb9dac551311737b967ce0987f78f32a19df77204548a0f64e5ff3fb4db7c647f1a3a9385c48f92ab6071b96b421ce695eed5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4a71436fc4283560f42cb42e7461c5a02bb4aba01f56e5db32210068e5dd979d693ab2bb83d92954a4c56c0c91c8210b700ba0360f83877c87f80f678839e8804009a198130880c78e77fa6d59917bcfb676edd46c7a15cdcb7bb4c5f0d0e726ab9a02ddace5cb5e8a7edbadef0b9777701b0383e2c0685c2fc1962cbef48f639ec47233f2cac63ff96eaedd20c70dd21552840c7c6f5ad36153d985b089ebbf7bcb7d44b1b61b04351b8e2335f079386e8717b4a0f9e6a920be0aec3ac399bbaa5ac492a4b0340670c7854d88473972248c9babe7acab619552388e2b3e0d5794508d00b42659c3691ef1af5686cb192e6168f9a26eb1880247d486d769007b082cdf74253a1b300f92770c324517539cac5b3b61e0e57c98cb3f8361c87bc1dc22ea718d4e8da9c5e7c98b57080a1beb284d151e29f78b9d2e9fb57dc8b88b3e3e15da77432bc59244338e90734b38db596ec5e9316dd798fa793ba48270ee53069e6f83785258cdacc555eddc0f8293be6c7551bd056eaee06191fb2ac48b0fdeeb01dece09d6069c76e0c8967d3931077154791af982e1bf1a3366776995cfd60e3b9008fa67c2df619408559c9c030e8cca271fda7d3a786db8202b79c009eefb61ca587cda7455fbd872422a07a37b15fa058c37f44a3e3968deff546af04c584f9e6a0d4ce1cea4f5535b79087ec6da9e21b459c62814dfcdc7c06222786274efc6a9ae2b5468f2c4a807e1f16dcbd0a328581993189f682dd28afc9d0caf56307222b0a154eeefd010f47c0dcb6249cc3e9782a0a530d7b67a38fb40489906c38a3bb949a914a2731a8624ab9e4bb66966e6fefa5920d0177ad2dad834b55d35b95dd1899c09ba65f9d07ec218988f23013a5a0031a4d56383bd428d1b52ea4f80ea1c03480afb80028c596639be50fb1e48bea49e70cda86d6daea0f1ba8e3864b4ab4395bc6969aaa034f400b9b4e2c6fd4cc5fc6a5658ab56314e4448b034ea0627faec8a827838960bfaf62679329fb306666d300e231092752f4474e172d94374a736fcdc5fff521bed4e87bd6a345bb864c103d5d30e65aaa879c23af5f33b47f3f4ed1470036d3f403ce263497caa7d7dd8e84e1b44c64dba47323b1990588dd741c2cb806101dce383e4b82075f741d0acb4fd039a4d174825dac8418669c5a16168264b1cbfd3ba774667b76615dba66cd75f879371049a2cc5523bbe87d295efc09f3bdfda09452f78e9c6d750b75c2881e0f2d3a37f2d4ff20b2a43172de7207bf2a1e43f884ada401eecc154a26e60e360fedb13e6f65ce072f776c9e877a69e0b791216d1f8313cc04bc23e7aa6bf7c4dca4ca34a9dd3b379ae12dfd03ffec1c89da6b1af4b52cc56f42cf5d63bada11dcfd31ab0a8466162237bb2ac81028c4d123f80c9e2f035c101c45e452c4c8430564c16b239d8c9c6ec5122eaba17f4d6a5df53bb84ba73a65cb07a4092b87ba55e0e52e5375a76bf7e21d7f79b046bc417af272e96060aaf0aaa9f7f0a28c229ebce0518abb7504d7e6fbfe02db6d1a172f00858a0c24c9faeb9b35ff5a526e2daa5c4526ef22afcdf1d810c17b41b3b7802d114f587e21f50e27538a47067df1e6c996ae6ce546e0a3e668c951da61d2f155d7a98fb46c802c6ea5080886ab4a3daf8c76b2765af3e3c0dcd6ae9938a97097842f8f627520084b78a2632f4482b0cd8df7fcd8f6066da8b810660e97b8479b57a222a6c740b6020c05da802e92a8a352205387075d195d5e6556a6f392b564d1907c8f819941b33dbf952b46eb88d6ecb6036e26c8e80e5aac36357b97fd763709033c611dea65b628c9c8ac1be068478ad67e57bd96e030270ca944e3bf196d4318825bb4a3e5d974157fd04b659fcb76ebd590f8c1f28d3734503436b2a24fce9e62a321b978169457d15e33db828620df0bb386bad6bb744d207ea204e759fe1f61ac9e982a2e4a157832382c9a7735d2cb851a239beeac112381cb5e3ea09f35bf60e7d5e277888498d8b61539d22e37299faa0f91795e78bbe60b50d733faaddb8ad2d8c5c7052b18c3a3cae72fdb972d9db56d3e2e9d2d8ecc8c6c2113b5ad1df2647ab5d0166046ecd4a774346ed0a2d0fcb243991b6da2a63d658fbed7046dc4e38e54604fa3b8d1c51f14055e08ef74f59b9f56cf54972315c38826deb2b5470685972793a59883b797cc4593beeee86033b3547ee5719fdd44339102e1f98ed6832c6f4baef1299bdd7b6a89baf49d100e1d4c4624025843cc42038a00cb44b157bd4cba6fb5dbbf32ce4a3fc396b56ccd7fcfb159f4cb3e7d1b643902b3f446abb624cbb542d80f17a4f526c4aa6b6287831a4074eede8c1030d31e49dc7795a6800dd10c3b246c77d5ef35159c67d02cda05bb13f36d799addc80cd7bb70620e8752f0b6496a88238b7e3503a11221b54a290843a7c9835ab5fd6505593c19e71974f6e817f5b86c0eb7af844db3dd44236af8e753c5a7358d6819f9fe00ceb1798c555c59f09b28aaad0da3dd20c9aab40441f8bf03f367ad8b7fe5013b0cd666d84119ed1d42d7a31083aa99f72730b48e4d01bcfba78561f2878e5ce7cc5fb6857072829f421d6ee242756928bea3ebba09ae7ba145bac723e3424e1400a629478d8c35afcc77a8f20825f34f9ab4a7fb3c717992210fd32e033413eeff4172c96b0e329f5fffd7a577b446b54205b3f802e07be32e31662417e698ab655ce6015cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd622e3557147096b1593ec08e17e0b8f74e7e43f157c42c05550ba7c51e280f752a98036344f592289fd23a6072f20845c85a7f93404542f5ee9c06d6c796c73b5025fe1268673b891245b861d17dd649f0bd5126ae8e2df0b39efb548d00f6166edf6b44007a72116f34ae47deb9f11fd478433a872c38f8710487500c1f3421b506fa5fdcd7af08a245da55f46e9a6201828e313e15b2840a318859fdc500991252a2d5a3c3152f963f4f7707b50d7bc5e41d10d70c6e626fea1a1aefa1a78e404d4c66579ba6dac0fb607049785bd7757d92d9ef3e685144d400c08e0488f6e4f22d09b3e8cb6dd6ac199a628cd29be372b8a92a676bee1585cc623e317c277728475a905330c28d22e4a44347a0945cfc74287e241705d13ce846fe8a09a8dfd163aa80194dfd017f1610bd087378f8833bded7a506b0c9f7c28cb530a63074859893f082315a117ce1a1c33d18ab9b9f070bb24a5723579789a3eb298b1b4e1c2a69e074ee91437fa548cccdcb57e5bbb82e47843e18e2844fbb91fc04c9680b019fcccd3fc519c961148dd73bd4bb5d6aa770ce769bd3e89d2d15797e4d672e29a32ebf39ec4d7d52e1662b0d8c6f289d698574533fb9c0d90fe6ce7e09f6db2098f176afbf7d154041f4ff897e46cf4eb4ecc662966a624307d02055d4a739d4e836b925691836d606c7c50e5aa67b984d29cc18681b3ab7173bda26ac5872c0a7d211c5d6572c62a8e51711340850b6a914992b5a72a24ebf5fc7c06416b91e146051f75179a3a93124f0c6d9c9a6b821ef5e03348619fc0a3615a2a2b813e4c49ceca579cea0d0409e321e0a55b96afd20fa3b8a645e5171f595e188dbc3c6aa35772c8ed9a5d4d46b18628dea17873bad989fb81919b6bd011dbd24490bb2e64d38671aedbca7c81056850d02454abdf27b52582c310c40ce1ae0d946e581a05f58a0068a48f118e80186e0376f984f262ddd080e7fbf3b08356dbf78017bd28c941c473f83aa8a780c8ec71febca2cc82bcbfa47b6bbf2bdb9284fb060f7226bd812df34c3e2df0980f9e75a5774f4bf833bef1b87190042d270436a98f4a0fc15be9263c979af4d071f2e4da90ee14c5f5cd29d11b5c66450590d9541af1c0d01e9f510260f4caaa54caf290d6bd7a87f47a21999b4acccdb78dbd5e811d022bd42a30f316e3bb76750e5b23612132885192cc195bf25fd4fe789e4ac11201eb231ac1e57e45855dcf7e4622ad2f7013029cf16b7219bca0c4e04a2fed7b0bbe40a5c33281a6182ecbd2c2e45bd7a83ea6d6a3122b0cb8c9afbe2a84eafc8186ccb435284feb6ccc1c9d760600dae38fa5e846ac2161c4fbc092e29762ea93837091e43ee01dbf4cf17ef7f018c3b053e4a8f59aea9c347cda0dc8392385da0622b69c5693f1f19aa1e4e67369a9d93c6d56ae0103002737b8e5da39ce06811f31ec68a4ba2f25682c800ff606c92c3e86e9388e3f338fca3d3855c1a89ddd4c5bdfef990515f5f7ff43c0e9659a935f331cd6d52e5303b940b585c6c1c787a82fcaa3ec9431465fbda7ebbaf02f4c799eeae6a2836c7b41c8c40ea591e01a18f5904d7b34782098f72e5e2c6d2c2ed9cc598cf01c921b5fdde102a9831f7cb1baa5167a34217ddb53bcc2232d654d2af385b2e4ad2ccd3bbd532ca2ccb65b30ad9b3a3dac8bbdfd1761e4595914c1221b2dc2125a4d30f038d0f7874a4c6f10ea12283d66527670a9c2a063621c69286bf9be30ea939da659321594ef9a6277acb0444fa7e5a4782a22a9d9404658d519f321fd8b52037cadf592a63b8b172d3a10866a2b0873163f12c926a06d2cb978fe81e48344fb8748ed4799e618ef8589366a2e8de9f8eeca55eb040fa1169e736adb7b592de4d591bca856e630b52d8cafda00b54cbdb69aebc9e0ce792e36ddac54f789f85dd2b04b602f7b4c1b2e826033ac0b68f55a7f6ba83cdb7accda92d3dc7baecc405ba222aa951d8b662c073650d304698e7632c72696598ec4e66d89098872c3d91a5a49e2b76ddcaa38b7cbc72b78efc5aba804551896d37b36031218b4c14bf81c9d34eb9021e606b37834a253d76070aea8a4ee511bcb0b22be4956938c5cd48768c5372136afbb9f6222b3a2688f5fe963f0f65ab244171daa063d6476fa8c49d6290cef0d227abf37f531e71b4c6efcae4fd862a5604cde364411d845b4fc1a7d69708e2b8a0cd4348a7c38391679b77ee7e8bed6c9e7bd70885c847a41b2f91be61b55bef7271efb189b3e29395983509bff8c08cc2d7bd0d0b206bb8e876f291ab6bc21ead1266ea2581d03e1f635a46cd50e9175a83790a68826365ca30af0fa3803ce4dcceffdc282e3ae7830dce28e4776b93c8a19a75c2033f0a98aba3717bf2bf394be37c64133872428c684b9e8ce587b211cdc271f8a8027f00abc7c7748e382b836baa9f7c39ab39bf50df522c2712fb323f5207b056381b58d58c2015ceedd066718f2830a9a06b14c3df9c96b62b72608a76cc88938b4a3d3f47153a382e1b84b5805dd186f77d1e91a3735cde7cc62de39b34963f7a396a54a3fdd0319d4fd4f16fbabab51e90a2be071554c85d9e10849228d73bbeb2f71f251765c075392f2aa8b41a74acde9331455639589914ff6b69b11f3ca4e7821e54341ef1aa56fc7b79687cf65695a677e526fd2d4a1c6faf80e93082bfeade8ee5a10165630bf6a9b406b639a5f02be47308c6ac7c74b64c19cf6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h506555527d016b1df135ed83425916d0607211ace7ce7b5b08a59cf3f62bbfc3cc1d44e71190b61759bd8e930599888b775357e2e687e21fb160fcbc7b66f1ef2893e7796d2e66981cd07510a282d93009d4326b49dc723aa4b9e0a7b30ebc2d1393e5568e82699a44a025c0812dcd89ba003db3baa02b3de45191e0a19d49dd609f9dfa0a59560c33306ed2b4b7a6abe85f42bba01462dc15c2a5a5773dd5a25d34949af4d525c967284328718931938241b8584942a65649112c1b279d93444426e934e07da41e84bb5d837b9f20620bc628c085ebfbd9160ec61f97f06e4822f5ea8d4dd38c96b0433e93a915f76d278f49c5a5d0929d264ad811abad47efedc4dd7c54c491b54fe98cc6573f787af828d1d9e7ce72a11fdaee30089c9d18c376e6aa1f623c2ea92f15003f1a00b9a4d0a76319193cab0f772de0e9367cef204097e769dac96ec232bee696af866cdd9f884461de25146a9a09123cc707ad54e5b3c0e0048c56120b8e05ce21ed94baeaf0af1d98fa9d418c5aacb29330b6f97a21285c9a1bb4099f50e3971f0066ef17791595a7e39ca64ce44acfd3fda953fa07b236bafad04763c7997eff9e4186f330015ebd6eb4dac3b56983eb6ed662e4f19405ef1095de9b6a12cdabb8954ca1d446811980e6e08e9f96d7a7b5dce16c38a0b28e92d87094041cf128fdd64681bae885be5818a518b3ca3857f8a9d1d6dc3626090b0498562a42c41508a164f34024074e5bc1066501552dbff12c3ee80afe2abfa1b372f32581679c37984cc890b6d827cbf3d08f700cd486a9c539ba829413396fd48c6b03ed1381d47d2e5ed8fc2b068be7dfdbb4794f635ac5cfa50a96238bf8a687f0d28fd569463fefc5a7a16b60c792f3b3a542be8fb72b2beb968808bb2d3134edad9c079ab1ff21f99a5d76534139932ae418d09841cfe3323303492cb2d66ad67f7c8f825fb1a39e71265a151f54a08a52308799bb704c43d80f42431bce84febc4477b7bc4eaea09b249ce7f2f6e6f343f556957f1c76bd6e29db74616263a93f09ee3aab19ccb4b6640dd7dd8fb6b805449f9b09b1ab2bc8d693b737fa3f291bf23ba085654b1d68fcace245f82e3ba296c7568c1c8452660ae04f7b8f3bc389a545b883face188cfa9034e7ba7cda5e6b8e35f58f39c249ec330644c48c0240757076e4cdbcc25b81ae8c5414fffae3da3c6f0f032a73605e1150a1278d187c1162c5ec90cbbada234a359c85a36164a17fd343cee616e9b0da2f42003ef7203d3eb13d1d2dbbc8252c69032ec3583c0c9d79a90ca4c8612ccb076f738e0759b6c1f2780f1c768f9885625e5c8baee2b69ab9d022370ba5179c53ee81fb427822d69a447c3fabbc34ea1af37aec88d152b9fcbc10a7389a7de4332fd695db8bca3c464058d779d32fd2521184e82a8ec4269105ea88ef3d9ad945358ef6fb0e7a6ac765844a02f15285e87adb30b7d77903e016e9e43d97d6997838a821fa2415f2fcdd4d09ebfe1372dc4ebb49e277e286cf87e219565b58731eca81c149a0a70f99238a31fb6e5699bc987251ef4bd8e112d98f1fb0481195d5b0d9ff491465eb704c9869808c92106a6fb0fc1cabe7f12ad8bbe12d6c2d26de382f4476ebc689cb89bb30e5ecd045998cd02d59134d5b56d6443dd1088cf0ce6dee3c8e131a51bc91ef78aeedcde33567688c173348575452f174c1197b467ca6498c0b6527cb1e8ca9ef34d46f89b33377c928137a6fc9df48a83cb61c0dd5519d4978944a4af5c0734d522d21db872085816a54c3d231928c96d83b04af4be782ac379aa3e2a28a9087d38402752b7577b82a6298636845e0db117bef92d451701fb15e577593855f0c1c5d7536d8f1637c545607b05880347f5167853929c2200201cac2d0ab61858c239fd73a50247a9ec49c55c44e90ad42179a78b59661bcb0b0e007bf8de308bd0655a2afdc9c251c1a70fa56eddf9b30d2c1cb0b7940746eb3fa5c65113a683453e63fa36d558d5dc632a6e9bfac5fdf85826d3214335fae97f7565982ee5ac575cf278225d180f6e735ff99614afaba93cf19ae6971a7eb2cef7307f20305ba4c1b93c6867a546b68efa52e3ee72dffa4635626888271bd1a2fc324205f8e96e8f3c6c071ac111a2ed3ad57c5b1875534b1932deca7f0d5478033ed1225d93fe0b603f38e364da2598d34697c62cc5da5ced3a418ebb0f30136fd847d1ab3408c06303dcd05bc3438c93788be66e60d9450b26273a826bbbbeffdf9d2e2e6a3da9ccf130ecaab70f4829a15d2a975b2ed6667006edc29a47d50a940f69a592d9386ad484fef1ca1258841e625e63a18c9c248305769990804ea55ce9cfbf39f1b76abd4f72fbe5640fadb7519cdbfe9da9d3ad128a480d07b4075ea09ad7ea7f6044f9dd3b805c785a66343121530ce326b8d2cb90a15462041d81fcf44dbb2b43ade7691cfd1ac9219e043272674653864c6064db0bf3259a50962e58067dff21e0e72100098c70199e375e19a9bb83f3f41ba4172e45fbf75269a7c9445349d931a7e3482ca8b0ab84f7cf58ca444cf27a175945966760f06bcc9217c65b349c1d8b314a2add6e68a675a770415b797bc8ab2946e5e44c4e6a879aa6c5c0621dfc23d9b1b922d7f3669565aca9a72c52c3e671178447313214a351b7df240fe2eb5eef053b1b7e0c6a8a88f4670cc88182ed4ec79f93a6b5e805a43286b9889723f6bbd04ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb3e02931f7508241fa24fff6c9a10b3fec4b84cc42277f64bb707afd4fb56151c0ac643193f12ff186204bb043c2559ed83815fa6c9f97e966df0a18702cdfb28979cc86334e5788bfe84d58238e81732a2f7a1fe32803c87da174f6a2f677401eda3b7be7a9e03b7ce148d750415c29290030d954496218c6bcbf942759714216128328f17bd29b93c073e754d555868f54be5ea27e58e5ac2771bc8b9005f5dfc27f3fdbaae779fa2cc1b1259f4f191a83804b87a840952d22ea42bd4d97f0ad16954bd91f2ba11bc9fa1ee1b2d7c73da46f0497e138a6627087e28609fe83fac0fe330f99dfe93c8b4e8526313e870a7d8abc3a9f1852f4d7d0c90b852644c8708357618ff660a6cdad72d76390cd6ea0ed6a318b54957863383bfea448d50991b01a7cad7b0ee334b8b18b6d1833f4f565835d597608f294ab6e4c5eed021f63e175486a796e9e263fa45003462c0c61c38ae5b7d836b0f50a91c256f0b046a3a7e298639cf395e4a7711eae197f5e5ed656cf27453c238883276b48f8a70b0dc01e5977840c213f966da87a87b432048d7258afe344551de38f45f91d721c09b8c5193d5b5e82c8668eb569582e6213405bb6cef6d4e3c3bbe58a82832dea59293e62280755d6d309b4f3ca119d11111f1bc67d8cb274065d64ab780240b1d560c4cd63cec04e0ce07698d5046e97731fc968530a03c7bff55588ade8e2d7b77be95c8004c5a502f921b5c44ef67e5b1935a9261547158e0d89700baea46518e7f03416f5aeaec3cc4679e4b91411563e95909dd8ebe06af0092fc2ed29c005d53c2a84cd59766f4d5e85be61dae16572e005ead5f22fb99fa5fcc0885ad14dfbe54c2ff9581d444b86ccb4947f662db9ea8dac1ed83c6f0d64327c151067fbeffe2309a5242650eefd23c45b270c09655592927168968c53be4c701d40ceede22544e123e51ed55ec880809ade2152623eb1bab5fcfac31c0dcf40aefa784e83df95a89f6de72c238c1949fa0cf682b3e3fd1ba95a5f96440570006fc98de3c7f75ec1cc7dcb777584ee6bc1f80f0896296bf918687001ac264abda6b6a4b778b322e74bd27697528d8226b56d5a59078407fb656fba37fe7332d56827b310463074b8e3fb2af1d09f9dea6afdfd794378184963dde150530a10e2c133b2b3d28e2469864944cee7d07c16e613d4ae6344d2fa9a8da55538bab1ae1998cdb385b6c811d4c337960f84037fe84dfad7b29f1a29dea186df755da66e5932f65624958cb5ffb9ac663a11ec0ab820b13fd61d8355c53d79380de62c3694110df2eeecfd6935e5fd6d3a9586af0f4c98ac09627c672dd30f1faba7a5ff1bfedaf5b360546453f84b8dc5ddc9f43ddab63a9ff75a7c7144af3362ae05ebabc6bcea2a1df0abf2e3ac2398b1d2c1dac40b2b295455494e67e2afd9972f8cd0ab7bd3cee8797a11c5e82d202b65f71ebf09e8b9b1a884cadb829a6a7d08be364dcbc5476a992b903fdf03f81a659304ad004c01af7f3a07c06584c70ee85d10f38d9d2c76a24691b6e1a6ec9f05beb26bf84f90a31e753040046aa33a49519594745306fee95e89dcc81b4fec36e839371900e34d2213cf3fb575cb99b2bd3551c7dbf52a31fba4478fac09ead31336c9610d328e8199124dd93d2a59531435f098cc52df2b83792daec6b74ce2ddcc07f1a55d0e6b270306d94791984eb7a8421cffc133cadac26f3872a14ce5278f4cf0b67920e7e57bbf28418a6c55b065913b10fdd253d47d6c7b697c625c9a317f3d8c0f0d98ba86afdfdabc3a4df496900e14fc6af4c55150bc921ef8993ec51dde1a678eb8f320c5ffda5fec78b4dadcf58db68e36f87b517f3b1ccd2894a1816483e5bb238d51260757ed85308c2dda294cc8ca3c2e306f4c05c27b418116d1f75248afec36281a3afca17d922605a7ef47053d2b55f41e8ee449c99708aee3b533d1b291c03f673dae2aa32a21e0bd599d63e059c4bf28dd41d2d1ce386befa3dcdca01bba2d337bf67103c69b24386eced9f20a935c03e6d86c7830af681214688712f8fdd9ba3f2921913aa45834977ca35dfa67119bfe93f95899756c970077643322ac8075cc888cfcb566c5500baa5e7e30303f7ec6c1e8e2fa8242a571f48ae2eaa91fd06adb384096d0b8a8de3fa96786025e7bb6dc8579d4273cf59f4c22d27d81da55069da5f8a900992dbda4497e608902107e5cae1029d5690e808a3c9472c61ad71c732e1c3c8a7a19aa208a1ef05b4233ebe8690dae26dc8c8f6208ab6d22924c627a3c27b9235738d951327afa0886271538a5877d6e0d4480d209d11b2a258d90968b5b6c34219d0fe3983029fab8911f5fd1d3fb75a1166623e40825a673153e197abf7e96e8478b802d5be2438867b39b16e5b3211b1d4ac9c79b0c14f9ce524eba03d530578cb985b21074be87ca1810fe50f4a0ce7d8b834ad68af49a8bd41de7edf4489b85a648a8c8f46abf425eeacf592d0586a41cc568239ad47d659af616b9f48bf914adc81872b546ebd9d31d8376991251cbe4c18ec98f641521a0a20ede54fb0cd186f889dbde80b1ab0573d5d8fd266f4750cd4b9b5660c3c33665eb0b461db1070d049c78dbce99ec7e2a73dadcc7443a04f983bf47a1c7d4631ac8eb8eec32b5d2e8696ed1dd5e0601fbb0303eb2b82d691f820b49f7f6bcca7803adf2951706fd7548bfdbd36d990544e290764f4dd253a482e091b29612;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h66c9487362083518aea5f534bbeb1810827c9b392d3dd3ade9b5ca557e7318fe266077968e8802d1c167a08c03d2a1944bd71ccc5cc429038edf9a195022eb94d68bbb02c88a58ef0ad2cab09b00037d71a5ebb67cf90a04a029d52090795336a7462a59c98886ebc14f98946761499cfb1639e057fec0f75766ba871771b64a0bce9e287f906091f19f48bf9f8052e0c6c4a647b2921bb1454d74f25fa4e4aff6bb6a36cbf3a6154599f643ccf579ffe0e13f46e4668a3d48f39a10207b323179f9d7c6bfc0303ca9a213f59c147f60356eafb6cc528fe6fae241d75cdd68e73c2fd7d5f9f245042a341cf6666bab5b11a28329c3e7f775707b7b5090a5811a92439ad4d3828ffb20394ebf35e09b6db1150f4c9c6a7e87eecaaa9ca21ecc14854efd39e89678184f9f2517d89621e1a7682bd84248f98ddefad2da30bedfada2c9e04e6973b5f87c00627e90421137e383f64572a134d94445ddfe81e2cdc32cd8e2b0d36e6de7143363b2d05d87131251da4891079ead5b0b022669cce30aa02fe2a851703f15571c574e0f980b143eaee85337d7710e66b6bf2549b78f6643e7fc27f8e776771df32358f9166435e2fb2e2d7fec7b821ffa13e9afea8dc847239f0e5480d98f6a03d301ef11bd8a94de8f0cf6872bd115a058122dbb31c6f6325d8e8b8569ab5fdcb9fa47c4c6f67e6adc0e65d51b27104fda2c25e5c7e7a3595c765efdef050134fa9c1df9b69c75d0cbb987e6c874c2cf62551bc7c1fd5957510adfcae870d805b8d0fcfa5b9b9fa1ff639d65db01ee2a89efa821d37cc4f6784a6a46c413ee1693e283d87607a76e8b2b4cc45ba7c039b87cb6fb1ac5d4d37ad4227c2eb10d07f7aa98b6a9c30d25e7d33038dc4abad854ec533fdca543f9995ec06c72dcf697ed1defdde0b851177fd305766ba7a36454cb08f4445833ffa03be9a9f3733b5e5f3bd265ecbc72157c398ff147dfd176a2b9d27492fbeddd0db487f651dd9d09ac61676126ab35e87c29861459041a556f7ac2f219d52218e501e158a96d402ebfb7b17d676a88eaff2a5d814f7f92d17a5d729e4e336cfbbd2e4a506243c66a785ee930c3a8c992188dd9bacde026ca5133cdb473b301dd19cca8de392dfc2cd6fc67dd110a6382f658a5cd02de2165e91fe18fc3ea43fa49ba861ce0d66da339c4aed16824d1fe11ab7e4a96714fba23955e19a37bd1fa23b738ade87523cc5519557119b5b99ac9d433562e10228bc8096c014bb0f0ca996a99d4fa0b86d20b14190a05584b4e9e958d0973a4f1202054b6fa6e3160700f98e2f95d064499a421c4d805af0959e990d97ecae106b88dd42e53acb14fb1679a2ee49dbb61b5318d36fddc0d3a7ba5ba1e07fc2e5a3e341b7d14d5a338d69c5fa4c368e5ac2c1124e69c14666d5700afb54f8e600fe60fd613c85075cb8169473cb26b756f46ba691efd162b66523f862b6d7ab4499f079810b7be6e5999093a4f1e3f314c66e64a9d989a51485cfa3d3a54d553c22e91e6565a65095d466a7bf40f31967b434d5b1846e967aab389c66295f6d4a8d397e009a2b2b0b9db364f4a83bc5cc920669df40efddbc641939d587a3ab8e47e6d65705d8216e2399c43193a61b6d6ab06508ee495871456016d0eb4558488e6d32fc0f2a4a61da0689b3835ff0c8f87c537bf7ad16cfd431b4d84b7a12520f5f3bba961efe40e54441a9aaec7b15d8582da2f53f98c492a5f4dd6cca4f477a42d4e490a1272e9d7d6d19dc2796a72fa14586179bd58913bb6380a1ff9f402b8babb66a7fb95e2ad08b3ea389af724ef2f8527c704d3adab88bc47d3a01aa2bb7ba6d5eab5668b1cf7d99b0499302c77da5f3a0fa0bab77a8be9cc40b12bbf873b8242cdb6159831f011cd2e0e245d179c60e98fdff6d8d0d8f6839e7cfa47467da56dbc411bc7b3320fda4ad6767dd8cd33b0f17479d7de3db0d757cb811ccf23551edcc906cb4ca935a76313036672d5b304585ef22c4ac09b847348a0eb0580ce93c39fe3862f10c8e9663e481545bb66fb879a76888d1dbb99842a02d78c49c45787e37b88edc584ca280cb6249943b2e8b253674cbe01e1ecf1552eeb1aa27828586e69f819d98dcb8a78f292d2e2b0eebba3205aa81d9184c3e09b8e39d96f101fb1f2813b94962a962e3da93f4ab61dbe8db97614b7e4ea7bb91883bf2df8601b6faa71997ef215d02f8b24f31e2701a69be221cf780f14c9577691d0d35a4458e7250fcd023ae6e4a72a3b998dbe882828c2552215e47b990899b627e0dfa76f413f54c93db365b4912d349eeab17ede014ea7afe3e99545324a0c1e6d1bb677d8894956d1765e7fa8b287d80d5a51a1fb8738c2891965b064a04361d5ee099207491ed8d4d3e3d7825ce3de3495bff08602aed5ab54e45a64dcd339b32bfbef963e089c9088a0d63b5b425db2098b7d08a4c4e41fcdaac7212540677e5909a0e443396a3abbd94ab1845626792ed44dd9d999e635824be328dbad6f33c22f11a39d70b3ab0ed4086a9fc22e5a3dcc0dc73b27f9a65a0cdf72f0e54e715ca8c5323a70f12b11aae295496f9576646c966f606308aa7bccca8d022b9f7ed2792c9b53917fa90e52a3b2bd03dd26df09c37d4c14b8d615efabaa235037dafdf85b0ef44c1f2695a9aea404c65bf0fe8c53460afba3c9494a8e9822b138f87115e97c400535f8ed324232195ce6b60130899407f32f0c42c7b65c1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h12fdcb99b328af80fd09e7f30882fb718c717a26c5e59c3b5671bf71a5596a3f345c3d312c8e952c5ab0a908533322cfd18e0d9cd89e52463e49cdf800ef5d67c62d10df9aef69b07c23eab0f5409e079a4f373b5b1b8d3f1f5c777d3bf876f4ba665a6c284efd2b3b470887c2f23d2518d8b4030eef9064626604b926371c39f2e4d9e48cde824db9ec3f7ca6250051de1b1ea2989d02bdbf2bced35d99ed08694476bf15236200af78c44ae065f89e02e1b58a1936753da2fa7ad26abed9bee62b37602ce1910da9fc95216bfb282e30d269c24861655983b8e17fd11cfa71f023321f0755d16bbb7255182f86dc86365a3b30da453d012948264eec6b4a53f7c9b24f710715a7ed16336e58cb616699bbcd10eb0631366bfbdcff4ffcea5cffb5cdbd6adc73bd554fd926c07cb5d26490ba90568cd995b8885ad9698dbfab9c42807e2952a537ed67c731982909afc13c4256474af5452e63e038dfa1014d15b15f453bcace08c6bf9ea4088681d9a088b4cc66b92883b71837b58707d008d9f927a4349338a01ceb8133813befa9a42ae8b9706cde25b6b4d8c720236da9b9e59fcfbe64bd2fe0230e618130499dc6dd1a1018434e4c915952bdde39e3e419c9734aa5c372ff3d640463709d6026952ac4442848ed3e4f9dde0c0f0ff833a0b1119ffea59d0e4b6c3d42b1c751310d60f571d7017061f2c5995414251567bbfda7476960c0ff0f1724b5a3cf1836d4ce6fd9202c17566d77774c9856c6256e784933be4462eb63387992ab2d0948e58afc020b695315f3193fcd117989a4f92ba56e10b4e8dda89209ee08db382cdec64e9fadda0636cb6de021d19a0e007d972aae1a77d2660f9313478e40424809fba1133881fd8b5f69b381b463e43a103c7ae49188ecbf0a579cdeec93e5e44bdf21fcfc2205c82dbf4dbc2f60685fc08a9bd5a2fac3daec2d529124636b3d4c53bb3c1fca11699aaed95fe8b76e0cce921cf43976b788af000fc76c7a7af3900f13814528fd04381bd7c9ed086122227a9a71dc8657cecf85f5a776c5bc591361d271a138ba62b20c122a2a1b57516b43631d6d4720f2a5d1bd0ae96977002d306a67bb8366b0544d456f3340fa2cf8d437c1c3d5cb20a693574af01b55637f6f7a0967ff1ab7664573defcb0ecad9f319c522ad1242163708ac852679ec3cc7b276296077b4d4768a3ec52c52c2c9db80ad45169d64abe45e5dfb4374d7058598c89b9ec0294cb9284e49a29ff7f4e8860272bfddc99f0037568d09b2d6f97907ca6b59af3b614d1123eff645f2f0e6144f65d420886f8e109a2c07f8c0b31f008fbab40f887b474f96f81ad74ec96049562afa4e473ee4e81b26d7130b1ad07ab943a70199146c88c92ec0e292fdf3ed514c466681eb50a7cb4c4173c692d9e19b5f81f294422e84c0d1abc64d1632557a27b8a384b2d4c0495131fd3b1882c03bd5ae2564931ab35a911a3655b912d9a005a0185eb195563c1245d3b11e1dfba66808662e41a1cf0307a59e7cd6a99809fd8ab8971c7c24b5ca6e3c5186d31a5247674981d6fdd34b453195bb8f6e6c33796e2531dd561226d2065044f8c970b799d73dc33ba1dfc123ea6e1729e5330436b9f1afbba4b9f7dd6497a322d339aeecfc0c7a96402f76a64f4a91f54cbc25324a7bb4228369b6337db82046e61b33382b081c62138484ba9daee284063c01f641e9c48938c46152780206325794092397c710b7cb3aebd0daabb6321df398b3efe0c8a551a72f2a6e7a0757857ad5074fb5a2ce5c7ff849bc4edbc14c370a77510d970d11c70c0cbf049e47ac3f5e8ec41d313d2e4301bad5abbcf3f8b4b4a45196bd80dbbdc1d0860141540e91c44e2cbe22b6b02f748264bbea7400439039b6cb1336af8922767d5e8317788668ee42906e78b66cd31f6e8f8808d137931a5221e3d2c050e3b5e951f4c09ef73f950530751dd8ca7e91e1a336f80f6e46b6ee76963da8ccb2c47a997b51810f75848c83b2b84742283fd9a1919bddaf9011246943fd6113d726d013ff8aa7331a597f678ed07f90846973b699b6e0d8134f87843b67aa32a77cfc7ddc025620fd6803f3cef44cfaa0ca4dfa05ff28bfb780b1133ca831920a9df82c10dcbd97cb8eba51a7ea9c8c87ca1c34068954c00e588786e0795ce829c010dc0d80c25865db0cea1dad47f6d4feee3bffd7ed9e5723d11009d4ed5ffec89463ee89751fabd34abe2adc8e9687adf0dd8a80ddd2c8fbc15c1620ebe5b96de6d12d037419f88a111e4f9dc3010ab907fc72630c161073278ad1b02e6a6c79d2829a99439fcd457076d5897ec4a028bfe857467082a99d2c1e39dabd4e7659cb871ecac54c647e285c1b77bd0a8f22c7814ee88d707b83cc138f4db773af25b7e042c06919d06aeabf9962949d4bd3cdaf84c31bf04690179412be8ee0cc98208422dd37d533895bdef197b83dc9183d0d422b91b9aa02251e4584fb540682cd2c7b4063e4a3275084d9277affe2dfcee80207de53f01f56b779d54a1a0dd92d06a1908d2f21a1e41696af695f3676ce0b9b67302fce1a554298ce2fc52cdced51f8d4aceca322f82bc3000e4f848b1c9c55b526e75455126a1e4d2cc6fcb455812b06560228319010b2acef7f5976605f009715676043859a34f158490f736a0d456b10e96416729e40096175802d0ae4b896ff3acfc47e8b6063b8f6b02295b043eb50d03550ee1e333;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6949be238a8e37f7f774e67760c7f2ae54a808fd21ca9df299e49660ee340f082166a3add54dc26ae860e748f257b28ff1d16d3fd8cf4da2f8cd1e6f031b34638964ad0af3611350f7e21cf209431eb16cd0bbbb89b6d0740ee45f0b8b4c843a344ec6aae8c0fbd0055daa44de95c063d5c92924381c4cd6f1f2cb339afed245cdd6d2bc3f26aee0a741199dc8dfcff4aaed808be1a08523a45c485c9fecda53866f167670732df5a7c86f20b3da75be3ac88b65944ea0109f75ef190241b97549ed00218ac5b23ff8f6eed0d999009602df53f163bdf1752be9d188424299d9c0416b14947ba6d328f693b1beb3541d5028323ef645ec0a6e1a02cc2c3c2bcf92395d79f50b9664199cc5f4fa9514e7a9703799cd784e5dbed2877a96e0cad82623733e9553e4caa41ffafe025f369f70e7d122328a114ce3c4d87cc25413752768239f6e0b98fef4879a923b7cbc9c3a861afab92e1d7fc24ea87101712284453289ee673494fe9e80805708a552e8dea23960feafdf7c7febcb43f4b73573c0f9f415bff56362fdc1337aab456cc13094e4261da4f59314c5bea0ae2c37b51b63c7b999ff9e4fa58beb0d9ac018af137ac0fdce0b2ed15447a81209068cae33d9ddec08d7b599b27b8daa411fcc9aed38ab1a59b20494fe3d0f348d1f0ee8dd5641b11982009f9d3f6153455c163338b9082d26a00e7a5dcb00702397b8739b11d9f2bfc28ee729f21c2e527dd124b90b3a6ab2576434279eb5215abf63189bbbdc060762089aed9208d316d9220877ca890e4096e82d67ba06980cb0052f1c91f6ef8539a079a99ff46e6aaaa4e6f8dd7795f82bd43e543fdb8aaeb93cca72d953bf20234b78a68add54c818bb4d63384a3ba763d3678999861e16985f1b98df93d2588a00a5349be96f591077273cdbf9e360184da4b85caadace77bdc24d2c31cebd145e1d7ca246f6c774b05749486ceb9467217c1f554655ef7f51e2c18ac5198aa962e48d2ed716ca3a6f4a52995fb1a09f02f519e2e2ff9819293a0367f6544650c98354fbd5289dc4254e8b152c93cd11a8ecc4a3474a7a1a4dd25e94a517845daebd90a8abd0c1adf2ef9bfd1535f6753e8d6dcd45466f424472a2d41eb250f8483ba2d37d27efce078322d7d758934ef49fa1a45239ccc144c3397cf15f3c4f3b88b249a4ed9dd07013c2d549134e97bd5bf84224448b26b4f9f3a1cb4d1cf5fc496fa7f77374ec2d6ee5aa8df453b1d76dacc1fc572939f7a8bf5ffe4e6aa4a00e0e6c27cef3db6dd8bcf24055f7f583f9ca3109121add21d0a790900abdafab7ef649662384c7db1e1d11ba05f34655ad6cf40caa33692886f9a003594537e4ec928ac1fdc14f75259a112af8e4cb98a9fd4f675e199c0e1ef8ae7d273424b756368f075b05bd382ad6845026211b89f9a35e0071ccf6d62e91bf4bdeead17a524fa8425a24cb35898be0af63f839de0e94674088166673bd973e4240c98c51d240a0ba99bc3f8e030c473b52c28e90fb4ec9f605b5a086b71e3e3062553cb5e595407ccc69868dc5e27f81a6464533df44e38f3ca4e04c23f400948c975a3cf9c62796a2075bb7744e324550dfe4ac832251810883678bf14e85a75b32b67590a6994f18b8fbfb7ae4fe3ab34a3657e9f31bdb766323c3643e9876483624f4e9cea0f54811e4c6800b1451513b15447f7482fa8531c0831c322a8f02268268ffa2199268d3c264e8fc148c38a2d67ba1cf75d9a994edf9efa4bb15ad2927c9ab9bed60d04a4ff2b30724ab00e684b7abcc729f3990af838befe480463c5cc5e29e68223fd207dfd4823cc3322cc5f87651d5896fd69a0b6f4469bf0b7b1406a4ab839d5dc529b09aed6b802776897fd40e5bf13f5a74079460226f9d4001ab93398080995892a293f2b813087a8c3fa53608dba09a9c5e53b6f2116c83a3ea81d2143595d3869d70f9ef23901f7de2e9352ebc14394da042a9f2c4df0a630cf22d15b2c352fd046cc52df4601e75c605278d81925c58e676bba5566ae3c5f2ac7f62374b6ac101040dc1a15fec4fc9bb64b5358a7fe799781eb4dd65d8911b7a25fc200ac2be4aea286e6c77f132049f20df25d0438e0d266ceea0310a24200688ab83aaef8a7f89d569f324e6f99936288999f07bee391681af94b853f50a798315ffa09c1a011374be3f140c61f66617b40abe85a10b28c2206d1fc45661d3e9f016c52bf4e1bbdb7da1a9c896b249d34934101f4079c6aece457cd980eb6861100e3df1d02cf1264b2506f7994228ce4d0ef85903f5b500a918b80803cdf40647cf020b64de162ce5bc343f04ec5450226fbbd0c29bca08c49811aaa1761b51a4de787e6ef2346cbe0c4aeb932667d68cdd61e5ce91069586cf7df0c674c000dae94e1003b34f7756722453a10177ef2d8e59d5975b7729e6c9caa9028aad2a5e8630247a666436d48a9d000f4661d32f2ad13bc2af171c2f51177c4bb8ca538380e4c6b864e97f626941152d039f24d21ac75c978e15f5545b514c8ea00b2ebe0dff295f8d35a35ef3a77c1b82a8e6f0038765c2428c5890c2a89564235208c7b63c7a46b2ad812e27c3daf5e2a39515d17bca59ad10a9e3f57489f350fdd8ac8ec393be5bfa2ffe275964c890d3ab170d8571a6a6b28a74168d9c45dad287eb998f9d751b0a0e896ef8623ecd09456fcc93bbb3dcc150f68b3647ff8171e73e2fbe414f66c9b0e86a39957b63cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3bf2a76e88eec27fc27260035e1ff354d89a7b37cb8e1525cd75f45efe163267036a85d327d54c1735534fc58b6a76308a02bf69d89b2e5800b502aa169f46d476280868180944ff98463143429e0f20d0ed07ae5324410fb3be935e02892d052c7532eb51f5e226a6224ddf6c52123d1e1a7844c89566ec51eb70ba885fbe21ca5c88544e538cf682bce07d47f5a1ad42e72ba2e1e26dde020aab683ef0c6b3a04c7000b0973f62a90708d91fb6ce9afedad94d72833adff6fc47655264adb734b05a35e60df4cf0718de326dbdd6c90d6d082b89f36200db87ade437984622317c8b06ba9fdde8c966b582b5c131ee09ce60f3802bfb645de0f1f14f07e1c29eb469edd167672c09ae6abee102d42f0c9a01165ae8b744c15c14765f2af618dbec63ebaf90f0bae4f1199c1dc2373e08fea7657518d30c7359aa43391d21d5ab3af9432873a08a7ae74fa6965b1a968576c444399cfa381f66126620d6f93ed341f3f113e71b7d62bf6f89e53f81a1e0556ba1442b7aaee8a61bab5e108d6e599e461ca78021884e10f476a58e4018425e81618b26877d741e864b46563bfdf30812f23aa19ea883a4b6048ea109e1478b40769fb6846b03609f99b1d5da4b5083153c3edc2b5d334a43b74519ac4af6fbefa2265ca5f1a774f767310f6bd5881cd18d59f3c5495547246f58ee05b85906c36454a8be57e79953bc13b51be289fd88f38ec4ffa55bd34033b60b71925c3b5373f49f03cfebc6154fd4fc0768739b7c391a7eea324ca8e817308018b0c6f00dc3498f322b6033a3e6c48a942552a7581f6d74440d127ded08083570cacc70d5dccf1f6586eeec21b16627752616af885fb8ea2492d9e116d1c830463a8cb5ff3933e7ad5f33141a3dd66593640dfb60a3d741dd883de9a36efb3fbbcfdcb640d39a8b9a00cfef4a13e9329aef200a26c984e4d1287a21b3ef90ebb2f45ed10d62050a79b85aed1f643eeda6507c4a573b4a6e08470e35a0aec2a2249c8ff8ea2fdddc549889d5e794dfc6a517f5ae6592930d2218ce98c726d671b67a4f556ac98f411fc65d8e0432d647a798077bf903e49ace70c064b7ef9c78e79530a5d0b596460c1e5a97be1eba7924b920f33e966d962a25b0bbe9fff9300c992bc8c841ec9d195cf36fbf2583702c555da54c26e360a1ff54c99a22b0714982154c4513e4b509b17a16eb6f5f03c80a5649f841a0614472bc0ba92f6116d0c2619c9e71dffc58bb9d3273ab3602a55391fc96dd13a9e10c703347d492d4e6ffa003c78a7f935003a8775683ccf23fad0b565011262119747096b34ef500224169d2602deb01b880376b69fd0061502579bd060cda9e449cee487b140810ac5a3df4ed25491c3396011b2eba6791fe23451dddcd1c1d59891eb1f6f56923584b4d5ea6ce0ace19202b3e7a91577bf5fe86287cbe955cc0ffc7eeddc3c945850a70da29b4d8e9acca997cda84b2e35ebffe2e6f316501d45fd99edef38ca042b66b427f4c07f2a6bbc642e0c24033d9041c816d67a2effa37d2bd63a6638d4cac7c8fc53ab6d4bbf7ed42f5607d352c8cb333432705cd683ea8ccac35cced25f2aa3cbe42f9d93e315ac778ecdc96aae68e1805e356a8d247853d02ad13884ac6bdf4f4f1b0be04a47ae85635436beecae0bae6bc17d92dee215916e427fb0ad7213b1efd085c887f86a3f88098dd457ceff50d56947e825f8bb87c53cc4c8badaf96f37ef8550ec46544e62d59793f3ebc361fdedcebc903b6a5f967dfb2aec3beb81ab27d53e2ceff20a09e4a5cab959f785f5fddf3c94d4fd52d77f40d4408ab33ed42ed558c1fb113b86fb5ed7e2d0a50b70bbf02eb2819956dfc121fddf2229ac292c1e2a310e9e292652eac378c0abaf9f78b1b34966b46528c8800f47c2cbbf7d0bda16cc1d7432571d0136034333871ce0d6d2b7bfb354613801e88f9fe84421f6e61c43cf5aa727ff6a3143b545c0391eec7d824dbd8861f20a34307a952cfc1bf012a3a6f9f19e54598a34162746aba83325aaefc6f98c2aff49d65fe938a56c2c06d6fae553a8b10edba99a8967647c4e5b95bcb1ea7e382c29edb0931d5e68bd62e6cc7e0f53177d1dcffd2cf4f6c155167637afba3f3ff95b46f16eb0b324fc3ff88ffce39955b089a31a59c910f56547bf3c324a78e2dbcad7f94fb7753d40cc4437e2a5df464d856d624805012f864b2be16b5b289a79d65ce9344eaddf9b3363a70f5e18442ab6ad7140b6281a03493b38bf1b648620b3e036a388021af440388b7ad996058414d66183f96611452b94581634d556f337b7d7d967074b10dc5e69fc6b7432b137b30c0e67ea1b932a7e732e812649e2e093620de05d20105a7597a30e4437f1caf629c4cf53f37d30df99ec8b203cc35e55e962f5a606474207e2ec75fd2d1b7445dadfd511cffe9b03b74aaf4a107a417df3d77ddd255fdfe7fa335037c9e1bb7a5a0134bc230d36767814734cda2a669fb967c3ba754ed1e90010a2e8b8cb7a74ff003abd7f12ed4d89754941f844d3a8bf61f484294f59b67fb6b2685e7ae759cfcdf0834fc91dc7eccc17164b110cd42b6ad9db75a8a2e78bc2c850c38d67ecc03e54616fb695a06b847f21c0b0e7d37ec519a8bb5be7ec19cc79eb70016882b1aef6b98cf23ccba6240c4148d04b7ea301724478cf6b29ec178529dcd7ba1de6a4be33a743ca6eac9fc6f15f795925e97554abddc275297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3bdfa43f9fc61f203aa143a3223bac9a40fee3fb6d6d7ccbfc5e495187a89ccdd4b3742ef963cbf13b97d8f0401ea5f81c8f2d4c4105749992999294514044d73ad2971645b85ca46b42cc9a3566ec10527c2bbb86af6b54c6e0af7478b77af3379743edefa5b342aa0adab0d48bd3a5793b0e85f49e2b787be21619e543b3a0ae3a948df83dadd3df043c1480ba38ca734d15dc7e0ca16e60dade80f0ac90471583429f8abddb5f4b0bce1d15119a4ab6f7b9c4a8f4db1d38f6c69bb42a5df16044020f638fc96483d085db9518eebe4198e6dcc7484fc97c2c3b30a7b990bd3d8404bf10094c6df23463218005487415809615ca52ad0ec8f7ca6636ecc330d437104e096dc244c265a86bf4aa6323899d9eff66490a85267e77e62d8847c06bfe090cacedbefc6b113f8bdd79ce5857fd0c79645d82c154eff058b3a9661b2691668ab8ead48a88321d4a256fb40851a545f5004cf3ea0545d75e80250689ebb13c7c7cc82df3f53cdc41ab166554a412b924a0d49a8efa540e502ed58e5731fcd71d3d7dfc26f56569b4045172c2dfb2f6d3d02e88e5e10d8500277eb2af0c8e14fa7302c9024c745c9e862efec742e4084c067eeb75c9da2032f874b0a00e1ba84482012c2235bc2b04ec72ca6386ca3c3753c7f97c8c5c2b1c09504c87d0513d984d5f2116c5c756eff7942380fb482a7ac08b81e052c0d0e7d998efaf33ba11398a79b80a1877b4e8d926e7a594f5bcaa17afaacb56b6b486c5e9906a18dd4446651f097f748e8c709457431b5c3676080f5b736a951371b20a951bcc840750d7d043dbd20036f770f7ae604c86978c881e643838c6741bd4a1bf245c382672a996d925e7297beb1988466fed81c647712b5fecf847713b0b9d17ae2d888b513c8c71ff3426b79f0fd5057540015e5d84066bf12d98bfaf4faea98c2099b46aff0d4bfc4bba898f2f7186b34cfc969f95ad619b3e5eb1c01d62986503ae8fb371d5f48b77775993ebcc93063a9d0b27938338f73c777e75393d778b7c3bd428239c89fae7e18057da1a86a6c15f235a158421c5b2ad8a9f5f80ca22a8d98da36b91a2b7887d8b535e2a75ed86056f6a10343fea2c405dfd1583013dfad2c849f375e59dbb8cf568be515db7daa1a514f98e743674264c60efb78635be89a2b4466aa88b1f06a8bf62c7db0a48a55304accabf2cbb042ba40fd50990e0cc6899bbaf8d848d6ddef98f7e17899d79be836f78eb2189135275bbd05aa7bfcdd649e334f0731f8e2c7c5ac3ef3f9c8f62641fa0da75e354d84a234f4616a3cb22d57c789dcd14b183774dbd0fe59a67cf97f20efe64a183753d81eeb752a245953b9470a5a79e933f1e960f12219c63e8ad2df205a7964b2bc418fe8e3ec47085ef8d3fc9730b2d1774ecfe40407f463b7909e9d9194e0ab466aa4b1291392209e80c91203d144b1ac0a7164a687df76bf24e4167b4ff011ee244efcd5f5ef867800960c30fa94a9032fd11b39a8edea2237f19f6b6ba36cd95a7081da6d688fc6e617d9bb8395618158e2dbaf40576655bb3560b3fa4947956950b250dfd5daff2fb03e08c62de2a679deca6d9d9d4b15368bf534e0367f6c44408dd5a0c6c92d1b946e5e436c41c86168dbeb5f9d826beb6b6a403f3581f4424b0b22864ecc45092f11cfe412c1241a2fa67f10d52b17171f45b9bd1fe2c11c2e8dcc6d830adfffa37b33fb332e2d92c78e3d33f2a885ea7ed113b1daba0277164060e168da9b631c325d575367dbeffac175c442fc2670b218b3080d49bde5b98d121510a719b5dc9174c060b0a8528aff6e8fd8fcfb0bdaedc502fddc32b66914a39482d8e66adb6710b0ce04b063c3a0aadaab81e3b516931540c7ede571de4bd91bf53dcbab51be0bec22be52667abdf47f08d6ca13e3157739bf6b4985a747ecb5f304ea8974b1e376394ca46b898c5996ebff107696d8606e36742a8d8abdd441e5b76832e89288cb00e284280b2d6e0f6ce962a7e3c37ecb2ce84624b9ef1e9e524af8468a3f460b6afddfb2a87d6e767e4e9e1449347ab0fc3471871b5df853ef1c6c225e20c076d0727d100c5f37ad68f39dca3b9a64edee3672b130b88f4e9f8d9b074560f68ed0fa9c4b141ac93f0109c3ec0e402e47fee0e8d24d2a88a251275237e6c7e144f33147ea5bf1817111b9b4ac209f2e24eb368850f012fda015f67ba5a51cbeccfc48757ce58b91c60ce431a60c5f567a7606013a3101419716af8f3b94f24e6c63b2ebfde21789c250db0bb735cd597a647b901a76d52440b3fc097061f1ea043a033b02ce95a20804349cb06768f189159ca6a57d5ec2fa8be74954b4a6c913acffe1807cb7f6d91bf343310a4e841c39fdd5116790ac85a57f93620d48c7c261e042d68a1335ce1faec21518c46acb50a68d729773fe2a0f794c198f3d200d1891b9c0153bb2909301401a03e5538b2d4036741717662fab61b6009cf79d4116f29bb28a33fa8ad99ece8d639ad79ee18855c6e6d156486e0802ca72355f83b867017aff1a5562cde24b9526a0817b69c095729bc681bed7dc5398bc928751977fd3a153d2c0b07048d0ea1f7a5655696035de53880d63d8cbb463c4702abf17037f5479b05e41ff2481bfe246649ef8582a67d14b8c2f4515a657dd79a2cce36d383239bf6442c92b876e4596386db25ba218943c7e800b2e72721ea7462253ec306f4f9886bbcef596d19ed697ba9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hde67ac20ee6867736dd036394407aac319d0fbb49eaadd6722d3b43a10ab629193004cab085ab0cba3bcd0a6bc35fa605cb705c471c7bd58e01b23c846edfe67097eacc8a6c0bb9051b52f534f9bd180eb472e9b7b3fa9592e6d5ac721a4bb2e4eb33ffe6ba631b1f065555b0cca07c878fd42d4795371198a334789a052359ae5330951554bccae4315267ff98f04a3e7e1b20e9838013a474d1fd5d403091e03f933cdab844da97ddec409e0485c25b2ce824261e05495de4f6c7af0be71144a12894a4726af23019dd8e978584277ee47e596c245b983dde10349f9a739ddb83d3e72456b758cf922e08837151cc3a450b0b3eada800aa287cd3d840ce6cbce9a91e97503f09ed41ab8402cc3b67a042225d34e2dde0794d8107e73b00d56d535c9ccc46ce9a57b807a277498a8c67dd9895eacd9d242d0b5d4e809ee987d8763d482359b2210b20b4afbef76cd191d952d3c362a23aa6ac3e42b147ac221cbfbc24ddee2781aab225295ba541f9fa11435a800cc47111fe985c3b381b4bed1f8224093beb6fda31558da756924bf63073d8f6221f15fb6c39451df98edb41cab165f65c6d02fed321a1c74ffcedbe9d0db34cde5d2e1c643313b204083c27dade064b94fdae429a2cfcdfac8bf3944632cb9608075ec7a4bfef43bab11f9c9c19a58a5fbcce72f25d4c14e79a0ba930bd9d0b629f2128b7fec2a01cfb840578309c276076b0ca264a984659fc40ac1e07ec146959601afe52e5cae5a4208294b4170f3341cc40e3d56cae65f7951ba2028209d84ca7004d54df379e388a53c74cbe2cf4ea1bfda8024517e44ab9198e141573997ec6f2ce9168909c7e67369f6ae885d9fca8100a75a893e921023d5b3fa7ec30065bdb35e482d0b50cdc673b29430585d2810aa4491a32cd03e4cfbbcd52d5b83b5b75b0bfe8386bffe48a8859c6dba4d6ef21a6cc5cd43d2c6baba4e0c13ad9749aa7cb9eaadaacf4a14251aa2b304fc520949ba0597afc596c7d43b75f816915156b66e58a0100daa3ed0cab5e18a1eb0b89d6c6f7b635b01d06008faf994271a766a8e83649b7809f3acfae82997aeccc2db214627a3dc76e1d2ba9045836bf206ee31aaf75140b1961f2934851443bbf3246f9bc79bc2763e1e0df85a08309c10fac84ca02506af1999313e67bc1283ebf7b040f54a58fbc893cc0b3708e557227f28f7e656e6379cc298b32de2a8a9531ff91f3639cc9794b420c1b84eb02b130c47b8a7b34ad6b774959ca53d33b17bcbfd4097d90530805863ceed42f4d4d07c6ac316f0d5457e00a26fbb5828e836fcfbad710e7973d7eb2eda3eef95101b5f8670d6744fb02c56d7e30cacacc0c854ec503e1dcfbfb475b83b2663e9a2a70c804ff178a3acab267164dd4ebac2597a12e43e3523dd15eda4f62588797dc48dd7728606ac2769182c4994d45919ea36c176326b8f283783dfb78e2150af686ef71fabbaa10c4fa4761ad34a09bb1cf4e3a3fd0e68c8401e1c3f4a6ed2ffdd2fccb0cb20e732e0f2afb276cf8cb0b0f9b59906948598049ee6f3b8dd33b49f76bb09ff55f6ed9df38ebe65fc06a92738362c7470d386cd0fbd8380efe79b6e4843945bffb2b66733baf84a28d359a95d5dc7cb3c6b36fc42a90d95a61a41c154fbedbb8ccebda0dba07c99a4e975cca5ac013e1405bb17853dfc6b6cc61092451d81b1b15185c97596bb52868ea7ed25adfc75e855925f79a16a6052683f9f14d13cfcbb77df4d27b1f4d586a39e4425401ab24b682febb34fa1e97895c8995def0d4b20c3b2b7af1e174fe81527bf937937f0227bd5332403cb028b5f961e58e70bb938cd1974b71c67564e7e71d055001a55d4d878321d4c8b5fe733b1f074f2cbf484fe1a1d94906cf7938d2ee80c4124f85379ae4ef2956a2ee80cdd7b3193ebd8561a48ed91ff41661cc721dda3a72b442913a6e2bbfb4780ee97609471a7c07a27aea37a1d4b2319ea8770dc1487d34d7716daefdd5d5b1ffaa74e91749c37bbb6547c87b3383780a2ace4047f50b062606a6097d69b6689e2396dcfc260772b39d57601c1d594be8d0e43c922e981b4c5b8b610727f3977d9c7fc02370421f0a6a8ece72e5cd9ffec8c040cf6788c08a7b7285f7a23ad20330abce3150fa14616f8567a61839bf9b20e1ce11a89db947baaeb27b7aa736efbae890a99fb448575d1111859f8a2c36707d6e4a58a913297c73e159ad61f727790d17820d78c71819cdcec2a94094fe1d05a32878efa463225cc5837f4145c5b3b55ce34d1aeab132c6e8091aed468ee84c664267c5d507ef002cfbc5f32c9dfa691f5ab87c72e6199b7f382f89344d5a82726e11b5d6659d6920586aa7fcb31c7ea09d779725c2570f29cd07684a83e23476f3b005b4e60a56cc7c7dddf894475e5471e79555ac182b7cb19ef834974df601ee81e32364e8778c81ab304d842353cd1c9d2a40cc71b8f080cd4386f89b6078c1632889dfa787e65746ae71eabbd522256d20ffb541a74d2787e9abf39f230f60c8bff620c3034ed5b1c695c7891442b0d224240a26801d0de1794ceede48e6c831f68a1f8fe3b869e55bfdef5f8571564f571681e9161a7bab338c900cd9e61d27c172cf1d91d6e4ee7ca24d0c333110d5dbe9d5102e3f2eb0793e36046065333233585b6b45e944003925fb288f728c35f3c684b6da5ccbae3d8b2b1647c006556177bdb5def49e42be4e8927bf5ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h65c9b832f639cc274c6779d8563e8be1004825a190c495e92525259cbe4cd27bec13570f310b9666a58961e2e520ecf9d2cf4f06a47a953c23461332b11c6ba7b93fcb9c46ce3b8c09a0a4857d7f214a1c14f7f9cb2d35813916feaa65df8a3e1ebaac4371fd6e326987d97b85fce3b209bde731b7baadf5127885757ae0b388601ec033a5c96798c97bcc9bce02b748659b38285a4fe7c84688a4840f1922495938592e356490f00e2e076a418b3a76bc86b71b88a4fef8adf226e3d2fa3bc0c662b81439543f72c91ada785b5492868f97cbfda6a3fae0abf94d242d480b01d8e40a44e4191ef0a18798fb3a008e082b729c3a3bec0e2d75d57bf6c2bce8c7baa458b70a411f8351380a38860096bf380941329cc568d03eedc3d2e1f3590e8808773db07819e9f0d857d5b95f5673c65408ee25d420e48ba38cea860260f33a65ab53f5ccce0390058ba9bc150b161f79914454406591fcba39a210189a65ba521f19d13c78adb219b0eabb810384a3c58ce8fa6f88661b93ec9420f39c76b578d7032ae9260e96a6e82c18c45730375e9b2fe9c891ed3cbc9218d35ae7d883af12c18f4a8ea597e2555468c7c879319e78b3457bf309b1d12dc08d26f7ebda823f9a9988c7a5fb524d3a29e0efb980cb8a52314e06e2651c0a7b251a0fe267f2358304a819df69efd80b9490d147e3e58e227d4bc140b3ffff5a4d60ced8d2b5cc76033970772725ba134e5f90ff0b5a035d2c7803f93a10edccb3dc1b054a43635230b7ae5d44d371cf8f0d498b3a08663ef13b1e42867505c878b68f5ba3f44037b478fd748ca384859b6460e67f36c0b51cc5238e10a0ee986b5bd97f37150c68588f6c6a6f0b2f25edd4f876759d725d6b518b822af5adc49030940241738119b495e4ca066e18a79d7433fd0c9952aff439be5ed214bd758f36eca862342cfda738d5926bb81d72f4948878a0f2da71868e2f83f1d8d39d4060d9ea470297559cc38bbdbf43275988173f0c75b0531e887ecb901fdf2233a746619b99981d93d5ea9dd6c6f7e4a16f2d81780d3fca612ed81e0662a553edfcbeaef2b1afed74d33d50bf79ec9483709dce46d3d1c6fa37bdb410103cca122471094fa804688c40f76e9650c235d42a2489af6f644d4c071888ebfb098cf033a0d03ebcdc81db2365f9afe74568b6e555b7768d9c056f5125490eba4b81ae4a0a55399bd96a3edcb7ae549c789b7c2c25d24dbc6ba5097955cd4eaf42429edc22dbe4749363717dac01556f3ab39494be697eb92c3aef4cef7751bef02031f4ffe6912428aa1ac5b35f13f5afcbe450ebd2c7729203ff16ed58033fbd5517b9f69fbf244144b79054fdef4290708cf0d64b95c2ca8dfe8d5100e9ef429e8ffbacb857eb3fbf32b25dd2850709b182fdf4e5feff172602c2cbe2b19e0776b9d629d5b5c611c0bd2c574e9eedf3f53636751f8f75efcbe113af1b4c5e853c87770c0dcd487543e194842a063910431182adb23828d026cf135f578aa806930e62e1c830371792a45e014c4291cbd152b85466f94639913fc3bef4c1df327e9cf8cfbb964f6722eed8ea998a6278b352aa7412abd66c0eb9c96e2376a9b9806d97e7f9aae1dce4cf532e137cca45c99a6ef6508d41a2caca099ae07e1000aad8aa861b74666dc93d334a287bb1dc0a2980c2d1dac2259f80b7061ceeb804770ad716bf15c5ead6a6129302f936e07499ec619fd77d94f8a9a95cecd24ab8238ec867fedb97e891ad2ed96828308103784f9f57e30452bf2daf68c3cb0a2bbcce9063713b513cf9c4a515ac338544ac376040440da05da3f4b12a1928daf8efdbc15ccb95af75683d942d332ea815971d8cc7334e07d954f99a9d15c926eb1651884a55e2d827e9798638c75b2bbf07cc522f0e181200d07cc8951016d04bd9f431bd44e0358b09f7269c3bebcfabc3e6f00ca73a9224424b337ac6a6cc7dbe5f5ebe1688ee592e532dde8a10065954a5e277a8211a6ac76c96d7484d4fba54a2abe8f31e98b164bfd4d0c7e02201b65e940453a4449a537624ee17fced7ce6c5f2d31e48216ebf7e892b6d3e7c581f59f37de19f0f9a911faebb74362d8b9c618a0ed1455e6c33e62d711209dad72450dadeb10187cc627dd3a0cd416e85e898f496b140ab97be5019135c3fd491cea3b1a5a45445119e19d4a70d7f2586120386a302fa20b0c66dd7509c967d91418f2b959507ea96945e071bb95591d4558d473a59872e3ea4246315ce8324575c2f6efc0ff6ef0131bbc59b489e6a22a010dff9f39108aef8b3e5ae9db7b8e4baf013a50158529e5e56069dc1e548832f05cbc61a5e15680f8796fb5573d9895ddc9480107e36cb69257473f52e79e2ab9b8a5c979f3a1cab2f75cd880ad8c4637373a5fb048a63f9f6f5d2f7647611b2a31056f905c12a96dbb0dad593a267a23adcaf4f0bebbf61ef003799fc6a0f6b7372b6d39a54e089a7927e416affc4fc0b86a4cf84307b0d190e824df4e15eca0611df28401e9260a3483b4b0e9cc3729cbbdbd9cd5336b02d0752469cf8384f599f3f2675fb64551a112bb1976e0a61167a1daa7bb343872396b856265d52cf96eb1dcf68487f43172c296baaab1c5daa03c8e9288d418cfd53f1499f2c6645a978dcc7e664fb9f9ad0ebb76ec8f1ec62287a0a6fac92d58745a5d77ba1b8d94be1692fdf0c9cd294fb911728b6ca52bb5d7f64312977c104860772aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6333c4a78be4283b1d5ba320f6c46f8fba3dc540122c53e52148568a6c621cb3baa884629c0bcaa318a22335b005fe69fb5162753988618cbcd9b3c7c0d1c41e7a5f437453d58be1025b2735af694d84963e9e4ef3fa9b7d55caec777f624c563d13c60a7f804fecab6207b1d14e60ae24cfda26b7ae28d35181297746fd6d5461e1856d44ef90e82a93454a9641f10a38f9cc526d582ee0f28158ee4cacc19aa026a98fd12f36bbec63e5c4eb97e5ed1aace61d66fa0e4094f1c8db51d2b45f8a9e3e2cfca09e9527a1a9b1dd3d72a01e845c7deddfbd7d5ca04de6bb6f1bc5dc7fbb7fdd37505a4b4d343216d015ef9e63075642324e3968516ebd67b9838435102ac4f45de681564653812b734259b68768a23e35541d8859334681ee0327e4a1c2c16aba1d756b8d13c8ba5d015fc0f10377c4603dce6f33e770a8ad55d4e7da2bf36d63c36b4243806568afd79642a7cee81a4ee4cc7ec99014b8a3c552768f00c71d7653cf7d5b0ba987901b3408cc4db47a82929b7ba7d7173e5c2040af00d41734d578eda4ac423213b3b84588405d5586fe44d7ae9eb8239cde5480cf9568a0295804cbf00d32d84919f464eee9749065aac3948bc76decb2f8c30447b1f359c839ce95c3ceec2aeccf3d8129e839c819ee7d39642c68f07f249b5e8052ca9c679c5b836663b6c3888db71b9b0745f44f6892adfd95326db08d62b5fb99a4fba830076dac4b7ec2031dbf561708528b694bc92352ccce0f066812569698d06cc19667fa1f7e31168692ce9015a749b2396f8541d6e177586994bdb944bc7f3a9f2bab63b384146eb913b11be294df957e2f40d8728807f3110f2622dd69105e1b357706f7706bae32471d77f018e5b3d229b3ea6634c667bf641cb6c92743289e364e9104e824e68ed5dedcbfdfee02274dcfe214287197356480a2bf4d55f7d8cb1be16cc7cd6cc6ac0de3b48baca23569b558fbe281a34da2f7ac2e60ee8f5eb12b204c4d73c48b041dfd53f094e1ed63e6ca91ff44cb4092f1c6a56b0cac4b972964a1170fb8b72a01878b9bc97ad38e9a87a8e0b9bfe00dc9776d5f740472fe7d27b2d535722aeb176d61ceecdd6a701fb4f4174ac3d05e0da63057b3dc1266f779fb7ecdf0baca396d94d4693b34e6889695e92b55b4d8f871c3dcdf633c4d4bf9cb189cc00ba325e2f94cd42204bfac799574531c363b191c55e2d126e92786976a4299399e691b3e5bfb42e0035e9bc585c40ee12f524599a3d8df85a31ad1d16c89110d70f20836521bd37c1459d89498c70462ad1ed9d62530ce24f567c4eb7fdc0d6780a75b4d37d045a9e57286d77dfac3c981e39a2cc118157ebd8feaca3a73866b57f48188aa1038f4273faddff8e35927ed39aedb44a8fecb348c5bdafc13350d23137868700624731dd26b831ecc711e03b33b7da596b9f5849d24c87bcd7cea13ff9fd27bdb214254e5e95072a132956f2191c2540afaed7a3f55f4af4d34529122e3c417c5d007f7686702880613cd07bd0fa95d1635bcbcaf212e4fab8764cdeaba02245900b4def0ed22c4726023937f075d9a8fc671ab7651f8ffb5175d0adaded0a7bde0c0863aab5acb2126aa42651d99d63c3f4c35603bbf6fd53576e1233fce8dd44f76589e39c55d0857d4ea9f84e7198a702479b1daa555716deb41435086e6ea4e13356ed503e41a2c560c372342d6b1e61908b1640e6e540b770e835288ec8e53ecdf1de1837a19bbd037fbe73f42887fb08dbbc9ef1431a100d941a15edc78b45ab4bfac34d1411ce8f9f487e1a2b2db6b84fcae47cd774d949130ce13c2c3cf9756a284361ac4916f5dd7135d463963733c660de127f5522beece8fe5e4abf2830a55345a0cdab6c4bf276f4574b0ce058f9b4b94a3a47c444cab6e219f6120ca446a05e380674b2a161f3e5f3c63bd9b5dbb8209f1c2b071a2e183a5bbd85bde1c605fe6bc64e2e1b73c81378ecbb19f460315d28b4a65c3658e568080296338cfcc35c9d5074759c3066d35ca613d072d34ecb6e010e38c61a15a5205f48b8387b470fdbf0408cae4b7b9ee4849f29f3871e91d4ee5eabed8daad78665f7baf5e34deadb266a25d77e8afdb6c0925872d2ee5db2c8d26e286169194414f2f83c3a72e9765a26116150b99260f58f1babc2a938c1f827925ad509be6f4ac9b6af2dcca8d7f74e2c1f3ff4ace2a88688d3f6037004071ec8f283d76c5648057d460224fcc0f42297650d7421acc413c5934bee2e48fc4c49df7e9b70634b8e5ed409c7615ff5aa3e8b1f00a748d6e7bc86fde60286c6338abdc30f1b67070b8a6ddd60fbb399afc2cb7f75b50e9dbd623102057340a762bc185c597d2c16e26d8b1667a5b3655a5bd876b1e33457fd4404980b293e4df477ed86def23d167a1934a730fe27fac54f4ac46e528a76fc4e4f29868b395ea80f309bc6af16b02560c317c5b5f169303724ba92e3317bcd1854968f2bb062aa9023478c7ab8239a523092247b869c7c38bac03626507048566dd806a56bb32a03aadf47987597fa322edd6dbb573c13ae8accad9e08ac5e190a7a0d4bf55c24b9f8a3ed735b4fafb7f9aa105df912be18e2991170510897065f5589fe99fb240923833044aecb7d2272026c5855d4ead7d9b9774d25c6252d58b12054e19c1ec9702ee2840e6c3feb4c39753a6fef6a64f38b984b2cdd103615a52e0412626f73128e4cdc95a57175b37e00d1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h35099b7ad4f07ac72c4db36ab50470e0e07ad4f05d585186174f7441e5759cca686570c3ef76c25ee5c0654ae7efe5676224af8771769408d59ef94bc7bd5e4badb9d4b985762e65c350bbd06b289a68a9f63d2c02242030b1276b2864d04b2d761f24c7c51022ea3f972add54559e108a42be561590dca318b72ec601b8386994d2729551df104f51054f46f75dab564c2cb66bdd4e22b0e2ae638d22c33fbc5a4b2b45ec529f722edda96d23fae9abb5af5c0096f00e94eec2a12ba48d60ba655a98936ecd3044207ca11b92684dfafbfeaf300a18341f44590f41224d1582a2a16bdea3006b8aed7548ba11f02e2a9a7fe6011a3acd09a0577ebe1c7a30bc70544fc61f39214ec84f70a8ac15afc2306a6112b8137c20d8b6a2061b6ebe3ba66b2d675f421bc5c6660e6aeb5954ada2ed34e71325c0a8657bb8b9fa00dca387624b0f9bcf5a01c634c75c2c8b8c546008fad9bd063607189c90feb95bcd4c86710606ae1f19528843a9b00218bbeeaa273d0f3dd0fd623b3afef943502fc2d95d549d192f3fbbdf1df82bc09a01663dd175264c6617b59e699647e70b8e87e12b0460efc00bc10fdcda51ee0e114541c07b1233d54f59553269d9f011a381d7edb84098e774cb396467068fce1229a0b6d02e67445161b2ad92c864b4c9166c1d56848972156807d20c517734fb83d70e7d69c90fde6d79448d14eca161e41ac2594981af2a2df973d2672590664f89d79f6276f4bf861f355a4a0d10f5b2b729a3db5e86bc3798824302676f8105b99b57756d6e2461738fc974f337ed92327c62b24bc8a2f9338f29974707034fcb3b60d40f9dc859f609717c136416cd4064f349c0aabcdc46ff092658ca94fb2295ea46b3a36a10ea388559b6e19df47d95ba77419af43294d2aaddeaea2b865e5ea42279b9379fef7dac367d44f400681f38853a43efaacfd217957a1592e77484f27446e3d61264e3b9dfe858eb3f6dfb3fa71b85f119b88ab6e0582a45225663b91b1c4eaa1592ae3f696f755906bbe7564874b2147f3739b5e92974bdbd415d7c245eea0909a85a54ebf62a5e2b8cc08ab0ebf08951e7ff56fcf04fba5d2d5b1cf404cd0d5a0ce28e4167b98c6eea60d6ca2d055c1d7f8413ecb702ace83cad8346c0c88236901b2fc0ac9a1e112b240d089a5c48f39a0e5e091eeb751b4f7007f29dc47d2b997836069923367b9f90d01ccf8b93ca0c5e432fb4bbaf47e76e65a8647a4645f4c6dc92ccaebb96b469691d073a51af5ed558b2a19a617214ce24c759c57065316dbe295bc09dfaf401fadda21fc065193d507f52346c1d8efec1611df69389139162172a5a8200f4a76e1543c4a535b03d3f92039bf8fa2e9cecba482b7bfe9bf2572d8e72c01e0710bacdab777ac94f3b21a01d9b2b9fcf0384a918d644e38c8afb9ad4afc11e011216db599e0182f64c1fa9856fc2e8185cc006ebcbbf9b6b9657095e66c7709e90eec6d53e904d3a0cafa4e31e125b19311d6c2711dbfc77e07b7a8f6237fd6b186eeef99039a59c9bb387951a4bf8cf3b10f0c45a56ac8b666cdf52b415ac99e38b9a4cffd022e37e80744e5f46c1e2d32f32de7c995b2f62faa530599f5fa29d7cfd832a694bdcf350060ffddf88678a3e925f114528640216a13b53445bbe3ea3f57c8ef0962963a9db8515e23b990cb0a3961699bc4348adac26f289d14f0281c3e8c190b78976bbfe98f1ee0d7a8b89bf6e0a318e161be0ebb4bfb532ce4f23dc4adf22ef1cee270eb7f90d1d40753b833a5429e297364169d279692c3c21a616e4856cffde43758e74f5444323c5741127cfeb574ecd1308d2a98adf101d1fae314bde14b65552fa6eab791cd19faec2db2a36d75ac14b0c9ec459eba9e6bfdd86868b7bf0802c2fee344ccf0a9d6769c7fffde4e9714f99a0ec05c8f85a5d1ddd656e65a65cf56d51d5e0f7b75dc1d4b238b46737ef9a2a39cb614b98c0d923cc0b1a19a5c463712a8bae25c77ee2e4caff11043217b4213d70253069f17462d310d5ec7e12aa984d0e906e864a2c4654194eaabf3cafad70525c1fecc6998d36739d54d1701442c0604f954c6f228bd463a8344d99765bad86f42cd11f8f93dfd9e9b9465cc5034b87315960e443353d778045663dac4c52a235c3ab16034cba4e41c6bd938541e189b7d3f05a2a66651d2735d4a6b1fe280c1f6be8b86bf3b3fce5bec119afb925528f4ce04362bb758809f24ccc7fc5ffaf2050b454109db98209ace4370d04cb76b0442c5ddca6bfb36428b97c22397ce976525872ca1e48a764fe000fae5f0867528b8de231974630068ff78bcaedf74812bb3af9e80b496552cb30d630c9eee936047977908c36fd6f9e2e5a173a41037f3f7d194cc16e53b094061cc0081f873f2ec7891b4eee6f1480e99d650afbc6a0dc15c67400c6793648942bf9d105420a59e0ef306549c2d9f38b3335eac71b8235b304b22dc0d3efd9d1ab4e254b4c057d264e3f12ed773cad14192d17d12e8521eb4fbf5c02d15c1bc38aeba5733e9ac7b5fc522308d740f6841ec58e61fc943daf03215cb8203a76b45376bff5abdef8560f6ea1aab3349602b2641b09d288ff7a4973bffca6faf1cb9ecb21251f11301ddde1fbaece2bc7f7bb6cf39212fd389ca0092a4563947ff1cbdd8bb912203228b125fbbdd6e670056f597b88fa237ed353d4d65e07f4b724d46a58b380f7e17887f4e14f2acb79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc8f1e2bae817f641836e8bb08b3b1c54aafc84db05185490dec9dc708375e8e696885222add8d249c8a8d9afd6028ab13aa119dcea835a7b6f7ae16f9e35bbdd68a0fd5d1034e1dc68633d84fdb01d5e5b1ed48e2be6d8a139a28c2a09685182fc84350ae10ef73f38d075f3c302760fb7e211fd2ab16ce3c202662b818376c1de22f6a45f904d1d33e692732b2467fa8dc76a6e7b4cd2e58498cca3c65f2fdcf51b5bf1e4997398d89367a43eb82db31f7ae177b923e0c4e57d62c0fdf084d35127473cc9b1782c2e4e4f708a41c56ac27655323a9b313db168aa14c3c1f8369aa9ab2ca24c072474c495c78ccff3fab0468e3a715403addb4b9520c4b347495549171281b23535df7032a662e19ddd32ffd657e799553561f10f975cf5c1ed02d5d494facebcf93d8c92c1a0df2ca778d5ac87768a2312a72d7d30a20e4f6ff109c5396b2f8d530fe62ea34e1c26f619f9a89bb06b65bfa42f555d13389aadc107ed9778caf2d3b1b218c47e27aaa992be35a282292319be2ae3429706937a65e9d876cad38dceefb3eca020d76d5dff8cba4edebc27421bef38c373d7313f0df8eefb347ff046830c282b954c2e605523b96ad8da215844b7c7fe2b64c38a38631e0d707319eabf4c031de0ed358f104f7031ec48e8eaed3bde4fe19ae45ac2d5d0e0edde8b3f2936459cacfefead2661234d516559830567b64b71a6b8f5cd2f944b2f6d0927e3d2233bd86b57e4dcd173c96465ed8e72ada941cd7350e7a5050a00196427a4246729009c31c3a9a18b288a81c49ec461ef730c4b91a81ea4a7157dfc95f0181f43c93c47591aac04bbbad9dbdd54d98ae4d44a9934c3bd5e6cf5c749f6a0ab71d7fa5e46d8bc145d2dc03e7e1453700d99abe6ae7ad291ed15c3022e5ccce66f50f67d24ce3c2fd3cc09eb44d6b64fb31e82e4af1b75fa6e72d970508238cd83dc2043985a26f0e93a02db39dfabb5c72e616b6888ddcc6eac2bfd259828e2fe11ae328b6150120048e9aa0c853c426f294016c6f856bdd744c2643ced111e8146ba3c94f3cc66fbba49979a054132fe1ed2ea8651d93b634eaf4a28624b2885dbdffd1d1050d8c6e4412380703483c8f5e10e21c28699df061627ab5a8f1b06d3cf5e0026783f80d9923827cae4b3ebcec3c1ffacabe2c0446f1d2d9c8acfcfda38a05d1029331822545334bd2e185b7db3ce88ac1e1402f9ea668883c001f65688b9c3fc1970226f45445e1fbd4cb42a97274f25625f55395fcb43003e29a51d78efd65b06587983e26fb1f7fd078dcc314f09f774500a690451c0d374fdb894ae38b8229297154c84a9f2ea188599e7e4c648e0a8c1ce02db04da1957c838154b16d53922daabbeb4c508baadbea4c28f6fc90419b94104882c01665d79bbae615c6d2a8768117eac095c3b737dfd65e941cfdfce219fd45c4b652b091c27908be4cb4a977695d216d9c297845fa2d34e7fc1a27b9deffd7c9c4eb7e2d295533bcb3cdd3ae575c805795d043a20a53d6ac6fd810f4849e7cbf694d803c8eaa1e1e35662f6f5183e3c267ea1ae983be3caf2da010c9f9008180075f2b90c946c944d4f4c7fdc0022ea6013668e279496f2028413607e10b770e81b134a833de00694670f792aef25d03e25a92b565ac89b4325922cfae143d9c8520ff70b1cfa73fc6a6f9d1a77f3b1847d699e3d0b8d622a70b3784075361a504e028e1ed2d422c92352231a454a5ede75c2c97f236e11975c177e505607d2009b0bb7cc9c7f252b9d7a794bdf481e0a840406a3a1ea2999bf64532e5f497702096fde630a84b11f70f46b9fdf16444e32317cd881e35d582c36ca4f1fd26063525385155db28e2445361856b684fb1a6937de2bb0a90b5e40df7f92db60e84cc7655eeb109ddc35d5d918a71aca7b071f18abbf061953476ce119a7ffcef8e06ff8bea3e8f7e41253b9fa347eb0fd5636c38ab5ef028602af634645dd38c0605f0fff27fc923ec5c3827e986e1a0b7b6d3aec9b305b5da60bdc56d3a4d138bf5135b2669a5b667fcf9122b1dd8c453e3caaed231c5bf96c2dd3d783dc05d6e9608755d53d4c0020311b4b2afe47746261368234b5340c551723547cc86fe31e3ef0fcb1f828621e517e48ae914e274c88edee4433d6a7e5cc6cabd6e22a3140b2a51ef067284442c773466f441b39a429b6a38c9a31afafbac5b590c063e53e26d5a4a967db3ebcb19c5203e9a1c20627ad0d4e2f9316130d5540473ac66a3c43151eda316022f8915aade7acec53daabf38610ea6215aa3192c0daa4f27824958cb0a46435691e99a4959ad85d2214972dce6041de081204ed257b146bbafbe5838dd96a3a005ba6fd8efb82a94c70852dccfe1a3f1881463f704ed2e7d021ed25feed2ffeaebb2a6c08afbfcfebd3435522b10464120e9969827a3b44f41417d0c22d09b4dc5d53a91aa3a031483a3b2d8229eabade18f7716c0f493cb0055599fa96045033be1d682382065813faa4a6b9058878d812253441cfaf13895b31ba4311c39e4d472b9ef2edd5b02311b3b962c86ef2d5eded8661cd79d00bd85b3a5c43b4165bed309776b0d47289b1b5f66da6a621eb91d8c74b036870b9b57eb1d784e1889c7dd01a746883014a208c36295472d123b538dffc9b21af2477a69405db791a888297ba3c4ec259fa15eadc89521077c6ee8b4048f7146c379848fb938d75d9b21400bd063f6c68cae5c5ccf405;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h14379827898c77f3dcdd43b44598cd4c97d54ca39e08cbfdc4861ed91f1203873a183f72402691c507de5c43cbdcc6211473d5a2efab173e01bf2844f02d7fa0f0e625a46aaf1f309f04232a871bb7f3f687e482e08492dd3b1542a61de75b708d16e5bcf7d6c4efc790dabc28c089f95d87d80cdfe18442cf0fe8c4d749404a03b569fa96b01fab6c337100550b81a881f7e2e46e86f1eb396d2c5b5046daf45c4dda1bc4aec610f3ef8fe9d68f0cda8eb91ad5d1cb7db2c4b7923bb38fcc938f83595a632c2664efe0174a0407668ba097cfcb12d7be55480719b372f4a60b3214c273b38c1df4692744631ba1bd6678bba48cfbd70e7ac2a38d2506a0dedc1bca353a7659350cf290399a24d21f2762bd770b8ca6d5bda83634c72992eebda6a8ee03a11f0ef63f7febbb704be5fb28a1c9f1721892986063eba4a324715c59959f8397e3bfeb2656c41ca8dc47d5b4713d08886883d6882f33b98e65fb05265b19d788ce96ff5e655669bc58c9a65d8d1c3ba10788c84c992cc6f30ddb5ada136b4e30bd3e149bca62489b9abd5f04ae4a2ab5f8049452dd78ef84a1d57983ab9acf9e229ffe2292a882235f847f8e9365be62d9df8bdb8cb04aac1ab92a73d06abe235e72bd0660fca9ab7ebcade23085cc667e20028c5409a5c01e9d4258788a638ca183235826519afc55a6963c58f8f54db04ae841a050224dfcc19dd7d9c282bc40a94230d6e589f5c146176935d20d7a75c9c11aa4d55df6c08d9bbf8cb529987a4147beaef5c88469ffd6dddd7672f3624ffeaac70e913ebbdc2a7dda620531979b1dee3be8a3da52d5982dc3a75047da7d7c5a3accf03668652dda1deb33c993adb8c2a471a2d386eec785e23f417f4cf24dcdcea852d2f53fe039b5348dcbef560e08ebbb7d5b85542879f67e944043736474a9ac742c3d1039b962eb5807a15472673bb2c9a24d8c611013b7c54982917483e5d668d54df37eeea3eebc56e3bfe7dc54ced9f149123c1f594532eb8e5e29a40bf32e989ef3c4bb468a864f34e2c7723a39929400e32bfc6243dfbb1332921f3bc57fa931614e1756291c14bb00b2828c99a31ba73a34dfd72f03ba071e29bb5a042fa6b727a8234252c1cdb305a01cce4a6455e15bfc78ce4de4c31e359e94ed56f1740c825ec3db95fc22ba977cbcdd42019c45150ee3ae25d8ef3afc9e91f24de71f9e7f480f6869c4144a961783e3e6ff5e69398904957ca4d7938ccfb009119f46bb4238167849d4dfb185bf14c6719b993a8fcddf84fa86507ad4d10191275ca4372d66d4ed8b5e2c2939c0e88cdf9d16536a034f4318c2e86b6c91123e2964d97eb39374835c2aed06a19aa72cb1d1217aa0a44f897a92e907e57f77ba60c31fab9d7aa9266ec622cbb09158ae822c2dff00658fdcc515ca2ae7467ebd16a14f6f863a37f164325a7ab2482ecc097caf051aa092c5c4c92ae84dec51dfb96e145a0bcc51b15c47e7c5cee8f3dc3d2c6c5edbb4d6c46601402dd30b0057b0894e04e76f33d3a24599045db9babb9d9fa1a3b10195de68c34c679e94e888fd85925951cd32a9495302a304ec6d87544017a801d9bdbea7a97310bd6b8a9b02afc7ad97844015fa4cc1bd08bb1ccb87727d2790bbfae2c0cdd5a43aebc489c3e3452f7321867604a0b527039aaceb70eee59990493d56d479e1558c1a5d94cc7707eb0a877d84b86d34e1484caa2d40c17670805ff795abef9f432c86e24900779cb1c4170e32b2acd88953c63a05de1f31636d5205fb6fcf945c717a72841276bba7fa76a99feb9a64e5f78e3f777a122ed81090b3fb79a8bf2adb77a1d33d0b605c6f6b975833e3b0647997e6df8cda6d21f42f8077794c734baff481699771e239ec485f1ae3331e18e7c0b9aed5bbde6134a443770c27c7df739420960d8ffe68c371e0385a23c84d22e66fa1e88f966a3cf1f4f1009ccbce3460b1618e09a58f5b5f40b87a1e3bae384dba055190c96f1e5e9769f3bebe904c9748d3873afd140e89f6e584152e0239f08100007faca41ce4d56b7cfc319c4b610cf9d5041a5072c5621eff398c5930fa1fec6cb0060bb739e155345ca9f721328828038845ff05223d29ce765f0f1aa789b5b6e715f773eb9dd92f49c8f8db8ae4b94b3c2cb06867a29559258ba4a370815e890cb690838836f72dc5567ea63933a518e9d6a19f7d868efba4f75f2cadc7f581fddffb4179547f6bca2acb62c2ed882ebe3a8a2eecb082e4f36bd1b1c3c9c935b564306f98fa871df93b79ae4186ecd0d66e54ecd4ec6bf1c8a6897ef6155bf30e00c6200e0a3d1199f3baf8e4151a903cf9113b86f2168df9365839b702d27b97dcd5b8bea1857034f8604ef59aea7a2ac2c14fdb516ddf40c503d5037a63ee0f6162dd4ac657fc40f8614e8f9a2baaa60c1c234acea45c8c1bd9cc1c7b86d07a5dd8b535e0738020f3d2425cb5d7dc87a325ad4ec0e255aa55a95290769896871e8d5faaff4661a6030a9e751da9c70cae3d4330439387655c80ee653ad3ab79ddef667d87c4bd3ebec4366628708b3c9dd833366f185f044f4ad7576d09ec922678ea46f4c5d401f2e37736f747a8f0489ee00c534e332422a871cdcadda7e83115c48dd957b44876b87bf7517b8e9c37fb00c11c81d6a850f77898b09eeb91e6c909584512d1420b18d8050a252bc3702b463996ec298ed0df91685ca0f2500da61cfdb23f1bd7107e10bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2edbdd4aa307e2572fb6c1ffb840bc6f9f6673ef7f1566dd3185606f154389766f0d16670051b7e0196d8781ba8b1dac9121e6323559e423e1d107cbc4ef15fb827e87900783113f517e48444277cebc73e342437023ecabf37b6e232be0569f82674262eeb952f52e99d3cf3b9e2c67dc5078de6f6756ca74dc30060abc55e7a11da79349c21234311592f39c13ead259d5d4afcb1f7108e7188b01a13e4409c5447df26c6c84fc9f66bd80e6ed16ecc5354500caf0099b8d3cd1595a60516e2cd212c4f57fe46d41a0596db9abaac10be9a91c3f8a281acb95e9a3674f1ae18cedb1b00ac6d3ff3bbf842053f6b718cf6d67a55eceb0f481cbf29c3b4656ad1236e9115f6a0efd055e0f25e5634cdd68efc046f2224267fa934796cd6b51f4840fa58dc581069eb43f4ed8cbfa88ba755f1f61b0d5e5958eb25c3246a6702622044337ae48b738ce14886b1b09fedb4160d9034edd5005708ac07b55f6908822b90d3eb869310d2024e69bc686da1a27b430a72b3c548ddb06e340ee88b2a2242e133b065dbe5a1c8dbf04c5546f034855ea709328856acd303aff50baf01b38bfc5acd6c9c581fb76ebd4873636489b3d862829dc9a5818e46b97d3ddea98752fb33dfedfe06f293b0d5dfa82a0213a1a322218c28cbb6783b7365e3618fa90d883bb420950eda16907f81a864e77da0096e481c9856841b1e362fb6696408ca274c13ab4cce7911fd33fce9dbcc9e2f776317942b728c96164acfb6fad3a79bd0159ab279d83f7fa620675a0265db62ff50a225cfbded4020b08770748113c2ec4d9dd86a7bb72ec9d0ceef68f6d26afaded5567ef57d272ffabd1c08ee0bcb80d8d01f56be420296771e12587ee0bc1f09fd994bb10f5209fc9a3b9528ade192429ae2ecb7fccd5609ea0b04c53aa9efc0bbc58589ea200c1df58f22278c992fd6eb6c4ca46168e7e0786fce4e504a00e8aae6dbfef12d25a75708f68bf45f505dd21459092b0d02d327f1ff373916f112d6a5d0e456c2126a275c114b8ee18f649d3ba6d4513f1884eec469929402912d0030c28e78138f91ac23b82cb5260073dfc331b7a93eeb30be6ec7c709e58f41dd3596121313f2b466b00010341b84d342ec8740e212d24b08a02f47ba756da607a8515f65936741160e26168f38e6ce90b95cdbd592b4e355c23a7150d882aa2c32f5185efc710038eaf2984a1a97bbf68fbb67ffaf434de3c6287b8040b58f367e7a759e64df27e17379bf8a08028973ac242cb38052f6c479f194c78122a5774638815f2429c170118485dc0ef9c8e36c1542f01f654e83447f3b4262805b3bb5836f25a75b968451d32320cd5d283160b655f805d9d6752658e3982eade8da927a690388dcda2dcef88d4f7ce6d3d1f55dcbda4c1af2f0c6d36ee236dc6b99f0d7d012436b9c2911efc55cdd62153a7c69632c65c33fbc8f1c17ecb70c2d9f7fda772bb3d4c8db14eb48fad5f2036c009a6d709c34b5dbb0f9ac21dffc2fee48ba98668945e0dbd6c9c30517d55b06fad3c0b6393fc0a89b5452d6bde039c48a563cfc652dcffd748e406d29c7d7e5b0a1c0ad29e731d6c7eebd45d34ee7a0482577e3dc0caed37da52aeec8a0db1717a1d7d07cc7da3b9b883e1e01dd3d886270dd9f1a57956f8b7b2758ae8a6001bfe2997de78bbd6cd2b43032db10a09f7a12f81ec830d9365cb7edd02c5b39aaec694f1ac988742dcb67464478ac16cdf19a017d45ca50a6f922e237d6619bcfbc84ed8a707fc18345a62dbebdbefe8489491eb5a8ae9937d27913fbc043fa70749ad9a8bccd03a098f2be099e8937455428c13c83a8ce60e28ab7d668c14ceab989497325bd6c781a2ebb9cbe04c871d0e8e02087c4eda7feee00fb76a08980d01138217e20f11330fdac6fe5f39ca1a21a937c99c3c34107fc7ad787dbe650fa129d13433bde3801bc5699c0f99d7d8e7c7789ad535f4e693ce94fa23adb2fd55340d3fab0d37650b43f4865c5f152047692a589704c026915aa00ba8f398420e92996627a1837f42f16b51633cdb009e56c9b398989ddb56076259569d7f95d0fa4a918b17625a21f69d000ea2fb367071239f0aea1d6668e3e979f77508d6576e7a02c301c7aeb59f422fec36c6850998a5c57f39660fda82a27391a586906f949287c100cd247f2756c0887ed6b807e7934bc8e3f01b1c590d91676da4e03d955b67a1f6d9e7a39e8279655695dbb98386815d47129e0d5071a8827cec722ad169aab8df79fee5a2160e66b0eccd523a32c07d88664555d5ad28ac2994f78d3e63a5af985b4bb3c4cf71e46c6c2ea021f8ae334881db599225630a01093274223468731722a9f01c7f5907064ece859b3bb9d48c85fcf976ae0e6dc3ca8d76f10217a1f485f0bf92d5b91e0bc5c4bf435e80a0ebaeaaf1e242987c325fdbffe567f605af89cba2f318325184f68bcce929eb2a991790dab4676a6317d147086cb32b844128fc74a9d4e3e72d1daa391c6a37d5a5ebf5a9d322fe5f403f77b9b2ed357c99926fe492b2629347580cab6b2a002a22c264002cf58d1516762bb1472393d98a639530b890a71dff3e63cf0ea1d8d8f145945f59fec0297ace154cfa238334355cd64cbdcc8fb82c89018fc5da238f3efbe02d8f5fb7ebe812b886b53f0415bc24b89ea67222b65b0d58aec279f3a43ce175eb844191ec7b84891f728afd9db14cf790a3fc788576a2e28cee5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'had925db399af55448acb58c98a5bf136ca29b9d27d85807670114b3b649f331d8d1a4ba0db32c29d6fb7a77010b07119c05c269f1fc5a500e591b7863d9866d4776216afe55412989a42253b1d08651fbf9b7aed6763fb9c03c6c4200f661592a71c6684f248e1ef2c8349f8e5255f834504f2f7adc63a39a7ea8324b48efb9cddc136ec3f043ba76cd323910b4fe355e1890996f74b08ad0c683f41227a7f8bf742e552e9d37a7a00989c27a20a3f5b1968f426b99f6621c65997344294cd59068bf95bffce0395b61b4507886c9e59452a539b299cc4486105a364cfb578e5de65e757e240663863c2c0b0a0cabe53efbc23201b12f2e72ff0203fdf9a3a119dbef5dc112cf5ec96cf95e342fe61dc7b2969e6abe6218bd395008eaabf3709290d676129a82cc55fae4726076d10bb18fffe1657e22181e1e95e2bb6afe61c115f708ed53a4c50408d9abcbd6066e1a648426048c1e76a392a780156152811f4ba5496f7be54e5f4c8ee7ad35055444a75a640febe53e156e0c5d1e1b1011ce97fead81a46a509f9ca29ff1b438964ec679d72b708c817dcdb571930bf251d21351ebfb3bb5b0a190b6b1dbb5d4303eaaf8e4453d06523300484888e82a4830df1369a2dca10a7512c44d98ee3773f932d2c2884bcd81eb947c76a0a6dd391113e756b31a62fa4392b4986a85313567985d574e0172187b4e1f78ed07c9d5347c56ab09d39b6f5cd5b10ca0235b7d2dd3753c9290d77f80e18b2be87031c99ff6ea37cafe99f75ab9da4f6049cc98fcc39a93f54871323b9c089b2f08c9c8e518845473470729715adb082a32643e4d8c6e444d6dcc1e3fa5270a7dbcdd22a249a6efab4cc4ea409d2a7ff1b21b9a2a36cabc1715a7b91d901444b03d18d8042837d1779a200cb840531077300f12e5ac96e507c54e2604c6f51d1b119b9ebc74df8c4a79f7c8c368c0ea8a7dc6c9478b8b24f010c0a6cb896e24d5dfe749ac526ff54acb12e295a9bff3a50ed1ea6428da8abe6cc55ce0f798fcd421924fd4c06474f5ec9c4703930eb7a5cd8462b4374b3185259467e6521ab92295fc11ae3a43e2582b0fcf50a3c8b904275ccdaf56b98a0a8ddd6f8a5dc9e609c6d87a008b46ff0d9267e5fc91e8d13ce492aebd0df88408fb1143ee2ded7566387e288c52e5a1f77b0807be7dc864ae1d58997bfbf525efbd53c7da4ac224cb2a5a10bb593daea8dcf48eadfe7f2d8ed1864ba40fec048e2f3d7f4fd18cab3468801cd1d9f44df478b29bdb489b5541bac88f51272c2e80beb4179cf64d662c58ee308bacd40ebe081c8f8e70b063bf0781500399a1559295e2c72730ca88b259cdb08b0c2c97f69bc41dd248db528777e38f6a33e0ad4f5e4e6ccfaf58060e04db910d5670803b2d45cbb4b63b1c4b66009c675d20e19ac16739ae8dfc8de653d4245b54b1fc923971d2314681032ef049d140d83981fa181a4a6e8e3b190d668f69b4c4cd015b81a4a6fc3aff1df1dd5381d7e4f7f1f0523c1b930c34c9b879f97194250799aabd77a7c3d45bb630624120eb2b83a423f2a0372b9a54346d22b92e4d618f1b0ce36c21aeb35d15b3f9f4ba625f68e50a0830f15bf4b61fe3df1140a51bee999c924d4b175c459edd9992c348dcd0568759505eabd51a7778c6bdeb1d2fef8ee844956ec5fc7535af969e0950faea437196f131b009c85504923732f236f403f65a5e5a65bdf97d0e44577d8386fe964a615bdcd1ef41c640eb88b05c17ae3588610898f4082d7f52ed2c4d2a5506cbc9ce15381a24062d113a9791251212ddcf42acbf4aedad47bcfe9d0ed8886e30d3c9d447cabdbbb2a57ab79620af3ab35be2abcc45a23fa59889d562ffab2b0e0c6563ed4be38375690b0bc45b9b7b49c0ac4955b31d07dadf1fee475d65afb77b1ea41d8d480263cb7cfc15a3157191dd0ff1f3e0a073b9b11b5e3c23a8a4ea18585136f356026266268f79275b1ddcba530fddacc0d124e37b1e39791ab206ecb44ac936e944dc0851a0bc2fd1b3aa746f84840ef94545e7e210dff482d14ac880380c802f1a723e63e8266e8ebd3930d73d01f0f695efc2ff2a126b373dd45e316e26f4d851513172f8784886edf23930d58b5995f8931657eb6dca7adbc7438b3d72f1858eab9063c433d9a0f2eafc4c1abc4a29df5b759c750252017437be59ceb12b0b795cf2c39fd28dc99f46af80b39f57059ca04254b6bd275bd9d6c13374f39e2ad4b6c6e95259cbe56ff68ddb694603988c2d2232e0213c0093f0d4022c554ff1435a4e27065f2447e3e0150df3f54cec8a4456a31831ced8b5fe45e341c7f865f833aaee01dce6c9a8dfe5250f5c0dce795628ba6631d2581433e15448d317269b4002071e7ff2226af0f7e71142da1e8810a61589de08a8b2d7c97569180f10fe79a25870068e341965fe3d043039d66bcbd57e9cdb236da3df64a0a09ecccef8e274b1d9415ee858e47af86d18d9dcffbe2ed2e44c6d9f30ff39b2c37a865c0be91384b1a4b0e8e77a2b1d7db15d31756c8c77c94fac2d786ee033a2249db7a760e2ce6002481aa9f8292b53074bba65d791797557cae7cba15702fd9562e434d95761ddbb47559d1f5c310e77bd671b6d050c43a14a6eba96eeffa6ef5cb0411e10d6816da3353fc03fdf26573ba95c18c40867c10fc342a45d623ee9b6b6a26e29cf01a1893cc431a40345d06e80809f88b48317ed26e07f63c006168;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha7af0907e9e7759bd6d40962ac87ebb0a8f66ce9a113495ab2d57a78c62d3ec95e9f233f5f8e8868169184de4c60cf38f49f35152ade9f34e2a5104d4140ba7bcfe18300707da820f7a1360f82ab28692bf4ac3a5a74333c6afafb0b9341ddaa40a1ba11bdecd5c65b0a91e8676aaf5f6c5783f89cbf2798aa2c3259e9c4df9bff64ee7d577fb48dce73695412531bc75f92eb13e2bdb96e938d5a25d4b17b83b53f9c5b317c8ce864a1540af4d317452243e4d6e8f756e7802d18998b2af3f58269ae63a4b1beb6cfbb8c899e555f19d6f0bbbaf23d4445ff1ba6d5e0f445eac591eabf66110ca2cd8ff65c5c6bf927273366984c852203029765792d337d2bc50ecdc2a9bf949dd311f515b338515c9914c8bd1c14dd4c5e8f42d5b51306ab87e40a9ab884b2743135e3c51deea581b2e0f2d670310f895f7dd1f97b1b1c04836d7bbf2c24495c44d8d63d060e81db6cc78c43f2583f4232df6db044e5319bfbc69f3a1d58311ae3435f7a99a4da328cc98f4ddaa3b73184ecba03c8d7a1906aae9f1aac0805b81f3797b50af72049708ddd3d069b10b5c98b39e4c0a4b18a81d051e7ed60027340ff7506bd4d177d18c8078bb1dac8be48facd372a9692ee32ee77af5d1c5023a18913b04170caa3f8a511949d895ceedc522659773caa6339f1e53bde4bc949b2a2c24d5da6c51084c25553bf7ef7b7a49cfe85b98976de40d60f79122960138674f362f7a859a921dea989f9b443961ab832b096e994a82792f5195ed927394172f474f534cb060a21278d74121395f53e2e7184b8c6c7ab50da0b2b0a71b1b637448805787857f8aeea748ea2ba2464a1c32395654caa8053b86b53df01bd507dce6e63292a44f2f0a5731d6a21a02a222098e22846f76120147007c96b67b3bd57150d36c4f5d5ccac56766b2c793f68fbaa6a0c5744cb6368aad14d3b6bcb0d53c7f1cefbc413330407a4afa677705713db6ade6ff332df5799bfa54a170ca9ba79c5bb906e19177475e8ea663fb1440551453dbd1517775fac872e24e6842ce406211ec2c0f3a86f1a4bae67f7bf69824b91b392112f1af931872a621ec8dd1d75df29da242d307fc3f18bd79098b744a28f43c6ca64038b0a6ff959854d9b23827f873e862559472b91d45eeb1be147f0f8b6199782ecfcb29deab6f227ba3de66003a9d4fcb6b286572e9b996cdc93d530ec530cef5595ebeb3fa9cb5a1a0b8422c5174946e99dba1272d9090fe0210d5f31490a6ff14aa8898cbe9f7f5315118526300f8fc6a613106c32a914c0f72c0e78274e0339f6609b55ba8cbfcc2ca08e34c9592f6d36be511a8948fc63b61f914fbdc7d199b17fafeda35ec269957db8af06c7c3e7a5008711b1ea07628c3692472d51f922e9f1f3f7a5764626a0850b52e3e9a85c47d0fae755e6643b32b204b2c2097951ef4952c3e0dfafda860c1fa1fcd22f0134f16e6d78fffa7678506389854ce3ba1e2c3da099170e543aa8b4482573f817105f720dfc9a8dcb1286dc79754e19213207058e73348753032c497ca5b35a8d748eecf5da01a105e857d7e33173026196e048fe8c367385c7dad90a938976d84bcb03a3f6216907278bf3eb9dec5c0e929a95b36fa408e7ab704e93e447f26289693d0d1314c8360c2c982d352902b560de561400979c6856cc32a405b5eb49d5125f6c2a93d2b20c24ef433f2011ca1a79fd198c0993ed0e36fde89d2f86d017793767ec7ce8cbbcdfeef1892b15a768d1df1291cba4e30ab3a98042c9f39d3ed7ef6595b0defff23685415b9184a102fced099ff98a997c2b59ccd12e334c95306b890049b1ccca642e0d36e4b26ae04ec998845c38fe6139fe4978f740cb54b110d9a5b30c7a72835a4b20348e8c431480bf0a53652c4e110d99279132128db109e804f9387cc897d8901cb6516a1f085de32a56caca7859bba3b0272c9df60d585ea18512c25ee1b6c158f50c2b8e81ef5d641098b026a79005471a96288d1650d9e4f311abed4b06726f72afb3bb618d228ee0985fc3cda935f533efa0d6434bc73411150bcf346af2c40795bcfaed73a760e44c2ce5f5d44d73db9888088b080963d0762d97feb29831a2a6f781d7ab104328c994e3ab0ac635904da28b03d204a643580a7437ea86d31ee3e3a7cd1f0f42bad5e719250df1003d88a5e6575bc32eb32fd2e594cbb4f1fdc49a3c7dee3a58b02cb3a0171e67db016740d37de677564ce302bde7fe99055ba418ea3c72d6810ec3ea1860d4678992134ddd8ffd0024cfd6554d3149abc24263364b1d7e9bd8b2b603bce0bfcf539613ccc050b0c4e81d91b7b79e6b10dc86f406d19dbe8dcaf2a2dba2bb42f663d4752cb169a5660a90cb83fc59a96882f1c92b574d3d3a1c2f5a06f30299d9c4d9b789c4a2bfdb77d959f0d365887f1355915793204767c9195f6197b77d9e9d60a0c4d0bfc8bdd8d81f861d5d3eec027e83d9cf963eef43fdb552ad16d74ee8299b8137a5299782fe5eb006f8be899b4feeeb71fe220cf8a9d1295f6c43bf3dd11b74ae442ab8ce4e0dd3f8db6a9dcfea2544c06eefe7aae03f6a5751199a321f587adab866007e599859e1833da03bef8703585f70008bf47ddee2e74619550c3b46a1f77be8a5457e2207441e4253f5a19c24ee460f8730512cb82ab808164440fddc0f30870b11debeb6462d212f0addeffabfcdce73652973f7eb39da843c2217bc87ea655dee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h72001987305ea2ad45e19b871db0773d9511c1bc3b6e124e85fad16b1ba997d6e8781b7d9b23ee2ab22b11a95e524094f93bd24896e40da97df41e64c39ff195ecc05cb69067141bfa333ed763c04d7b93b9ad00fb173a779619e8b84704192b35406aabcfc19a847ce83bd39197c26dfd6f4d5f7606fd9a00aaa128f1a2110313283465b5e25501d396a8a1937951473255f9158d2b9f566a9769701da54bee273448cfb82f9777246763e560fd1fbd5ad28d04c61019d1e6523a5f38a563d323ffa6c22ca9a9d80f3fd0323885aa11c5589a4c1d00bc765ab8097bea526b1d519268309fb65ad004e9c27a4b62d01f6fd3f106f4ef55077f97f1767df519e486b27a634c85ec9965fccea3f5d7857d8fd00b3d2a4086cf7baf8c704126de8d6dc0d47c2da50af38187766c14d01c51f62f5e556cdfc77e4b12342a077ad34dbd3975e4e328b09b0cd2eb00a8d099f5b2f6761489bcce7b5b39a1eacb2d330d9c6dfa4b95521459ed90bf39cdb2b2f86bcd61dfb2cc13f6b26167a3c2543c7e14970fa5bfc50e5191172f926bb697b1c93d7918deb3c17442d29fbbd3f1d823d7234d28431dfc455dbf64de25ae02ca672eada120ed4469f9a07e4de0f486b35cb3efaf6f1142b5cd1e879554a7e2f567a8e4cfbb6ea66626ef9e6a534add7133615ae33e61226c5cac8f2d97354329e830ae7de22ef073048bb3cacbdc28a9eb9abbb7261491775922d9df9964154400010c343a157a3094269064f92b7790e07a9f7fc2fd70aab92d3344150999f144c96fa573332d679f4592b282e3d9b42a160571fc811b9fce46044e161575f15ff9873aeb47772d095e3d95c8c4ce9e29b9bf5592233ad57421a5ab8cf125e93ae8bb30bccbfe43a3fdbe8f4080d9685bff8427af73d721bdcd25363e35d7b12ecb849c5ac436a86f94faa3e3d463477d9ae3899e09f91aaf8bcb87217056ed51fdd18f108708771ef543819f4801d57ee6f479cd31739044b6840c6b62c6c1eb5683421f0d7779f62cb19d9585d7344950a33121f7e8003b508aaad1211708d7888bbb61ea727dc7c5b8b178acffd8d75ed4585c4c8159e47ba38bf7a5d571c806fbcbf3cc39fcd5a9e7f08c0eb0891487c4ab4d60e2a711c3d1448aa377b3150917fdf3334aea571d14551e55bdfa1a21284191581bb43914381ac9757cb33bfe58c0cbad04eb95bba93c66c3bc373fa59c1d55e034f16dd953e6a0f915f2c133f7adfd8cfd78f052899efb50564e918ff49968447142b19c5475b886fdf06487214abc0ebd858f60f4764b8bd469079bba1710ba16a2c447f190da5a1b19328159b400b707d846f77b6c95a0fe4500b50a4be0e9068485319596de63d932e43d4727342185a47abc355b222d753ef9dc8407fe964acfdbc075eab5d9933411c5686be9ba28afe50b6d2379da065d48f3070010d577707a858cd126b0959ad31d9811c1a2a6a9b55d3798211b5305f886480d88bd265c2fd0455e8a49cbdf29d24f02832353e889cb6e72d1003b639c5da68a5d858162e462bb72dc0685df8e85b6b496ab47cf592720e3988ac8ea81986f2269bcc03ba1180045d42e39507b3955b71ac86d2e23a757a4b1d0c719e981b68196069d25b941980b0b0f3fb9db62a2fe0e70a810854519a8b39df7c9eaf97ce673e3f7e23c568dc8b0ebdea12ac547349ef259299e3666173c668e8b231bbcc8d0b56c8034d1c56add3209b1b2058a5561b45fe97ea5bacd6432e3f94173268686be143c657261d45e8e9523401da6b3aa0c8e69eaf2d7ce0d03d9176b7d15dcfeab06dba9b505bc4a31d7ad2cf1a32373ec034abbc83f8c66b207f4d3d4aa8e8586c0c2ea93b4589c2b2f03d391957ffad12c328b237f2a56a6a295ea6853f302a5ec1a282d2cb0125ae7b868c7ef9efcb9b22a73f17f61ebde265f11d00239f9ecd2b6c888ef22f30c20bf075b943d009f059163d44fa2aecd885f6005c8efb800dd37ab972d1b7d5d351e94fbfde9e0475897c329228b3170c1bf9a85f5e0f7c3588f2ba3ae4e772171ae85214cc43d7048894f58c92c5a13e9b6c6e1471343fb0aac670e42f5104f63e1cd6ba3bf87ffc5e7fd4dadd9375001789c41c0f146168618e688c6a6bc0a41db1013e450f07b2a38343b652006e99562aac17e4aeb32e71f921dd7d7d375f02782d77694941a5f9b20d2e9d0f45e11ca068e4d0c3a0aec107f0a734f53eaa5966b81b9c83c5400b2373aaa2c2356a968f38fa8c1ebe455dcc4ef5c901b8f6078eb22afd32b1dc4a72c4f2ae2fdc0e0d26e7ea8b3d3c3ffad4fedb723676b415a094d601e32413041f7a20857a9ca8286a42be864db41757c84845f0545d6455801e0810fc85d30d1f4bad3e5b0c0afac7ef8e88681a11f8fe578d437c207e423fcf56e5ea9c137548a84bb1e86ad6ecc9722f9b4c6d63fcd2540ba20118b4dbe30bf232e8e031311361dbaf9007b35e3d2a8190a66781e0a62dd9a2a3ef6c0e48dc6dc29913d598671b469cc69a5e3e0abd71acfec4b393e939ba8cb8cc40d383d5537201759477d166637d3178e2916000efc0dcc0bf0fa2ddf790e2311596451d0159fbb36212976274f05e8adef49d246b1317ef5f2d75f9ae95cf2b54d29558de3e16f9438f73ac281021e9c4aef96f9ad718f70065a726b73eaf90e92cb7d2d8ad97cdf1bdfdca1c77062e687beec1d7c022ca38680a4d7165720b81da0fbc6d2e5f6ccc221;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h55098e9d2476e732bdc2d63e727bbf3515d33621fe4b8faa8d9eae35eafa41b31dab3845305f1fb5c57842a1a03f8891ae0cdc1f22a00fd73ba00cf9f766b3b549769887c385d9c1e0005e8601e691ee55baa5e3b009bca4a6287499e468fb948be859db9194a5d5b1821b811e5827fba0ba1cc77609a494ecae2ff4031cf13854c5f33ba1e27fa775ece1e9d3bd6330c9fb1400532d74402ff0e6a54b822e236bf4ece595a8bf2ad574205fb2bf9778f603a193b74f459eaadbd1c37f66e18fcb868b683a312412b23b1c52f29faa43a3dfaa2339f4ff2e3e5e57532ddd092bce8fdc518114f429552cc4d60e2c45c2a32bfe69de07c4172a2de16e60eb9e89fbea51052f681b7280caed0a110e5755b38d0396f8acdf4f57ab83ca1042968ade6af89e04b005d605c2dfa21a42a1ed22c01b1a266a77fae8b57352cc9167e2a8b7e0c1b9ed2e27a6cfe5ad50058fc397d353b9e0dd427dd3c2e8dc4a9f27a0b1299e7acb43ae9703faecdf165227905b0cae82f9f9c3c871083e9c4be19a92fe1e787698d60d892681bda36117c591d7a4d05afc9de384478d92a16257dd059944ade4b2458a83987849298cc381b18d88fbb73b1355eb887fe5ef920fcf0608a7e7c641f753e2e5dcbb16fc30f4b59273dedaa5137d467bed1b0269309bc57df4b262445a77ae988b0c1759bb5a97f67d59d85e9f91c2553bd815fbb88d93dec569e474ac3cca329bca278a3ca52d1b6039619a4b34d6196c707d58be095c38233c1b6830a62dfb8d532d54a3f37b7d4e7807a1d99b7dcbc803b5b525c532ece3e2f20d4760bd417a5083e348ea7d8e918ac8a66a583b55ba4bd5879074ddf0a6935f6b4e07f1a72eb7a6aba8b5424af5504346028bdae8acda03afa781b9dfc4cc857946f3f8010a256c9c9be8585e56a7f33505de73b4d03ece51579b4c755b299429c41c06972439f798fb216c03f0c8ba5674dd9dd0b59a24b341ffbbf756a7386b23653705b23dc83754d5e9115a5c30786967a6cfb9d7a02e79b3b164b351e6a4236e4589af01e330489c9a45715cc428ab52cfc1a02a1a6dbc27b4be7b7f8da4380ab994a079a49c0b8d07fb531c973c1deb037280a3a8093b9d72608224010aed1d4d82971469231bde65d06cb81bc30521afde319a4ab440a22aa85a24e79ed696a45e7fb79997d9cbefe24db4781012896ea77c725dc6c769d9213906928d838389206dfe87e5ea1ceaedfd9626580b879889cda52185c4f8abbaa0d53e9ef7b165d0db6019118cb44c40057b64c00726081726b1b22cc882ecfa3a5ea3f34c13f04538d7c5741758d0577a99e33c21e791b8202bac89e12c86d4333cc4e56a8163ce5fca6c0a49eb5cc20363ce7dc5782fb32cfe3f259e83af46c015ee14655a7b028d23c0a88bac6f90b246a28fe87530a8e23e02c33c8a31c177bd07ae151e793a076b6e52444065ace0b7ab4c1ff3ae543361cb5a09ae046b363ca41a08918cde7f399f9a9a0017c28aeac52800e89bf93f1a9d6b679fc18a320b55ab35477a5e16f0f05b178ebe6e67fc79cc618932fe0f68c78e2dca33b8551ecce196f40136d723d0e56632e589c578f1649600b2faf8a8bb6ae2d87e51b884bff922cd292ca37197effe010c4012f0dad4018aeb1f044fd36c6cb0f19dec748c37ceaad3b08c8f0739cf931a15f1b3bea7820c949b04ca023bfa1b8b4ab4f7cd11114adb6da609e572efb7e440aa95bb7b9a87f99ed586d899daeb8b34e0e7f6c033d66513cef470cfb5806927b0018bbbf52f1ca78d364fac95379108b84212c3f91077adf4409232c21fb03fadd9586ba59ba362d992653ef10585456b134332402efa98ace76dadc2e93f74d1dcb0b12378dbc7a799f49a139c0cf7108bbd831e8fcdd5b9f838246fadcc8e6c023191f7165837b609f551cf5cb8096e4f79e97f789f79906e71109fbbefab3184962ee5f4b4371bd7ed0fac844720c6d57482fe714312f76aa17e1f73c441315a1d898e3e7e53a4c3e41dcb92b9e34adb061a13d6a2976c55f9689f78f33b158c6cacc3ca02d0e26bcd25ae14bc849acf16013c5794bfe280e76da361495931d8c35aac62b78481c162490362d029befe493be28ea583ccac75a5f38d73f8de56472efa7a3eb17ea4838d32f768d3be4f3aed205b5c7f8dc4ed59338f5d6e414734ef3b9f87a1a5cfd3bb07792523c3e1c823b08a12e8b8917e6937f5083e3269a40333ed5dda52e6b17370e7b9bd1070cf4cc6368a7c58790e96131084d39015125336e164b11c4072d2de4fc283a8e6ea1b36c8ba311f6c839dc85db0fae0990dd5c4001899efe96a77e174e6717307211b9e9ce36cfce9813670fb3b492309eebd7e89ad108c0a622ddfbd3943045c06defb5ec74cc59a934f2bb656bd7e1f790ce5a868395835aba641c3ce64e55a9c266b859bb88a5205f9a302fff13bea79759e46a89dcf0f1db0b7e7ba593fa1373bdb0b1fb5b8ddf067e5139bd57154a7f3cce15972c1490dbc577be731c10c29dad6ddce622eff60f2558baac4d36893214c72e607d8cb236eb6a70e1e15b26f1653355b40a8ffa47ead195a897794d778f76de44bdc985bc5d1b93209f5c9a1c6d6ddd4aee5df58929c5396b6e49b0efab72c9daa653532d8b780492dae3bef4b7da8f569f66ed948cc809036bdbdadb8bfa0e4d97d6eef5459f4c871cda7feca0a2f4a7cb4a6fd395479d10143b52cb1aeabcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8e28a50ac098a1170a305839ea9a4b2059600c0832bcc63243fd8839cec6dfa7da5675abde5133c72c3e889e8693de15233eef50648b57806492dd716bc3c01fab238a6af4b13ac1d524a9a78cc9b5617e6fe4cf22fbc2e09b4b3d6cf909c7b99a3640cc59a9bed4875f904d21f64bc7f782553d6af580b1ef91aba384ade328bacd86f2da37a0bd06ac5e93de648de5d8f4318ef8bed336af3be7e634f1f35ebd53daef1778b5b56a3e0ceb9f642e6294362593876cb1d0c7798ffd6dc96dd6e8ccf81277935b421d87a8382bf252bf7a48698f0c7af65f52f3d9a1173cd3e7c46fd88676fbded78084c12e7668e9594bb88c8cb2eb09bb2c90654a08ac383bde5892beb8ba2bccc2546dc45a32493178f6ef4dffecf569f37ec83e0630f01b4ba07bd10bc4dbb332423b74730d82730ac012906244c842e4dec68fef24fc0e9a7df716fb9c762ec03917c29cb853ed8a07553985656ee5c8fb5d392aaab47fda9d9aef1af2f331a2214f2933f709d4c92b3b29faeae128dba82a26209611a15a92c3300aea3c98b8fc65f7cb16b148691822e41c76488a3344c8171d46c9be0c34e7e2a056c1d66c9e3af8f86277f16d6886323111c08332b2266ac8ba1d67139a061e98e9c3661a6e381301a3be48304bd7315ca2e6068048f768ad4fbf687641e078e712ebb42369813334d5c3e2e6a2e72f1cf5e9fcbfaea141e11c3e7b736e71b9496354a46d3beab8999908e39fd5c6a3caab7e65d9a66f3b4d237d06f2864e1e0b42b73f1e921ec9a0360bfe42716baedabe7627b1d7ec5c9868c67a45111ed30aa836aef5747bafb0bf2f2c052c288f788ff19d499df35ac22696979251947e9422dd2a08de1158b199699f9215e94df040df1ee42bc0c470df0295d086bceef0b8a2e5113dd1961f6fd02de0563457ab030e349407d99aef02d95dbeb4eeffe8545eaa169bc0e430a6debcb0ade3e758e360937788b3a1e8dceed69b4b4e0a3eb50d08cf0b72055b208653f8022f3ff288cbe9944cd68d16305d87c869568d950576648545768430115ce5a21ff9d81a034787b2db79ab3c144f3cdb443de9defbb690e57a2859f61a1e2d44297930d80a19e9b1bc511caea765acb619018ca0f3d59f481f9dac11bfb2736f43e102ee3033f080f5972bab57ec909be5be97fa3f9341b6cc08ddd81f816d3e3d7bff62a47286b66c33d56c3af05c30d38a26ca8b943da526c01e4e2aa856d52791e972fb82b8c53cb347b8f9bdc77445f54b37c1a65535443830a07ac61e79baf90f9095b9f768b8790838cda7801f2074101640f435c13a14a5a872200eee5bf733efa9581c1af94cd1b8c29150f399d79db0261e88a198611cc9084d9233dc4d0b8900c8d8ef0f8a4403786775b3836a5af3255f6356ebf82093eb62011e98918c6a13f0092bd32638f7dfc1d0030b3fd7da8dd399652fadcd80982286918084ab70e695d7544aad0ed07f460f17be8cf64a5329f884394e194b7bb353fa81b9bdf1541d63c7f15959974010fdb9e0bae433dc5173da1960bc567f435b229449ac19778d8932c63cb61049648ae90baf78c3f239110c1b0acad9965331de82a8d2ccffdd7673d61c7422c13733b3d4faf6816d84f856017847a383bb98ab2408196f3138b2c9678e75c6ea86caf627262c293559cfec7ec19554236709791bfbcc3c0b3c2cce58ab2332acc23efa382521f99559d585dd5284d2d657526edd9b4aca02cb02c6f133b7b7582dcba4231fb0cbee1f9cab915915ea8a8ea1dd1d3da64d8df7150fd7a2421b2ac35b66eeb824ec58946e2032f5ae449108aff589a9585d383f035aa8628dea85bc14b2e7466ba3fa52a3eb569b8c9e9f37acb0ca60e43a678f7b359214a3b3b049a39339db6f9cbe8cda01e75a545120d4567e890dcf44ef138b24c8903d8b643c74463efb447d6a1bf4998ed2a769147580b8b2ceeb189364fac2d2e919759c8969b26a3a4f534631d8d14bcfad3af29de3e50675bad48e43d50e703201657bacfbd1ff0d3d0e5a296470ab21a13ba6e9b3483889b3baa3ec76824bf39cc2cac070e0e4ad24f3490659707064a0e7806f125a4788ee021b3d4f5d24a9ddad7b5a93c0bc43d3a4d0a24b2f96fd18a481c5e2e28c1438aee75d00828864e20b4e5fbd909d9555c7683dd4992cc0d5d99a1fdbe8606a0ae452f45fc2ad84e02cfeec9c9c4f4c5d234047a3ca62a7ffacd6c0d75c3c0476cc6e0b5642b1b71fe07cf15b87d97e120ad305015aa6f9f6efe7c28fb793317c65abf565fd7cc24fa08104ecbec5d50330b91966164dfec21b204f41854e373b24c432d3a16fe473fc9509e3c7b1e0ce4af1960809ed3e576c6db56faa0c7751165525b1ed1248088e40ca68c467b07b5dd89b4bbd3c9c0e70328233f40102efa12bc1837cd2bbcac005b286bb5296fa5da2a6725c4a65f2ff88c99d112838e4a896c748a5c231fed3545641646238b8bf0bf45925621d95308c409a7359efb7e7c262a9e7e704c4aab11f64b1a39920e0586591614bc4c7b56dc1ebea3170ba4f3dc3766f07a4e2f23012f99097d0a7bb763f412e6a2c4bf84ce39af8a2b0a01eabc44743298f88380ff1685cea4bc20cc9a9fcea78ccff38bf96c776625a779cbadcde06008d97cd255a8da2dd9aef00b0158cd55831ef8674dac45ba04048a2c1bc645accf880020cc4b260a1c58829da6cae3d62f4c43e54881c2c9f47abcac252d7;
        #1
        $finish();
    end
endmodule
