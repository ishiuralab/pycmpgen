module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    compressor2_1_512_16 compressor2_1_512_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_512_16(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    rowadder2_1_25 rowadder2_1inst(
        .src0({comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [100:0] stage1_0;
   wire [179:0] stage1_1;
   wire [172:0] stage1_2;
   wire [245:0] stage1_3;
   wire [240:0] stage1_4;
   wire [217:0] stage1_5;
   wire [206:0] stage1_6;
   wire [206:0] stage1_7;
   wire [217:0] stage1_8;
   wire [263:0] stage1_9;
   wire [209:0] stage1_10;
   wire [189:0] stage1_11;
   wire [221:0] stage1_12;
   wire [281:0] stage1_13;
   wire [244:0] stage1_14;
   wire [271:0] stage1_15;
   wire [126:0] stage1_16;
   wire [63:0] stage1_17;
   wire [22:0] stage2_0;
   wire [40:0] stage2_1;
   wire [59:0] stage2_2;
   wire [102:0] stage2_3;
   wire [116:0] stage2_4;
   wire [93:0] stage2_5;
   wire [103:0] stage2_6;
   wire [84:0] stage2_7;
   wire [86:0] stage2_8;
   wire [137:0] stage2_9;
   wire [85:0] stage2_10;
   wire [143:0] stage2_11;
   wire [84:0] stage2_12;
   wire [140:0] stage2_13;
   wire [124:0] stage2_14;
   wire [84:0] stage2_15;
   wire [104:0] stage2_16;
   wire [61:0] stage2_17;
   wire [25:0] stage2_18;
   wire [10:0] stage2_19;
   wire [5:0] stage3_0;
   wire [11:0] stage3_1;
   wire [16:0] stage3_2;
   wire [28:0] stage3_3;
   wire [39:0] stage3_4;
   wire [47:0] stage3_5;
   wire [37:0] stage3_6;
   wire [45:0] stage3_7;
   wire [40:0] stage3_8;
   wire [51:0] stage3_9;
   wire [63:0] stage3_10;
   wire [60:0] stage3_11;
   wire [52:0] stage3_12;
   wire [41:0] stage3_13;
   wire [57:0] stage3_14;
   wire [56:0] stage3_15;
   wire [49:0] stage3_16;
   wire [31:0] stage3_17;
   wire [25:0] stage3_18;
   wire [13:0] stage3_19;
   wire [5:0] stage3_20;
   wire [1:0] stage3_21;
   wire [5:0] stage4_0;
   wire [1:0] stage4_1;
   wire [10:0] stage4_2;
   wire [10:0] stage4_3;
   wire [26:0] stage4_4;
   wire [14:0] stage4_5;
   wire [21:0] stage4_6;
   wire [16:0] stage4_7;
   wire [25:0] stage4_8;
   wire [24:0] stage4_9;
   wire [37:0] stage4_10;
   wire [21:0] stage4_11;
   wire [23:0] stage4_12;
   wire [25:0] stage4_13;
   wire [18:0] stage4_14;
   wire [21:0] stage4_15;
   wire [30:0] stage4_16;
   wire [21:0] stage4_17;
   wire [12:0] stage4_18;
   wire [10:0] stage4_19;
   wire [11:0] stage4_20;
   wire [3:0] stage4_21;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [6:0] stage5_2;
   wire [5:0] stage5_3;
   wire [12:0] stage5_4;
   wire [7:0] stage5_5;
   wire [16:0] stage5_6;
   wire [5:0] stage5_7;
   wire [9:0] stage5_8;
   wire [8:0] stage5_9;
   wire [14:0] stage5_10;
   wire [12:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [11:0] stage5_14;
   wire [14:0] stage5_15;
   wire [16:0] stage5_16;
   wire [6:0] stage5_17;
   wire [8:0] stage5_18;
   wire [8:0] stage5_19;
   wire [5:0] stage5_20;
   wire [3:0] stage5_21;
   wire [1:0] stage5_22;
   wire [0:0] stage5_23;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [6:0] stage6_4;
   wire [2:0] stage6_5;
   wire [5:0] stage6_6;
   wire [4:0] stage6_7;
   wire [3:0] stage6_8;
   wire [8:0] stage6_9;
   wire [9:0] stage6_10;
   wire [2:0] stage6_11;
   wire [3:0] stage6_12;
   wire [7:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [7:0] stage6_20;
   wire [4:0] stage6_21;
   wire [1:0] stage6_22;
   wire [0:0] stage6_23;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [2:0] stage7_5;
   wire [0:0] stage7_6;
   wire [5:0] stage7_7;
   wire [0:0] stage7_8;
   wire [2:0] stage7_9;
   wire [6:0] stage7_10;
   wire [2:0] stage7_11;
   wire [1:0] stage7_12;
   wire [2:0] stage7_13;
   wire [4:0] stage7_14;
   wire [3:0] stage7_15;
   wire [1:0] stage7_16;
   wire [6:0] stage7_17;
   wire [2:0] stage7_18;
   wire [1:0] stage7_19;
   wire [3:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [0:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [0:0] stage8_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_1[13]},
      {stage0_2[13]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[14]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[15]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[16]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[17]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[110], stage0_0[111], stage0_0[112]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[18]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[19]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[20]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[21]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[22]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[23]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[128], stage0_0[129], stage0_0[130]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[24]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[25]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[134], stage0_0[135], stage0_0[136]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[26]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[137], stage0_0[138], stage0_0[139]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[27]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[140], stage0_0[141], stage0_0[142]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[28]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[143], stage0_0[144], stage0_0[145]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[29]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[30]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[31]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[32]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[155], stage0_0[156], stage0_0[157]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[33]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[158], stage0_0[159], stage0_0[160]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[34]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[161], stage0_0[162], stage0_0[163]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[35]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[164], stage0_0[165], stage0_0[166]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[36]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[167], stage0_0[168], stage0_0[169]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[37]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[170], stage0_0[171], stage0_0[172]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[38]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[173], stage0_0[174], stage0_0[175]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[39]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[176], stage0_0[177], stage0_0[178]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[40]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[179], stage0_0[180], stage0_0[181]},
      {stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181]},
      {stage0_2[41]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[182], stage0_0[183], stage0_0[184]},
      {stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187]},
      {stage0_2[42]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[185], stage0_0[186], stage0_0[187]},
      {stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193]},
      {stage0_2[43]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[188], stage0_0[189], stage0_0[190]},
      {stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199]},
      {stage0_2[44]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[31],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[32],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[33],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[34],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[35],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[36],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[37],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[38],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[39],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[40],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[41],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[42],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[43],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[44],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[45],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[46],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[47],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[48],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[49],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[50],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[51],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[52],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[53],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[54],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[55],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[56],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[57],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[58],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[59],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[60],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[61],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[62],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[63],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[64],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[65],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[66],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[67],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[68],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[69],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[70],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[71],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[72],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[73],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[74],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[75],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[76],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[77],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[78],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[79],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489], stage0_0[490]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[80],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[81],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[82],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507], stage0_0[508]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[83],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[0],stage1_4[84],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[1],stage1_4[85],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[2],stage1_4[86],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[3],stage1_4[87],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[4],stage1_4[88],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[5],stage1_4[89],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[6],stage1_4[90],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[7],stage1_4[91],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[8],stage1_4[92],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[9],stage1_4[93],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[10],stage1_4[94],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[11],stage1_4[95],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[12],stage1_4[96],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[13],stage1_4[97],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[14],stage1_4[98],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[15],stage1_4[99],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[16],stage1_4[100],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[17],stage1_4[101],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[18],stage1_4[102],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[19],stage1_4[103],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[20],stage1_4[104],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[21],stage1_4[105],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[22],stage1_4[106],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[23],stage1_4[107],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[24],stage1_4[108],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[25],stage1_4[109],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[26],stage1_4[110],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[27],stage1_4[111],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[28],stage1_4[112],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[29],stage1_4[113],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[30],stage1_4[114],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[31],stage1_4[115],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[32],stage1_4[116],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[33],stage1_4[117],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[34],stage1_4[118],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[35],stage1_4[119],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[36],stage1_4[120],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[37],stage1_4[121],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[38],stage1_4[122],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[39],stage1_4[123],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[40],stage1_4[124],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[41],stage1_4[125],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[42],stage1_4[126],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[43],stage1_4[127],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[44],stage1_4[128],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[45],stage1_4[129],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[46],stage1_4[130],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[47],stage1_4[131],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[48],stage1_4[132],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[49],stage1_4[133],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[50],stage1_4[134],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397]},
      {stage0_3[307]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[51],stage1_4[135],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage0_3[308]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[52],stage1_4[136],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_3[309]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[53],stage1_4[137],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412]},
      {stage0_3[310]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[54],stage1_4[138],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417]},
      {stage0_3[311]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[55],stage1_4[139],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage0_3[312]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[56],stage1_4[140],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427]},
      {stage0_3[313]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[57],stage1_4[141],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432]},
      {stage0_3[314]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[58],stage1_4[142],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_3[315]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[59],stage1_4[143],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442]},
      {stage0_3[316]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[60],stage1_4[144],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447]},
      {stage0_3[317]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[61],stage1_4[145],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[448], stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452]},
      {stage0_3[318]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[62],stage1_4[146],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[453], stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457]},
      {stage0_3[319]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[63],stage1_4[147],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462]},
      {stage0_3[320]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[64],stage1_4[148],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_3[321]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[65],stage1_4[149],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472]},
      {stage0_3[322]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[66],stage1_4[150],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[473], stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477]},
      {stage0_3[323]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[67],stage1_4[151],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_2[478], stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482]},
      {stage0_3[324]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[68],stage1_4[152],stage1_3[166],stage1_2[166]}
   );
   gpc615_5 gpc167 (
      {stage0_2[483], stage0_2[484], stage0_2[485], stage0_2[486], stage0_2[487]},
      {stage0_3[325]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[69],stage1_4[153],stage1_3[167],stage1_2[167]}
   );
   gpc615_5 gpc168 (
      {stage0_2[488], stage0_2[489], stage0_2[490], stage0_2[491], stage0_2[492]},
      {stage0_3[326]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[70],stage1_4[154],stage1_3[168],stage1_2[168]}
   );
   gpc615_5 gpc169 (
      {stage0_2[493], stage0_2[494], stage0_2[495], stage0_2[496], stage0_2[497]},
      {stage0_3[327]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[71],stage1_4[155],stage1_3[169],stage1_2[169]}
   );
   gpc615_5 gpc170 (
      {stage0_2[498], stage0_2[499], stage0_2[500], stage0_2[501], stage0_2[502]},
      {stage0_3[328]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[72],stage1_4[156],stage1_3[170],stage1_2[170]}
   );
   gpc615_5 gpc171 (
      {stage0_2[503], stage0_2[504], stage0_2[505], stage0_2[506], stage0_2[507]},
      {stage0_3[329]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[73],stage1_4[157],stage1_3[171],stage1_2[171]}
   );
   gpc615_5 gpc172 (
      {stage0_2[508], stage0_2[509], stage0_2[510], stage0_2[511], 1'b0},
      {stage0_3[330]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[74],stage1_4[158],stage1_3[172],stage1_2[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[75],stage1_4[159],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[76],stage1_4[160],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[77],stage1_4[161],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[78],stage1_4[162],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[79],stage1_4[163],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[80],stage1_4[164],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[81],stage1_4[165],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[82],stage1_4[166],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[83],stage1_4[167],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[84],stage1_4[168],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[85],stage1_4[169],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[86],stage1_4[170],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[87],stage1_4[171],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[88],stage1_4[172],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[89],stage1_4[173],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[90],stage1_4[174],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[91],stage1_4[175],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[92],stage1_4[176],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[93],stage1_4[177],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[94],stage1_4[178],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[95],stage1_4[179],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[96],stage1_4[180],stage1_3[194]}
   );
   gpc615_5 gpc195 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[97],stage1_4[181],stage1_3[195]}
   );
   gpc615_5 gpc196 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[98],stage1_4[182],stage1_3[196]}
   );
   gpc615_5 gpc197 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[99],stage1_4[183],stage1_3[197]}
   );
   gpc615_5 gpc198 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[100],stage1_4[184],stage1_3[198]}
   );
   gpc615_5 gpc199 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[101],stage1_4[185],stage1_3[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[27],stage1_6[56],stage1_5[102],stage1_4[186]}
   );
   gpc606_5 gpc201 (
      {stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[28],stage1_6[57],stage1_5[103],stage1_4[187]}
   );
   gpc606_5 gpc202 (
      {stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[29],stage1_6[58],stage1_5[104],stage1_4[188]}
   );
   gpc606_5 gpc203 (
      {stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[30],stage1_6[59],stage1_5[105],stage1_4[189]}
   );
   gpc606_5 gpc204 (
      {stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[31],stage1_6[60],stage1_5[106],stage1_4[190]}
   );
   gpc606_5 gpc205 (
      {stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[32],stage1_6[61],stage1_5[107],stage1_4[191]}
   );
   gpc606_5 gpc206 (
      {stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[33],stage1_6[62],stage1_5[108],stage1_4[192]}
   );
   gpc606_5 gpc207 (
      {stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[34],stage1_6[63],stage1_5[109],stage1_4[193]}
   );
   gpc606_5 gpc208 (
      {stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[35],stage1_6[64],stage1_5[110],stage1_4[194]}
   );
   gpc606_5 gpc209 (
      {stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[36],stage1_6[65],stage1_5[111],stage1_4[195]}
   );
   gpc606_5 gpc210 (
      {stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[37],stage1_6[66],stage1_5[112],stage1_4[196]}
   );
   gpc606_5 gpc211 (
      {stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[38],stage1_6[67],stage1_5[113],stage1_4[197]}
   );
   gpc606_5 gpc212 (
      {stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[39],stage1_6[68],stage1_5[114],stage1_4[198]}
   );
   gpc606_5 gpc213 (
      {stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[40],stage1_6[69],stage1_5[115],stage1_4[199]}
   );
   gpc606_5 gpc214 (
      {stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[41],stage1_6[70],stage1_5[116],stage1_4[200]}
   );
   gpc606_5 gpc215 (
      {stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[42],stage1_6[71],stage1_5[117],stage1_4[201]}
   );
   gpc606_5 gpc216 (
      {stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[43],stage1_6[72],stage1_5[118],stage1_4[202]}
   );
   gpc606_5 gpc217 (
      {stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[44],stage1_6[73],stage1_5[119],stage1_4[203]}
   );
   gpc606_5 gpc218 (
      {stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[45],stage1_6[74],stage1_5[120],stage1_4[204]}
   );
   gpc606_5 gpc219 (
      {stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[46],stage1_6[75],stage1_5[121],stage1_4[205]}
   );
   gpc606_5 gpc220 (
      {stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[47],stage1_6[76],stage1_5[122],stage1_4[206]}
   );
   gpc606_5 gpc221 (
      {stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[48],stage1_6[77],stage1_5[123],stage1_4[207]}
   );
   gpc606_5 gpc222 (
      {stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[49],stage1_6[78],stage1_5[124],stage1_4[208]}
   );
   gpc606_5 gpc223 (
      {stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[50],stage1_6[79],stage1_5[125],stage1_4[209]}
   );
   gpc606_5 gpc224 (
      {stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[51],stage1_6[80],stage1_5[126],stage1_4[210]}
   );
   gpc606_5 gpc225 (
      {stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[52],stage1_6[81],stage1_5[127],stage1_4[211]}
   );
   gpc606_5 gpc226 (
      {stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[53],stage1_6[82],stage1_5[128],stage1_4[212]}
   );
   gpc606_5 gpc227 (
      {stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[54],stage1_6[83],stage1_5[129],stage1_4[213]}
   );
   gpc606_5 gpc228 (
      {stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[55],stage1_6[84],stage1_5[130],stage1_4[214]}
   );
   gpc606_5 gpc229 (
      {stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[56],stage1_6[85],stage1_5[131],stage1_4[215]}
   );
   gpc606_5 gpc230 (
      {stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[57],stage1_6[86],stage1_5[132],stage1_4[216]}
   );
   gpc606_5 gpc231 (
      {stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[58],stage1_6[87],stage1_5[133],stage1_4[217]}
   );
   gpc606_5 gpc232 (
      {stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[59],stage1_6[88],stage1_5[134],stage1_4[218]}
   );
   gpc606_5 gpc233 (
      {stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[60],stage1_6[89],stage1_5[135],stage1_4[219]}
   );
   gpc606_5 gpc234 (
      {stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[61],stage1_6[90],stage1_5[136],stage1_4[220]}
   );
   gpc606_5 gpc235 (
      {stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[62],stage1_6[91],stage1_5[137],stage1_4[221]}
   );
   gpc615_5 gpc236 (
      {stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_5[162]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[63],stage1_6[92],stage1_5[138],stage1_4[222]}
   );
   gpc615_5 gpc237 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_5[163]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[64],stage1_6[93],stage1_5[139],stage1_4[223]}
   );
   gpc615_5 gpc238 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431]},
      {stage0_5[164]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[65],stage1_6[94],stage1_5[140],stage1_4[224]}
   );
   gpc615_5 gpc239 (
      {stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_5[165]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[66],stage1_6[95],stage1_5[141],stage1_4[225]}
   );
   gpc615_5 gpc240 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_5[166]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[67],stage1_6[96],stage1_5[142],stage1_4[226]}
   );
   gpc615_5 gpc241 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446]},
      {stage0_5[167]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[68],stage1_6[97],stage1_5[143],stage1_4[227]}
   );
   gpc615_5 gpc242 (
      {stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_5[168]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[69],stage1_6[98],stage1_5[144],stage1_4[228]}
   );
   gpc615_5 gpc243 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_5[169]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[70],stage1_6[99],stage1_5[145],stage1_4[229]}
   );
   gpc615_5 gpc244 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461]},
      {stage0_5[170]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[71],stage1_6[100],stage1_5[146],stage1_4[230]}
   );
   gpc615_5 gpc245 (
      {stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_5[171]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[72],stage1_6[101],stage1_5[147],stage1_4[231]}
   );
   gpc615_5 gpc246 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_5[172]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[73],stage1_6[102],stage1_5[148],stage1_4[232]}
   );
   gpc615_5 gpc247 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[173]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[74],stage1_6[103],stage1_5[149],stage1_4[233]}
   );
   gpc615_5 gpc248 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[174]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[75],stage1_6[104],stage1_5[150],stage1_4[234]}
   );
   gpc615_5 gpc249 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[175]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[76],stage1_6[105],stage1_5[151],stage1_4[235]}
   );
   gpc615_5 gpc250 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[176]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[77],stage1_6[106],stage1_5[152],stage1_4[236]}
   );
   gpc615_5 gpc251 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[177]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[78],stage1_6[107],stage1_5[153],stage1_4[237]}
   );
   gpc615_5 gpc252 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[178]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[79],stage1_6[108],stage1_5[154],stage1_4[238]}
   );
   gpc615_5 gpc253 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[179]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[80],stage1_6[109],stage1_5[155],stage1_4[239]}
   );
   gpc615_5 gpc254 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[180]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[81],stage1_6[110],stage1_5[156],stage1_4[240]}
   );
   gpc606_5 gpc255 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[82],stage1_6[111],stage1_5[157]}
   );
   gpc606_5 gpc256 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[83],stage1_6[112],stage1_5[158]}
   );
   gpc606_5 gpc257 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[84],stage1_6[113],stage1_5[159]}
   );
   gpc606_5 gpc258 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[85],stage1_6[114],stage1_5[160]}
   );
   gpc606_5 gpc259 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[86],stage1_6[115],stage1_5[161]}
   );
   gpc606_5 gpc260 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[87],stage1_6[116],stage1_5[162]}
   );
   gpc606_5 gpc261 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[88],stage1_6[117],stage1_5[163]}
   );
   gpc606_5 gpc262 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[89],stage1_6[118],stage1_5[164]}
   );
   gpc606_5 gpc263 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[90],stage1_6[119],stage1_5[165]}
   );
   gpc606_5 gpc264 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[91],stage1_6[120],stage1_5[166]}
   );
   gpc606_5 gpc265 (
      {stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[92],stage1_6[121],stage1_5[167]}
   );
   gpc606_5 gpc266 (
      {stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[93],stage1_6[122],stage1_5[168]}
   );
   gpc606_5 gpc267 (
      {stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[94],stage1_6[123],stage1_5[169]}
   );
   gpc606_5 gpc268 (
      {stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[95],stage1_6[124],stage1_5[170]}
   );
   gpc606_5 gpc269 (
      {stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[96],stage1_6[125],stage1_5[171]}
   );
   gpc606_5 gpc270 (
      {stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[97],stage1_6[126],stage1_5[172]}
   );
   gpc606_5 gpc271 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[98],stage1_6[127],stage1_5[173]}
   );
   gpc606_5 gpc272 (
      {stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[99],stage1_6[128],stage1_5[174]}
   );
   gpc606_5 gpc273 (
      {stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[100],stage1_6[129],stage1_5[175]}
   );
   gpc606_5 gpc274 (
      {stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[101],stage1_6[130],stage1_5[176]}
   );
   gpc606_5 gpc275 (
      {stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[102],stage1_6[131],stage1_5[177]}
   );
   gpc606_5 gpc276 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[103],stage1_6[132],stage1_5[178]}
   );
   gpc606_5 gpc277 (
      {stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[104],stage1_6[133],stage1_5[179]}
   );
   gpc606_5 gpc278 (
      {stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[105],stage1_6[134],stage1_5[180]}
   );
   gpc606_5 gpc279 (
      {stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[106],stage1_6[135],stage1_5[181]}
   );
   gpc606_5 gpc280 (
      {stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[107],stage1_6[136],stage1_5[182]}
   );
   gpc606_5 gpc281 (
      {stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[108],stage1_6[137],stage1_5[183]}
   );
   gpc606_5 gpc282 (
      {stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[109],stage1_6[138],stage1_5[184]}
   );
   gpc606_5 gpc283 (
      {stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[110],stage1_6[139],stage1_5[185]}
   );
   gpc606_5 gpc284 (
      {stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[111],stage1_6[140],stage1_5[186]}
   );
   gpc606_5 gpc285 (
      {stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[112],stage1_6[141],stage1_5[187]}
   );
   gpc606_5 gpc286 (
      {stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[113],stage1_6[142],stage1_5[188]}
   );
   gpc606_5 gpc287 (
      {stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[114],stage1_6[143],stage1_5[189]}
   );
   gpc606_5 gpc288 (
      {stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[115],stage1_6[144],stage1_5[190]}
   );
   gpc606_5 gpc289 (
      {stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[116],stage1_6[145],stage1_5[191]}
   );
   gpc606_5 gpc290 (
      {stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[117],stage1_6[146],stage1_5[192]}
   );
   gpc606_5 gpc291 (
      {stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[118],stage1_6[147],stage1_5[193]}
   );
   gpc606_5 gpc292 (
      {stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[119],stage1_6[148],stage1_5[194]}
   );
   gpc606_5 gpc293 (
      {stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[120],stage1_6[149],stage1_5[195]}
   );
   gpc606_5 gpc294 (
      {stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[121],stage1_6[150],stage1_5[196]}
   );
   gpc606_5 gpc295 (
      {stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[122],stage1_6[151],stage1_5[197]}
   );
   gpc606_5 gpc296 (
      {stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[123],stage1_6[152],stage1_5[198]}
   );
   gpc606_5 gpc297 (
      {stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[124],stage1_6[153],stage1_5[199]}
   );
   gpc606_5 gpc298 (
      {stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[125],stage1_6[154],stage1_5[200]}
   );
   gpc606_5 gpc299 (
      {stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[126],stage1_6[155],stage1_5[201]}
   );
   gpc606_5 gpc300 (
      {stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[127],stage1_6[156],stage1_5[202]}
   );
   gpc606_5 gpc301 (
      {stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[128],stage1_6[157],stage1_5[203]}
   );
   gpc606_5 gpc302 (
      {stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[129],stage1_6[158],stage1_5[204]}
   );
   gpc606_5 gpc303 (
      {stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[130],stage1_6[159],stage1_5[205]}
   );
   gpc606_5 gpc304 (
      {stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[131],stage1_6[160],stage1_5[206]}
   );
   gpc606_5 gpc305 (
      {stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[105],stage1_7[132],stage1_6[161],stage1_5[207]}
   );
   gpc606_5 gpc306 (
      {stage0_5[487], stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[106],stage1_7[133],stage1_6[162],stage1_5[208]}
   );
   gpc606_5 gpc307 (
      {stage0_5[493], stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[107],stage1_7[134],stage1_6[163],stage1_5[209]}
   );
   gpc606_5 gpc308 (
      {stage0_5[499], stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[108],stage1_7[135],stage1_6[164],stage1_5[210]}
   );
   gpc615_5 gpc309 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[324]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[54],stage1_8[109],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc310 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[325]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[55],stage1_8[110],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc311 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[326]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[56],stage1_8[111],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc312 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[327]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[57],stage1_8[112],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc313 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[328]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[58],stage1_8[113],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc314 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[329]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[59],stage1_8[114],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc315 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[330]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[60],stage1_8[115],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc316 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[331]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[61],stage1_8[116],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc317 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[332]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[62],stage1_8[117],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc318 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[333]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[63],stage1_8[118],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc319 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[334]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[64],stage1_8[119],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc320 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[335]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[65],stage1_8[120],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc321 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[336]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[66],stage1_8[121],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc322 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[337]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[67],stage1_8[122],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc323 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[338]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[68],stage1_8[123],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc324 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[339]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[69],stage1_8[124],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc325 (
      {stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414]},
      {stage0_7[340]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[70],stage1_8[125],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc326 (
      {stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage0_7[341]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[71],stage1_8[126],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc327 (
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424]},
      {stage0_7[342]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[72],stage1_8[127],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc328 (
      {stage0_6[425], stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429]},
      {stage0_7[343]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[73],stage1_8[128],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc329 (
      {stage0_6[430], stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434]},
      {stage0_7[344]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[74],stage1_8[129],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc330 (
      {stage0_6[435], stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439]},
      {stage0_7[345]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[75],stage1_8[130],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc331 (
      {stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444]},
      {stage0_7[346]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[76],stage1_8[131],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc332 (
      {stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage0_7[347]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[77],stage1_8[132],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc333 (
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454]},
      {stage0_7[348]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[78],stage1_8[133],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc334 (
      {stage0_6[455], stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459]},
      {stage0_7[349]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[79],stage1_8[134],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc335 (
      {stage0_6[460], stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464]},
      {stage0_7[350]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[80],stage1_8[135],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc336 (
      {stage0_6[465], stage0_6[466], stage0_6[467], stage0_6[468], stage0_6[469]},
      {stage0_7[351]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[81],stage1_8[136],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc337 (
      {stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473], stage0_6[474]},
      {stage0_7[352]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[82],stage1_8[137],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc338 (
      {stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_7[353]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[83],stage1_8[138],stage1_7[165],stage1_6[194]}
   );
   gpc615_5 gpc339 (
      {stage0_6[480], stage0_6[481], stage0_6[482], stage0_6[483], stage0_6[484]},
      {stage0_7[354]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[84],stage1_8[139],stage1_7[166],stage1_6[195]}
   );
   gpc615_5 gpc340 (
      {stage0_6[485], stage0_6[486], stage0_6[487], stage0_6[488], stage0_6[489]},
      {stage0_7[355]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[85],stage1_8[140],stage1_7[167],stage1_6[196]}
   );
   gpc615_5 gpc341 (
      {stage0_6[490], stage0_6[491], stage0_6[492], stage0_6[493], stage0_6[494]},
      {stage0_7[356]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[86],stage1_8[141],stage1_7[168],stage1_6[197]}
   );
   gpc615_5 gpc342 (
      {stage0_6[495], stage0_6[496], stage0_6[497], stage0_6[498], stage0_6[499]},
      {stage0_7[357]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[87],stage1_8[142],stage1_7[169],stage1_6[198]}
   );
   gpc615_5 gpc343 (
      {stage0_6[500], stage0_6[501], stage0_6[502], stage0_6[503], stage0_6[504]},
      {stage0_7[358]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[88],stage1_8[143],stage1_7[170],stage1_6[199]}
   );
   gpc606_5 gpc344 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[35],stage1_9[89],stage1_8[144],stage1_7[171]}
   );
   gpc606_5 gpc345 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[36],stage1_9[90],stage1_8[145],stage1_7[172]}
   );
   gpc606_5 gpc346 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[37],stage1_9[91],stage1_8[146],stage1_7[173]}
   );
   gpc606_5 gpc347 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[38],stage1_9[92],stage1_8[147],stage1_7[174]}
   );
   gpc606_5 gpc348 (
      {stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[39],stage1_9[93],stage1_8[148],stage1_7[175]}
   );
   gpc606_5 gpc349 (
      {stage0_7[389], stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[40],stage1_9[94],stage1_8[149],stage1_7[176]}
   );
   gpc606_5 gpc350 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[41],stage1_9[95],stage1_8[150],stage1_7[177]}
   );
   gpc606_5 gpc351 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[42],stage1_9[96],stage1_8[151],stage1_7[178]}
   );
   gpc606_5 gpc352 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[43],stage1_9[97],stage1_8[152],stage1_7[179]}
   );
   gpc606_5 gpc353 (
      {stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[44],stage1_9[98],stage1_8[153],stage1_7[180]}
   );
   gpc606_5 gpc354 (
      {stage0_7[419], stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[45],stage1_9[99],stage1_8[154],stage1_7[181]}
   );
   gpc606_5 gpc355 (
      {stage0_7[425], stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[46],stage1_9[100],stage1_8[155],stage1_7[182]}
   );
   gpc606_5 gpc356 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[47],stage1_9[101],stage1_8[156],stage1_7[183]}
   );
   gpc606_5 gpc357 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[48],stage1_9[102],stage1_8[157],stage1_7[184]}
   );
   gpc606_5 gpc358 (
      {stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[49],stage1_9[103],stage1_8[158],stage1_7[185]}
   );
   gpc606_5 gpc359 (
      {stage0_7[449], stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[50],stage1_9[104],stage1_8[159],stage1_7[186]}
   );
   gpc606_5 gpc360 (
      {stage0_7[455], stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[51],stage1_9[105],stage1_8[160],stage1_7[187]}
   );
   gpc615_5 gpc361 (
      {stage0_7[461], stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465]},
      {stage0_8[210]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[52],stage1_9[106],stage1_8[161],stage1_7[188]}
   );
   gpc615_5 gpc362 (
      {stage0_7[466], stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470]},
      {stage0_8[211]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[53],stage1_9[107],stage1_8[162],stage1_7[189]}
   );
   gpc615_5 gpc363 (
      {stage0_7[471], stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475]},
      {stage0_8[212]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[54],stage1_9[108],stage1_8[163],stage1_7[190]}
   );
   gpc615_5 gpc364 (
      {stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480]},
      {stage0_8[213]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[55],stage1_9[109],stage1_8[164],stage1_7[191]}
   );
   gpc615_5 gpc365 (
      {stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_8[214]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[56],stage1_9[110],stage1_8[165],stage1_7[192]}
   );
   gpc615_5 gpc366 (
      {stage0_7[486], stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490]},
      {stage0_8[215]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[57],stage1_9[111],stage1_8[166],stage1_7[193]}
   );
   gpc615_5 gpc367 (
      {stage0_7[491], stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495]},
      {stage0_8[216]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[58],stage1_9[112],stage1_8[167],stage1_7[194]}
   );
   gpc615_5 gpc368 (
      {stage0_7[496], stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500]},
      {stage0_8[217]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[59],stage1_9[113],stage1_8[168],stage1_7[195]}
   );
   gpc606_5 gpc369 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[25],stage1_10[60],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc370 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[26],stage1_10[61],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc371 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[27],stage1_10[62],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc372 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[28],stage1_10[63],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc373 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[29],stage1_10[64],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc374 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[30],stage1_10[65],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc375 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[31],stage1_10[66],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc376 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[32],stage1_10[67],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc377 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[33],stage1_10[68],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc378 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[34],stage1_10[69],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc379 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[35],stage1_10[70],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc380 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[36],stage1_10[71],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc381 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[37],stage1_10[72],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc382 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[38],stage1_10[73],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc383 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[39],stage1_10[74],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc384 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[40],stage1_10[75],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc385 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[41],stage1_10[76],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc386 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[42],stage1_10[77],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc387 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[43],stage1_10[78],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc388 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[44],stage1_10[79],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc389 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[45],stage1_10[80],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc390 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[46],stage1_10[81],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc391 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[47],stage1_10[82],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc392 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[48],stage1_10[83],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc393 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[49],stage1_10[84],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc394 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[50],stage1_10[85],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc395 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[51],stage1_10[86],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc396 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[52],stage1_10[87],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc397 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[53],stage1_10[88],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc398 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[54],stage1_10[89],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc399 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[55],stage1_10[90],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc400 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[56],stage1_10[91],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc401 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[57],stage1_10[92],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc402 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[58],stage1_10[93],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc403 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[59],stage1_10[94],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc404 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[60],stage1_10[95],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc405 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[61],stage1_10[96],stage1_9[150],stage1_8[205]}
   );
   gpc606_5 gpc406 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[62],stage1_10[97],stage1_9[151],stage1_8[206]}
   );
   gpc606_5 gpc407 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[63],stage1_10[98],stage1_9[152],stage1_8[207]}
   );
   gpc606_5 gpc408 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[64],stage1_10[99],stage1_9[153],stage1_8[208]}
   );
   gpc606_5 gpc409 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[65],stage1_10[100],stage1_9[154],stage1_8[209]}
   );
   gpc606_5 gpc410 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[66],stage1_10[101],stage1_9[155],stage1_8[210]}
   );
   gpc606_5 gpc411 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[67],stage1_10[102],stage1_9[156],stage1_8[211]}
   );
   gpc606_5 gpc412 (
      {stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480], stage0_8[481]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[68],stage1_10[103],stage1_9[157],stage1_8[212]}
   );
   gpc606_5 gpc413 (
      {stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486], stage0_8[487]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[69],stage1_10[104],stage1_9[158],stage1_8[213]}
   );
   gpc606_5 gpc414 (
      {stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492], stage0_8[493]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[70],stage1_10[105],stage1_9[159],stage1_8[214]}
   );
   gpc606_5 gpc415 (
      {stage0_8[494], stage0_8[495], stage0_8[496], stage0_8[497], stage0_8[498], stage0_8[499]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[71],stage1_10[106],stage1_9[160],stage1_8[215]}
   );
   gpc606_5 gpc416 (
      {stage0_8[500], stage0_8[501], stage0_8[502], stage0_8[503], stage0_8[504], stage0_8[505]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[72],stage1_10[107],stage1_9[161],stage1_8[216]}
   );
   gpc606_5 gpc417 (
      {stage0_8[506], stage0_8[507], stage0_8[508], stage0_8[509], stage0_8[510], stage0_8[511]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[73],stage1_10[108],stage1_9[162],stage1_8[217]}
   );
   gpc606_5 gpc418 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[49],stage1_11[74],stage1_10[109],stage1_9[163]}
   );
   gpc615_5 gpc419 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[294]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[50],stage1_11[75],stage1_10[110],stage1_9[164]}
   );
   gpc615_5 gpc420 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[295]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[51],stage1_11[76],stage1_10[111],stage1_9[165]}
   );
   gpc615_5 gpc421 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[296]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[52],stage1_11[77],stage1_10[112],stage1_9[166]}
   );
   gpc615_5 gpc422 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[297]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[53],stage1_11[78],stage1_10[113],stage1_9[167]}
   );
   gpc615_5 gpc423 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[298]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[54],stage1_11[79],stage1_10[114],stage1_9[168]}
   );
   gpc615_5 gpc424 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[299]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[55],stage1_11[80],stage1_10[115],stage1_9[169]}
   );
   gpc615_5 gpc425 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[300]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[56],stage1_11[81],stage1_10[116],stage1_9[170]}
   );
   gpc615_5 gpc426 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[301]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[57],stage1_11[82],stage1_10[117],stage1_9[171]}
   );
   gpc615_5 gpc427 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[302]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[58],stage1_11[83],stage1_10[118],stage1_9[172]}
   );
   gpc615_5 gpc428 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[303]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[59],stage1_11[84],stage1_10[119],stage1_9[173]}
   );
   gpc615_5 gpc429 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[304]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[60],stage1_11[85],stage1_10[120],stage1_9[174]}
   );
   gpc615_5 gpc430 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[305]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[61],stage1_11[86],stage1_10[121],stage1_9[175]}
   );
   gpc615_5 gpc431 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[306]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[62],stage1_11[87],stage1_10[122],stage1_9[176]}
   );
   gpc615_5 gpc432 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[307]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[63],stage1_11[88],stage1_10[123],stage1_9[177]}
   );
   gpc615_5 gpc433 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[308]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[64],stage1_11[89],stage1_10[124],stage1_9[178]}
   );
   gpc615_5 gpc434 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[309]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[65],stage1_11[90],stage1_10[125],stage1_9[179]}
   );
   gpc615_5 gpc435 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[310]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[66],stage1_11[91],stage1_10[126],stage1_9[180]}
   );
   gpc615_5 gpc436 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[311]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[67],stage1_11[92],stage1_10[127],stage1_9[181]}
   );
   gpc615_5 gpc437 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[312]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[68],stage1_11[93],stage1_10[128],stage1_9[182]}
   );
   gpc615_5 gpc438 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[313]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[69],stage1_11[94],stage1_10[129],stage1_9[183]}
   );
   gpc615_5 gpc439 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_10[314]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[70],stage1_11[95],stage1_10[130],stage1_9[184]}
   );
   gpc615_5 gpc440 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265]},
      {stage0_10[315]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[71],stage1_11[96],stage1_10[131],stage1_9[185]}
   );
   gpc615_5 gpc441 (
      {stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_10[316]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[72],stage1_11[97],stage1_10[132],stage1_9[186]}
   );
   gpc615_5 gpc442 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_10[317]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[73],stage1_11[98],stage1_10[133],stage1_9[187]}
   );
   gpc615_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280]},
      {stage0_10[318]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[74],stage1_11[99],stage1_10[134],stage1_9[188]}
   );
   gpc615_5 gpc444 (
      {stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_10[319]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[75],stage1_11[100],stage1_10[135],stage1_9[189]}
   );
   gpc615_5 gpc445 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_10[320]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[76],stage1_11[101],stage1_10[136],stage1_9[190]}
   );
   gpc615_5 gpc446 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295]},
      {stage0_10[321]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[77],stage1_11[102],stage1_10[137],stage1_9[191]}
   );
   gpc615_5 gpc447 (
      {stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_10[322]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[78],stage1_11[103],stage1_10[138],stage1_9[192]}
   );
   gpc615_5 gpc448 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_10[323]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[79],stage1_11[104],stage1_10[139],stage1_9[193]}
   );
   gpc615_5 gpc449 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310]},
      {stage0_10[324]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[80],stage1_11[105],stage1_10[140],stage1_9[194]}
   );
   gpc615_5 gpc450 (
      {stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_10[325]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[81],stage1_11[106],stage1_10[141],stage1_9[195]}
   );
   gpc615_5 gpc451 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_10[326]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[82],stage1_11[107],stage1_10[142],stage1_9[196]}
   );
   gpc615_5 gpc452 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325]},
      {stage0_10[327]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[83],stage1_11[108],stage1_10[143],stage1_9[197]}
   );
   gpc615_5 gpc453 (
      {stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_10[328]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[84],stage1_11[109],stage1_10[144],stage1_9[198]}
   );
   gpc615_5 gpc454 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_10[329]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[85],stage1_11[110],stage1_10[145],stage1_9[199]}
   );
   gpc615_5 gpc455 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340]},
      {stage0_10[330]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[86],stage1_11[111],stage1_10[146],stage1_9[200]}
   );
   gpc615_5 gpc456 (
      {stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_10[331]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[87],stage1_11[112],stage1_10[147],stage1_9[201]}
   );
   gpc615_5 gpc457 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_10[332]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[88],stage1_11[113],stage1_10[148],stage1_9[202]}
   );
   gpc615_5 gpc458 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355]},
      {stage0_10[333]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[89],stage1_11[114],stage1_10[149],stage1_9[203]}
   );
   gpc615_5 gpc459 (
      {stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_10[334]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[90],stage1_11[115],stage1_10[150],stage1_9[204]}
   );
   gpc615_5 gpc460 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_10[335]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[91],stage1_11[116],stage1_10[151],stage1_9[205]}
   );
   gpc615_5 gpc461 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370]},
      {stage0_10[336]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[92],stage1_11[117],stage1_10[152],stage1_9[206]}
   );
   gpc615_5 gpc462 (
      {stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_10[337]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[93],stage1_11[118],stage1_10[153],stage1_9[207]}
   );
   gpc615_5 gpc463 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_10[338]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[94],stage1_11[119],stage1_10[154],stage1_9[208]}
   );
   gpc615_5 gpc464 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385]},
      {stage0_10[339]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[95],stage1_11[120],stage1_10[155],stage1_9[209]}
   );
   gpc615_5 gpc465 (
      {stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_10[340]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[96],stage1_11[121],stage1_10[156],stage1_9[210]}
   );
   gpc615_5 gpc466 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_10[341]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[97],stage1_11[122],stage1_10[157],stage1_9[211]}
   );
   gpc615_5 gpc467 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400]},
      {stage0_10[342]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[98],stage1_11[123],stage1_10[158],stage1_9[212]}
   );
   gpc615_5 gpc468 (
      {stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_10[343]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[99],stage1_11[124],stage1_10[159],stage1_9[213]}
   );
   gpc615_5 gpc469 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410]},
      {stage0_10[344]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[100],stage1_11[125],stage1_10[160],stage1_9[214]}
   );
   gpc615_5 gpc470 (
      {stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415]},
      {stage0_10[345]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[101],stage1_11[126],stage1_10[161],stage1_9[215]}
   );
   gpc615_5 gpc471 (
      {stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_10[346]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[102],stage1_11[127],stage1_10[162],stage1_9[216]}
   );
   gpc615_5 gpc472 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[347]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[103],stage1_11[128],stage1_10[163],stage1_9[217]}
   );
   gpc615_5 gpc473 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[348]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[104],stage1_11[129],stage1_10[164],stage1_9[218]}
   );
   gpc615_5 gpc474 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[349]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[105],stage1_11[130],stage1_10[165],stage1_9[219]}
   );
   gpc615_5 gpc475 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[350]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[106],stage1_11[131],stage1_10[166],stage1_9[220]}
   );
   gpc615_5 gpc476 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[351]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[107],stage1_11[132],stage1_10[167],stage1_9[221]}
   );
   gpc615_5 gpc477 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[352]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[108],stage1_11[133],stage1_10[168],stage1_9[222]}
   );
   gpc615_5 gpc478 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[353]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[109],stage1_11[134],stage1_10[169],stage1_9[223]}
   );
   gpc615_5 gpc479 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[354]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[110],stage1_11[135],stage1_10[170],stage1_9[224]}
   );
   gpc615_5 gpc480 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[355]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[111],stage1_11[136],stage1_10[171],stage1_9[225]}
   );
   gpc615_5 gpc481 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[356]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[112],stage1_11[137],stage1_10[172],stage1_9[226]}
   );
   gpc615_5 gpc482 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[357]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[113],stage1_11[138],stage1_10[173],stage1_9[227]}
   );
   gpc606_5 gpc483 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[65],stage1_12[114],stage1_11[139],stage1_10[174]}
   );
   gpc606_5 gpc484 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[66],stage1_12[115],stage1_11[140],stage1_10[175]}
   );
   gpc606_5 gpc485 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[67],stage1_12[116],stage1_11[141],stage1_10[176]}
   );
   gpc606_5 gpc486 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[68],stage1_12[117],stage1_11[142],stage1_10[177]}
   );
   gpc606_5 gpc487 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[69],stage1_12[118],stage1_11[143],stage1_10[178]}
   );
   gpc606_5 gpc488 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[70],stage1_12[119],stage1_11[144],stage1_10[179]}
   );
   gpc615_5 gpc489 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[71],stage1_12[120],stage1_11[145],stage1_10[180]}
   );
   gpc615_5 gpc490 (
      {stage0_10[399], stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[72],stage1_12[121],stage1_11[146],stage1_10[181]}
   );
   gpc615_5 gpc491 (
      {stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[73],stage1_12[122],stage1_11[147],stage1_10[182]}
   );
   gpc615_5 gpc492 (
      {stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[74],stage1_12[123],stage1_11[148],stage1_10[183]}
   );
   gpc615_5 gpc493 (
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[75],stage1_12[124],stage1_11[149],stage1_10[184]}
   );
   gpc615_5 gpc494 (
      {stage0_10[419], stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[76],stage1_12[125],stage1_11[150],stage1_10[185]}
   );
   gpc615_5 gpc495 (
      {stage0_10[424], stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[77],stage1_12[126],stage1_11[151],stage1_10[186]}
   );
   gpc615_5 gpc496 (
      {stage0_10[429], stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[78],stage1_12[127],stage1_11[152],stage1_10[187]}
   );
   gpc615_5 gpc497 (
      {stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[79],stage1_12[128],stage1_11[153],stage1_10[188]}
   );
   gpc615_5 gpc498 (
      {stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[80],stage1_12[129],stage1_11[154],stage1_10[189]}
   );
   gpc615_5 gpc499 (
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448]},
      {stage0_11[400]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[81],stage1_12[130],stage1_11[155],stage1_10[190]}
   );
   gpc615_5 gpc500 (
      {stage0_10[449], stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453]},
      {stage0_11[401]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[82],stage1_12[131],stage1_11[156],stage1_10[191]}
   );
   gpc615_5 gpc501 (
      {stage0_10[454], stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458]},
      {stage0_11[402]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[83],stage1_12[132],stage1_11[157],stage1_10[192]}
   );
   gpc615_5 gpc502 (
      {stage0_10[459], stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463]},
      {stage0_11[403]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[84],stage1_12[133],stage1_11[158],stage1_10[193]}
   );
   gpc615_5 gpc503 (
      {stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468]},
      {stage0_11[404]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[85],stage1_12[134],stage1_11[159],stage1_10[194]}
   );
   gpc615_5 gpc504 (
      {stage0_10[469], stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473]},
      {stage0_11[405]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[86],stage1_12[135],stage1_11[160],stage1_10[195]}
   );
   gpc615_5 gpc505 (
      {stage0_10[474], stage0_10[475], stage0_10[476], stage0_10[477], stage0_10[478]},
      {stage0_11[406]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[87],stage1_12[136],stage1_11[161],stage1_10[196]}
   );
   gpc615_5 gpc506 (
      {stage0_10[479], stage0_10[480], stage0_10[481], stage0_10[482], stage0_10[483]},
      {stage0_11[407]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[88],stage1_12[137],stage1_11[162],stage1_10[197]}
   );
   gpc615_5 gpc507 (
      {stage0_10[484], stage0_10[485], stage0_10[486], stage0_10[487], stage0_10[488]},
      {stage0_11[408]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[89],stage1_12[138],stage1_11[163],stage1_10[198]}
   );
   gpc615_5 gpc508 (
      {stage0_10[489], stage0_10[490], stage0_10[491], stage0_10[492], stage0_10[493]},
      {stage0_11[409]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[90],stage1_12[139],stage1_11[164],stage1_10[199]}
   );
   gpc615_5 gpc509 (
      {stage0_10[494], stage0_10[495], stage0_10[496], stage0_10[497], stage0_10[498]},
      {stage0_11[410]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[91],stage1_12[140],stage1_11[165],stage1_10[200]}
   );
   gpc615_5 gpc510 (
      {stage0_10[499], stage0_10[500], stage0_10[501], stage0_10[502], stage0_10[503]},
      {stage0_11[411]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[92],stage1_12[141],stage1_11[166],stage1_10[201]}
   );
   gpc606_5 gpc511 (
      {stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[28],stage1_13[93],stage1_12[142],stage1_11[167]}
   );
   gpc606_5 gpc512 (
      {stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[29],stage1_13[94],stage1_12[143],stage1_11[168]}
   );
   gpc606_5 gpc513 (
      {stage0_11[424], stage0_11[425], stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[30],stage1_13[95],stage1_12[144],stage1_11[169]}
   );
   gpc606_5 gpc514 (
      {stage0_11[430], stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[31],stage1_13[96],stage1_12[145],stage1_11[170]}
   );
   gpc606_5 gpc515 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[32],stage1_13[97],stage1_12[146],stage1_11[171]}
   );
   gpc606_5 gpc516 (
      {stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[33],stage1_13[98],stage1_12[147],stage1_11[172]}
   );
   gpc606_5 gpc517 (
      {stage0_11[448], stage0_11[449], stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[34],stage1_13[99],stage1_12[148],stage1_11[173]}
   );
   gpc606_5 gpc518 (
      {stage0_11[454], stage0_11[455], stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[35],stage1_13[100],stage1_12[149],stage1_11[174]}
   );
   gpc606_5 gpc519 (
      {stage0_11[460], stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[36],stage1_13[101],stage1_12[150],stage1_11[175]}
   );
   gpc615_5 gpc520 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[168]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[37],stage1_13[102],stage1_12[151],stage1_11[176]}
   );
   gpc615_5 gpc521 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[169]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[38],stage1_13[103],stage1_12[152],stage1_11[177]}
   );
   gpc615_5 gpc522 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[170]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[39],stage1_13[104],stage1_12[153],stage1_11[178]}
   );
   gpc615_5 gpc523 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[171]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[40],stage1_13[105],stage1_12[154],stage1_11[179]}
   );
   gpc615_5 gpc524 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[172]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[41],stage1_13[106],stage1_12[155],stage1_11[180]}
   );
   gpc615_5 gpc525 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[173]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[42],stage1_13[107],stage1_12[156],stage1_11[181]}
   );
   gpc615_5 gpc526 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[174]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[43],stage1_13[108],stage1_12[157],stage1_11[182]}
   );
   gpc615_5 gpc527 (
      {stage0_11[501], stage0_11[502], stage0_11[503], stage0_11[504], stage0_11[505]},
      {stage0_12[175]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[44],stage1_13[109],stage1_12[158],stage1_11[183]}
   );
   gpc606_5 gpc528 (
      {stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[17],stage1_14[45],stage1_13[110],stage1_12[159]}
   );
   gpc606_5 gpc529 (
      {stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[18],stage1_14[46],stage1_13[111],stage1_12[160]}
   );
   gpc606_5 gpc530 (
      {stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[19],stage1_14[47],stage1_13[112],stage1_12[161]}
   );
   gpc606_5 gpc531 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[20],stage1_14[48],stage1_13[113],stage1_12[162]}
   );
   gpc606_5 gpc532 (
      {stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[21],stage1_14[49],stage1_13[114],stage1_12[163]}
   );
   gpc606_5 gpc533 (
      {stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[22],stage1_14[50],stage1_13[115],stage1_12[164]}
   );
   gpc606_5 gpc534 (
      {stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[23],stage1_14[51],stage1_13[116],stage1_12[165]}
   );
   gpc606_5 gpc535 (
      {stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[24],stage1_14[52],stage1_13[117],stage1_12[166]}
   );
   gpc606_5 gpc536 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[25],stage1_14[53],stage1_13[118],stage1_12[167]}
   );
   gpc606_5 gpc537 (
      {stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[26],stage1_14[54],stage1_13[119],stage1_12[168]}
   );
   gpc606_5 gpc538 (
      {stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[27],stage1_14[55],stage1_13[120],stage1_12[169]}
   );
   gpc606_5 gpc539 (
      {stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[28],stage1_14[56],stage1_13[121],stage1_12[170]}
   );
   gpc606_5 gpc540 (
      {stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[29],stage1_14[57],stage1_13[122],stage1_12[171]}
   );
   gpc606_5 gpc541 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[30],stage1_14[58],stage1_13[123],stage1_12[172]}
   );
   gpc606_5 gpc542 (
      {stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[31],stage1_14[59],stage1_13[124],stage1_12[173]}
   );
   gpc606_5 gpc543 (
      {stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[32],stage1_14[60],stage1_13[125],stage1_12[174]}
   );
   gpc606_5 gpc544 (
      {stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[33],stage1_14[61],stage1_13[126],stage1_12[175]}
   );
   gpc606_5 gpc545 (
      {stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[34],stage1_14[62],stage1_13[127],stage1_12[176]}
   );
   gpc606_5 gpc546 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[35],stage1_14[63],stage1_13[128],stage1_12[177]}
   );
   gpc606_5 gpc547 (
      {stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[36],stage1_14[64],stage1_13[129],stage1_12[178]}
   );
   gpc606_5 gpc548 (
      {stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[37],stage1_14[65],stage1_13[130],stage1_12[179]}
   );
   gpc615_5 gpc549 (
      {stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306]},
      {stage0_13[102]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[38],stage1_14[66],stage1_13[131],stage1_12[180]}
   );
   gpc615_5 gpc550 (
      {stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_13[103]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[39],stage1_14[67],stage1_13[132],stage1_12[181]}
   );
   gpc615_5 gpc551 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_13[104]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[40],stage1_14[68],stage1_13[133],stage1_12[182]}
   );
   gpc615_5 gpc552 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[105]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[41],stage1_14[69],stage1_13[134],stage1_12[183]}
   );
   gpc615_5 gpc553 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[106]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[42],stage1_14[70],stage1_13[135],stage1_12[184]}
   );
   gpc615_5 gpc554 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[107]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[43],stage1_14[71],stage1_13[136],stage1_12[185]}
   );
   gpc615_5 gpc555 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[108]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[44],stage1_14[72],stage1_13[137],stage1_12[186]}
   );
   gpc615_5 gpc556 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[109]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[45],stage1_14[73],stage1_13[138],stage1_12[187]}
   );
   gpc615_5 gpc557 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[110]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[46],stage1_14[74],stage1_13[139],stage1_12[188]}
   );
   gpc615_5 gpc558 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[111]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[47],stage1_14[75],stage1_13[140],stage1_12[189]}
   );
   gpc615_5 gpc559 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[112]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[48],stage1_14[76],stage1_13[141],stage1_12[190]}
   );
   gpc615_5 gpc560 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[113]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[49],stage1_14[77],stage1_13[142],stage1_12[191]}
   );
   gpc615_5 gpc561 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[114]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[50],stage1_14[78],stage1_13[143],stage1_12[192]}
   );
   gpc615_5 gpc562 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[115]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[51],stage1_14[79],stage1_13[144],stage1_12[193]}
   );
   gpc615_5 gpc563 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[116]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[52],stage1_14[80],stage1_13[145],stage1_12[194]}
   );
   gpc615_5 gpc564 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[117]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[53],stage1_14[81],stage1_13[146],stage1_12[195]}
   );
   gpc615_5 gpc565 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[118]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[54],stage1_14[82],stage1_13[147],stage1_12[196]}
   );
   gpc615_5 gpc566 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[119]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[55],stage1_14[83],stage1_13[148],stage1_12[197]}
   );
   gpc615_5 gpc567 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[120]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[56],stage1_14[84],stage1_13[149],stage1_12[198]}
   );
   gpc615_5 gpc568 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[121]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[57],stage1_14[85],stage1_13[150],stage1_12[199]}
   );
   gpc615_5 gpc569 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[122]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[58],stage1_14[86],stage1_13[151],stage1_12[200]}
   );
   gpc615_5 gpc570 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[123]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[59],stage1_14[87],stage1_13[152],stage1_12[201]}
   );
   gpc615_5 gpc571 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[124]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[60],stage1_14[88],stage1_13[153],stage1_12[202]}
   );
   gpc615_5 gpc572 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[125]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[61],stage1_14[89],stage1_13[154],stage1_12[203]}
   );
   gpc615_5 gpc573 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[126]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[62],stage1_14[90],stage1_13[155],stage1_12[204]}
   );
   gpc615_5 gpc574 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[127]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[63],stage1_14[91],stage1_13[156],stage1_12[205]}
   );
   gpc615_5 gpc575 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[128]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[64],stage1_14[92],stage1_13[157],stage1_12[206]}
   );
   gpc615_5 gpc576 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[129]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[65],stage1_14[93],stage1_13[158],stage1_12[207]}
   );
   gpc615_5 gpc577 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[130]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[66],stage1_14[94],stage1_13[159],stage1_12[208]}
   );
   gpc615_5 gpc578 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[131]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[67],stage1_14[95],stage1_13[160],stage1_12[209]}
   );
   gpc615_5 gpc579 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[132]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[68],stage1_14[96],stage1_13[161],stage1_12[210]}
   );
   gpc615_5 gpc580 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[133]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[69],stage1_14[97],stage1_13[162],stage1_12[211]}
   );
   gpc615_5 gpc581 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[134]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[70],stage1_14[98],stage1_13[163],stage1_12[212]}
   );
   gpc615_5 gpc582 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[135]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[71],stage1_14[99],stage1_13[164],stage1_12[213]}
   );
   gpc615_5 gpc583 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[136]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[72],stage1_14[100],stage1_13[165],stage1_12[214]}
   );
   gpc615_5 gpc584 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[137]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[73],stage1_14[101],stage1_13[166],stage1_12[215]}
   );
   gpc615_5 gpc585 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[138]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[74],stage1_14[102],stage1_13[167],stage1_12[216]}
   );
   gpc615_5 gpc586 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[139]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[75],stage1_14[103],stage1_13[168],stage1_12[217]}
   );
   gpc615_5 gpc587 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[140]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[76],stage1_14[104],stage1_13[169],stage1_12[218]}
   );
   gpc615_5 gpc588 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[141]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[77],stage1_14[105],stage1_13[170],stage1_12[219]}
   );
   gpc615_5 gpc589 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[142]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[78],stage1_14[106],stage1_13[171],stage1_12[220]}
   );
   gpc615_5 gpc590 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[143]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[79],stage1_14[107],stage1_13[172],stage1_12[221]}
   );
   gpc606_5 gpc591 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[63],stage1_15[80],stage1_14[108],stage1_13[173]}
   );
   gpc606_5 gpc592 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[64],stage1_15[81],stage1_14[109],stage1_13[174]}
   );
   gpc606_5 gpc593 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[65],stage1_15[82],stage1_14[110],stage1_13[175]}
   );
   gpc615_5 gpc594 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166]},
      {stage0_14[378]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[66],stage1_15[83],stage1_14[111],stage1_13[176]}
   );
   gpc615_5 gpc595 (
      {stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_14[379]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[67],stage1_15[84],stage1_14[112],stage1_13[177]}
   );
   gpc615_5 gpc596 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_14[380]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[68],stage1_15[85],stage1_14[113],stage1_13[178]}
   );
   gpc615_5 gpc597 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181]},
      {stage0_14[381]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[69],stage1_15[86],stage1_14[114],stage1_13[179]}
   );
   gpc615_5 gpc598 (
      {stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186]},
      {stage0_14[382]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[70],stage1_15[87],stage1_14[115],stage1_13[180]}
   );
   gpc615_5 gpc599 (
      {stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_14[383]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[71],stage1_15[88],stage1_14[116],stage1_13[181]}
   );
   gpc615_5 gpc600 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196]},
      {stage0_14[384]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[72],stage1_15[89],stage1_14[117],stage1_13[182]}
   );
   gpc615_5 gpc601 (
      {stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_14[385]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[73],stage1_15[90],stage1_14[118],stage1_13[183]}
   );
   gpc615_5 gpc602 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_14[386]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[74],stage1_15[91],stage1_14[119],stage1_13[184]}
   );
   gpc615_5 gpc603 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211]},
      {stage0_14[387]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[75],stage1_15[92],stage1_14[120],stage1_13[185]}
   );
   gpc615_5 gpc604 (
      {stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216]},
      {stage0_14[388]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[76],stage1_15[93],stage1_14[121],stage1_13[186]}
   );
   gpc615_5 gpc605 (
      {stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_14[389]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[77],stage1_15[94],stage1_14[122],stage1_13[187]}
   );
   gpc615_5 gpc606 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226]},
      {stage0_14[390]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[78],stage1_15[95],stage1_14[123],stage1_13[188]}
   );
   gpc615_5 gpc607 (
      {stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231]},
      {stage0_14[391]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[79],stage1_15[96],stage1_14[124],stage1_13[189]}
   );
   gpc615_5 gpc608 (
      {stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_14[392]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[80],stage1_15[97],stage1_14[125],stage1_13[190]}
   );
   gpc615_5 gpc609 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241]},
      {stage0_14[393]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[81],stage1_15[98],stage1_14[126],stage1_13[191]}
   );
   gpc615_5 gpc610 (
      {stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246]},
      {stage0_14[394]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[82],stage1_15[99],stage1_14[127],stage1_13[192]}
   );
   gpc615_5 gpc611 (
      {stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_14[395]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[83],stage1_15[100],stage1_14[128],stage1_13[193]}
   );
   gpc615_5 gpc612 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256]},
      {stage0_14[396]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[84],stage1_15[101],stage1_14[129],stage1_13[194]}
   );
   gpc615_5 gpc613 (
      {stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261]},
      {stage0_14[397]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[85],stage1_15[102],stage1_14[130],stage1_13[195]}
   );
   gpc615_5 gpc614 (
      {stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_14[398]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[86],stage1_15[103],stage1_14[131],stage1_13[196]}
   );
   gpc615_5 gpc615 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271]},
      {stage0_14[399]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[87],stage1_15[104],stage1_14[132],stage1_13[197]}
   );
   gpc615_5 gpc616 (
      {stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276]},
      {stage0_14[400]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[88],stage1_15[105],stage1_14[133],stage1_13[198]}
   );
   gpc615_5 gpc617 (
      {stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_14[401]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[89],stage1_15[106],stage1_14[134],stage1_13[199]}
   );
   gpc615_5 gpc618 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286]},
      {stage0_14[402]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[90],stage1_15[107],stage1_14[135],stage1_13[200]}
   );
   gpc615_5 gpc619 (
      {stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291]},
      {stage0_14[403]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[91],stage1_15[108],stage1_14[136],stage1_13[201]}
   );
   gpc615_5 gpc620 (
      {stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_14[404]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[92],stage1_15[109],stage1_14[137],stage1_13[202]}
   );
   gpc615_5 gpc621 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301]},
      {stage0_14[405]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[93],stage1_15[110],stage1_14[138],stage1_13[203]}
   );
   gpc615_5 gpc622 (
      {stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306]},
      {stage0_14[406]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[94],stage1_15[111],stage1_14[139],stage1_13[204]}
   );
   gpc615_5 gpc623 (
      {stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_14[407]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[95],stage1_15[112],stage1_14[140],stage1_13[205]}
   );
   gpc615_5 gpc624 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316]},
      {stage0_14[408]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[96],stage1_15[113],stage1_14[141],stage1_13[206]}
   );
   gpc615_5 gpc625 (
      {stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321]},
      {stage0_14[409]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[97],stage1_15[114],stage1_14[142],stage1_13[207]}
   );
   gpc615_5 gpc626 (
      {stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_14[410]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[98],stage1_15[115],stage1_14[143],stage1_13[208]}
   );
   gpc615_5 gpc627 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331]},
      {stage0_14[411]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[99],stage1_15[116],stage1_14[144],stage1_13[209]}
   );
   gpc615_5 gpc628 (
      {stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336]},
      {stage0_14[412]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[100],stage1_15[117],stage1_14[145],stage1_13[210]}
   );
   gpc615_5 gpc629 (
      {stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_14[413]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[101],stage1_15[118],stage1_14[146],stage1_13[211]}
   );
   gpc615_5 gpc630 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346]},
      {stage0_14[414]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[102],stage1_15[119],stage1_14[147],stage1_13[212]}
   );
   gpc615_5 gpc631 (
      {stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351]},
      {stage0_14[415]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[103],stage1_15[120],stage1_14[148],stage1_13[213]}
   );
   gpc615_5 gpc632 (
      {stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_14[416]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[104],stage1_15[121],stage1_14[149],stage1_13[214]}
   );
   gpc615_5 gpc633 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361]},
      {stage0_14[417]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[105],stage1_15[122],stage1_14[150],stage1_13[215]}
   );
   gpc615_5 gpc634 (
      {stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366]},
      {stage0_14[418]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[106],stage1_15[123],stage1_14[151],stage1_13[216]}
   );
   gpc615_5 gpc635 (
      {stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_14[419]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[107],stage1_15[124],stage1_14[152],stage1_13[217]}
   );
   gpc615_5 gpc636 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376]},
      {stage0_14[420]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[108],stage1_15[125],stage1_14[153],stage1_13[218]}
   );
   gpc615_5 gpc637 (
      {stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381]},
      {stage0_14[421]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[109],stage1_15[126],stage1_14[154],stage1_13[219]}
   );
   gpc615_5 gpc638 (
      {stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_14[422]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[110],stage1_15[127],stage1_14[155],stage1_13[220]}
   );
   gpc615_5 gpc639 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391]},
      {stage0_14[423]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[111],stage1_15[128],stage1_14[156],stage1_13[221]}
   );
   gpc615_5 gpc640 (
      {stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396]},
      {stage0_14[424]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[112],stage1_15[129],stage1_14[157],stage1_13[222]}
   );
   gpc615_5 gpc641 (
      {stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_14[425]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[113],stage1_15[130],stage1_14[158],stage1_13[223]}
   );
   gpc615_5 gpc642 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406]},
      {stage0_14[426]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[114],stage1_15[131],stage1_14[159],stage1_13[224]}
   );
   gpc615_5 gpc643 (
      {stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411]},
      {stage0_14[427]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[115],stage1_15[132],stage1_14[160],stage1_13[225]}
   );
   gpc615_5 gpc644 (
      {stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_14[428]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[116],stage1_15[133],stage1_14[161],stage1_13[226]}
   );
   gpc615_5 gpc645 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421]},
      {stage0_14[429]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[117],stage1_15[134],stage1_14[162],stage1_13[227]}
   );
   gpc615_5 gpc646 (
      {stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426]},
      {stage0_14[430]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[118],stage1_15[135],stage1_14[163],stage1_13[228]}
   );
   gpc615_5 gpc647 (
      {stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_14[431]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[119],stage1_15[136],stage1_14[164],stage1_13[229]}
   );
   gpc615_5 gpc648 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436]},
      {stage0_14[432]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[120],stage1_15[137],stage1_14[165],stage1_13[230]}
   );
   gpc615_5 gpc649 (
      {stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441]},
      {stage0_14[433]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[121],stage1_15[138],stage1_14[166],stage1_13[231]}
   );
   gpc615_5 gpc650 (
      {stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_14[434]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[122],stage1_15[139],stage1_14[167],stage1_13[232]}
   );
   gpc615_5 gpc651 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451]},
      {stage0_14[435]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[123],stage1_15[140],stage1_14[168],stage1_13[233]}
   );
   gpc615_5 gpc652 (
      {stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456]},
      {stage0_14[436]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[124],stage1_15[141],stage1_14[169],stage1_13[234]}
   );
   gpc615_5 gpc653 (
      {stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_14[437]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[125],stage1_15[142],stage1_14[170],stage1_13[235]}
   );
   gpc615_5 gpc654 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466]},
      {stage0_14[438]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[126],stage1_15[143],stage1_14[171],stage1_13[236]}
   );
   gpc1_1 gpc655 (
      {stage0_0[509]},
      {stage1_0[98]}
   );
   gpc1_1 gpc656 (
      {stage0_0[510]},
      {stage1_0[99]}
   );
   gpc1_1 gpc657 (
      {stage0_0[511]},
      {stage1_0[100]}
   );
   gpc1_1 gpc658 (
      {stage0_1[476]},
      {stage1_1[144]}
   );
   gpc1_1 gpc659 (
      {stage0_1[477]},
      {stage1_1[145]}
   );
   gpc1_1 gpc660 (
      {stage0_1[478]},
      {stage1_1[146]}
   );
   gpc1_1 gpc661 (
      {stage0_1[479]},
      {stage1_1[147]}
   );
   gpc1_1 gpc662 (
      {stage0_1[480]},
      {stage1_1[148]}
   );
   gpc1_1 gpc663 (
      {stage0_1[481]},
      {stage1_1[149]}
   );
   gpc1_1 gpc664 (
      {stage0_1[482]},
      {stage1_1[150]}
   );
   gpc1_1 gpc665 (
      {stage0_1[483]},
      {stage1_1[151]}
   );
   gpc1_1 gpc666 (
      {stage0_1[484]},
      {stage1_1[152]}
   );
   gpc1_1 gpc667 (
      {stage0_1[485]},
      {stage1_1[153]}
   );
   gpc1_1 gpc668 (
      {stage0_1[486]},
      {stage1_1[154]}
   );
   gpc1_1 gpc669 (
      {stage0_1[487]},
      {stage1_1[155]}
   );
   gpc1_1 gpc670 (
      {stage0_1[488]},
      {stage1_1[156]}
   );
   gpc1_1 gpc671 (
      {stage0_1[489]},
      {stage1_1[157]}
   );
   gpc1_1 gpc672 (
      {stage0_1[490]},
      {stage1_1[158]}
   );
   gpc1_1 gpc673 (
      {stage0_1[491]},
      {stage1_1[159]}
   );
   gpc1_1 gpc674 (
      {stage0_1[492]},
      {stage1_1[160]}
   );
   gpc1_1 gpc675 (
      {stage0_1[493]},
      {stage1_1[161]}
   );
   gpc1_1 gpc676 (
      {stage0_1[494]},
      {stage1_1[162]}
   );
   gpc1_1 gpc677 (
      {stage0_1[495]},
      {stage1_1[163]}
   );
   gpc1_1 gpc678 (
      {stage0_1[496]},
      {stage1_1[164]}
   );
   gpc1_1 gpc679 (
      {stage0_1[497]},
      {stage1_1[165]}
   );
   gpc1_1 gpc680 (
      {stage0_1[498]},
      {stage1_1[166]}
   );
   gpc1_1 gpc681 (
      {stage0_1[499]},
      {stage1_1[167]}
   );
   gpc1_1 gpc682 (
      {stage0_1[500]},
      {stage1_1[168]}
   );
   gpc1_1 gpc683 (
      {stage0_1[501]},
      {stage1_1[169]}
   );
   gpc1_1 gpc684 (
      {stage0_1[502]},
      {stage1_1[170]}
   );
   gpc1_1 gpc685 (
      {stage0_1[503]},
      {stage1_1[171]}
   );
   gpc1_1 gpc686 (
      {stage0_1[504]},
      {stage1_1[172]}
   );
   gpc1_1 gpc687 (
      {stage0_1[505]},
      {stage1_1[173]}
   );
   gpc1_1 gpc688 (
      {stage0_1[506]},
      {stage1_1[174]}
   );
   gpc1_1 gpc689 (
      {stage0_1[507]},
      {stage1_1[175]}
   );
   gpc1_1 gpc690 (
      {stage0_1[508]},
      {stage1_1[176]}
   );
   gpc1_1 gpc691 (
      {stage0_1[509]},
      {stage1_1[177]}
   );
   gpc1_1 gpc692 (
      {stage0_1[510]},
      {stage1_1[178]}
   );
   gpc1_1 gpc693 (
      {stage0_1[511]},
      {stage1_1[179]}
   );
   gpc1_1 gpc694 (
      {stage0_3[466]},
      {stage1_3[200]}
   );
   gpc1_1 gpc695 (
      {stage0_3[467]},
      {stage1_3[201]}
   );
   gpc1_1 gpc696 (
      {stage0_3[468]},
      {stage1_3[202]}
   );
   gpc1_1 gpc697 (
      {stage0_3[469]},
      {stage1_3[203]}
   );
   gpc1_1 gpc698 (
      {stage0_3[470]},
      {stage1_3[204]}
   );
   gpc1_1 gpc699 (
      {stage0_3[471]},
      {stage1_3[205]}
   );
   gpc1_1 gpc700 (
      {stage0_3[472]},
      {stage1_3[206]}
   );
   gpc1_1 gpc701 (
      {stage0_3[473]},
      {stage1_3[207]}
   );
   gpc1_1 gpc702 (
      {stage0_3[474]},
      {stage1_3[208]}
   );
   gpc1_1 gpc703 (
      {stage0_3[475]},
      {stage1_3[209]}
   );
   gpc1_1 gpc704 (
      {stage0_3[476]},
      {stage1_3[210]}
   );
   gpc1_1 gpc705 (
      {stage0_3[477]},
      {stage1_3[211]}
   );
   gpc1_1 gpc706 (
      {stage0_3[478]},
      {stage1_3[212]}
   );
   gpc1_1 gpc707 (
      {stage0_3[479]},
      {stage1_3[213]}
   );
   gpc1_1 gpc708 (
      {stage0_3[480]},
      {stage1_3[214]}
   );
   gpc1_1 gpc709 (
      {stage0_3[481]},
      {stage1_3[215]}
   );
   gpc1_1 gpc710 (
      {stage0_3[482]},
      {stage1_3[216]}
   );
   gpc1_1 gpc711 (
      {stage0_3[483]},
      {stage1_3[217]}
   );
   gpc1_1 gpc712 (
      {stage0_3[484]},
      {stage1_3[218]}
   );
   gpc1_1 gpc713 (
      {stage0_3[485]},
      {stage1_3[219]}
   );
   gpc1_1 gpc714 (
      {stage0_3[486]},
      {stage1_3[220]}
   );
   gpc1_1 gpc715 (
      {stage0_3[487]},
      {stage1_3[221]}
   );
   gpc1_1 gpc716 (
      {stage0_3[488]},
      {stage1_3[222]}
   );
   gpc1_1 gpc717 (
      {stage0_3[489]},
      {stage1_3[223]}
   );
   gpc1_1 gpc718 (
      {stage0_3[490]},
      {stage1_3[224]}
   );
   gpc1_1 gpc719 (
      {stage0_3[491]},
      {stage1_3[225]}
   );
   gpc1_1 gpc720 (
      {stage0_3[492]},
      {stage1_3[226]}
   );
   gpc1_1 gpc721 (
      {stage0_3[493]},
      {stage1_3[227]}
   );
   gpc1_1 gpc722 (
      {stage0_3[494]},
      {stage1_3[228]}
   );
   gpc1_1 gpc723 (
      {stage0_3[495]},
      {stage1_3[229]}
   );
   gpc1_1 gpc724 (
      {stage0_3[496]},
      {stage1_3[230]}
   );
   gpc1_1 gpc725 (
      {stage0_3[497]},
      {stage1_3[231]}
   );
   gpc1_1 gpc726 (
      {stage0_3[498]},
      {stage1_3[232]}
   );
   gpc1_1 gpc727 (
      {stage0_3[499]},
      {stage1_3[233]}
   );
   gpc1_1 gpc728 (
      {stage0_3[500]},
      {stage1_3[234]}
   );
   gpc1_1 gpc729 (
      {stage0_3[501]},
      {stage1_3[235]}
   );
   gpc1_1 gpc730 (
      {stage0_3[502]},
      {stage1_3[236]}
   );
   gpc1_1 gpc731 (
      {stage0_3[503]},
      {stage1_3[237]}
   );
   gpc1_1 gpc732 (
      {stage0_3[504]},
      {stage1_3[238]}
   );
   gpc1_1 gpc733 (
      {stage0_3[505]},
      {stage1_3[239]}
   );
   gpc1_1 gpc734 (
      {stage0_3[506]},
      {stage1_3[240]}
   );
   gpc1_1 gpc735 (
      {stage0_3[507]},
      {stage1_3[241]}
   );
   gpc1_1 gpc736 (
      {stage0_3[508]},
      {stage1_3[242]}
   );
   gpc1_1 gpc737 (
      {stage0_3[509]},
      {stage1_3[243]}
   );
   gpc1_1 gpc738 (
      {stage0_3[510]},
      {stage1_3[244]}
   );
   gpc1_1 gpc739 (
      {stage0_3[511]},
      {stage1_3[245]}
   );
   gpc1_1 gpc740 (
      {stage0_5[505]},
      {stage1_5[211]}
   );
   gpc1_1 gpc741 (
      {stage0_5[506]},
      {stage1_5[212]}
   );
   gpc1_1 gpc742 (
      {stage0_5[507]},
      {stage1_5[213]}
   );
   gpc1_1 gpc743 (
      {stage0_5[508]},
      {stage1_5[214]}
   );
   gpc1_1 gpc744 (
      {stage0_5[509]},
      {stage1_5[215]}
   );
   gpc1_1 gpc745 (
      {stage0_5[510]},
      {stage1_5[216]}
   );
   gpc1_1 gpc746 (
      {stage0_5[511]},
      {stage1_5[217]}
   );
   gpc1_1 gpc747 (
      {stage0_6[505]},
      {stage1_6[200]}
   );
   gpc1_1 gpc748 (
      {stage0_6[506]},
      {stage1_6[201]}
   );
   gpc1_1 gpc749 (
      {stage0_6[507]},
      {stage1_6[202]}
   );
   gpc1_1 gpc750 (
      {stage0_6[508]},
      {stage1_6[203]}
   );
   gpc1_1 gpc751 (
      {stage0_6[509]},
      {stage1_6[204]}
   );
   gpc1_1 gpc752 (
      {stage0_6[510]},
      {stage1_6[205]}
   );
   gpc1_1 gpc753 (
      {stage0_6[511]},
      {stage1_6[206]}
   );
   gpc1_1 gpc754 (
      {stage0_7[501]},
      {stage1_7[196]}
   );
   gpc1_1 gpc755 (
      {stage0_7[502]},
      {stage1_7[197]}
   );
   gpc1_1 gpc756 (
      {stage0_7[503]},
      {stage1_7[198]}
   );
   gpc1_1 gpc757 (
      {stage0_7[504]},
      {stage1_7[199]}
   );
   gpc1_1 gpc758 (
      {stage0_7[505]},
      {stage1_7[200]}
   );
   gpc1_1 gpc759 (
      {stage0_7[506]},
      {stage1_7[201]}
   );
   gpc1_1 gpc760 (
      {stage0_7[507]},
      {stage1_7[202]}
   );
   gpc1_1 gpc761 (
      {stage0_7[508]},
      {stage1_7[203]}
   );
   gpc1_1 gpc762 (
      {stage0_7[509]},
      {stage1_7[204]}
   );
   gpc1_1 gpc763 (
      {stage0_7[510]},
      {stage1_7[205]}
   );
   gpc1_1 gpc764 (
      {stage0_7[511]},
      {stage1_7[206]}
   );
   gpc1_1 gpc765 (
      {stage0_9[476]},
      {stage1_9[228]}
   );
   gpc1_1 gpc766 (
      {stage0_9[477]},
      {stage1_9[229]}
   );
   gpc1_1 gpc767 (
      {stage0_9[478]},
      {stage1_9[230]}
   );
   gpc1_1 gpc768 (
      {stage0_9[479]},
      {stage1_9[231]}
   );
   gpc1_1 gpc769 (
      {stage0_9[480]},
      {stage1_9[232]}
   );
   gpc1_1 gpc770 (
      {stage0_9[481]},
      {stage1_9[233]}
   );
   gpc1_1 gpc771 (
      {stage0_9[482]},
      {stage1_9[234]}
   );
   gpc1_1 gpc772 (
      {stage0_9[483]},
      {stage1_9[235]}
   );
   gpc1_1 gpc773 (
      {stage0_9[484]},
      {stage1_9[236]}
   );
   gpc1_1 gpc774 (
      {stage0_9[485]},
      {stage1_9[237]}
   );
   gpc1_1 gpc775 (
      {stage0_9[486]},
      {stage1_9[238]}
   );
   gpc1_1 gpc776 (
      {stage0_9[487]},
      {stage1_9[239]}
   );
   gpc1_1 gpc777 (
      {stage0_9[488]},
      {stage1_9[240]}
   );
   gpc1_1 gpc778 (
      {stage0_9[489]},
      {stage1_9[241]}
   );
   gpc1_1 gpc779 (
      {stage0_9[490]},
      {stage1_9[242]}
   );
   gpc1_1 gpc780 (
      {stage0_9[491]},
      {stage1_9[243]}
   );
   gpc1_1 gpc781 (
      {stage0_9[492]},
      {stage1_9[244]}
   );
   gpc1_1 gpc782 (
      {stage0_9[493]},
      {stage1_9[245]}
   );
   gpc1_1 gpc783 (
      {stage0_9[494]},
      {stage1_9[246]}
   );
   gpc1_1 gpc784 (
      {stage0_9[495]},
      {stage1_9[247]}
   );
   gpc1_1 gpc785 (
      {stage0_9[496]},
      {stage1_9[248]}
   );
   gpc1_1 gpc786 (
      {stage0_9[497]},
      {stage1_9[249]}
   );
   gpc1_1 gpc787 (
      {stage0_9[498]},
      {stage1_9[250]}
   );
   gpc1_1 gpc788 (
      {stage0_9[499]},
      {stage1_9[251]}
   );
   gpc1_1 gpc789 (
      {stage0_9[500]},
      {stage1_9[252]}
   );
   gpc1_1 gpc790 (
      {stage0_9[501]},
      {stage1_9[253]}
   );
   gpc1_1 gpc791 (
      {stage0_9[502]},
      {stage1_9[254]}
   );
   gpc1_1 gpc792 (
      {stage0_9[503]},
      {stage1_9[255]}
   );
   gpc1_1 gpc793 (
      {stage0_9[504]},
      {stage1_9[256]}
   );
   gpc1_1 gpc794 (
      {stage0_9[505]},
      {stage1_9[257]}
   );
   gpc1_1 gpc795 (
      {stage0_9[506]},
      {stage1_9[258]}
   );
   gpc1_1 gpc796 (
      {stage0_9[507]},
      {stage1_9[259]}
   );
   gpc1_1 gpc797 (
      {stage0_9[508]},
      {stage1_9[260]}
   );
   gpc1_1 gpc798 (
      {stage0_9[509]},
      {stage1_9[261]}
   );
   gpc1_1 gpc799 (
      {stage0_9[510]},
      {stage1_9[262]}
   );
   gpc1_1 gpc800 (
      {stage0_9[511]},
      {stage1_9[263]}
   );
   gpc1_1 gpc801 (
      {stage0_10[504]},
      {stage1_10[202]}
   );
   gpc1_1 gpc802 (
      {stage0_10[505]},
      {stage1_10[203]}
   );
   gpc1_1 gpc803 (
      {stage0_10[506]},
      {stage1_10[204]}
   );
   gpc1_1 gpc804 (
      {stage0_10[507]},
      {stage1_10[205]}
   );
   gpc1_1 gpc805 (
      {stage0_10[508]},
      {stage1_10[206]}
   );
   gpc1_1 gpc806 (
      {stage0_10[509]},
      {stage1_10[207]}
   );
   gpc1_1 gpc807 (
      {stage0_10[510]},
      {stage1_10[208]}
   );
   gpc1_1 gpc808 (
      {stage0_10[511]},
      {stage1_10[209]}
   );
   gpc1_1 gpc809 (
      {stage0_11[506]},
      {stage1_11[184]}
   );
   gpc1_1 gpc810 (
      {stage0_11[507]},
      {stage1_11[185]}
   );
   gpc1_1 gpc811 (
      {stage0_11[508]},
      {stage1_11[186]}
   );
   gpc1_1 gpc812 (
      {stage0_11[509]},
      {stage1_11[187]}
   );
   gpc1_1 gpc813 (
      {stage0_11[510]},
      {stage1_11[188]}
   );
   gpc1_1 gpc814 (
      {stage0_11[511]},
      {stage1_11[189]}
   );
   gpc1_1 gpc815 (
      {stage0_13[467]},
      {stage1_13[237]}
   );
   gpc1_1 gpc816 (
      {stage0_13[468]},
      {stage1_13[238]}
   );
   gpc1_1 gpc817 (
      {stage0_13[469]},
      {stage1_13[239]}
   );
   gpc1_1 gpc818 (
      {stage0_13[470]},
      {stage1_13[240]}
   );
   gpc1_1 gpc819 (
      {stage0_13[471]},
      {stage1_13[241]}
   );
   gpc1_1 gpc820 (
      {stage0_13[472]},
      {stage1_13[242]}
   );
   gpc1_1 gpc821 (
      {stage0_13[473]},
      {stage1_13[243]}
   );
   gpc1_1 gpc822 (
      {stage0_13[474]},
      {stage1_13[244]}
   );
   gpc1_1 gpc823 (
      {stage0_13[475]},
      {stage1_13[245]}
   );
   gpc1_1 gpc824 (
      {stage0_13[476]},
      {stage1_13[246]}
   );
   gpc1_1 gpc825 (
      {stage0_13[477]},
      {stage1_13[247]}
   );
   gpc1_1 gpc826 (
      {stage0_13[478]},
      {stage1_13[248]}
   );
   gpc1_1 gpc827 (
      {stage0_13[479]},
      {stage1_13[249]}
   );
   gpc1_1 gpc828 (
      {stage0_13[480]},
      {stage1_13[250]}
   );
   gpc1_1 gpc829 (
      {stage0_13[481]},
      {stage1_13[251]}
   );
   gpc1_1 gpc830 (
      {stage0_13[482]},
      {stage1_13[252]}
   );
   gpc1_1 gpc831 (
      {stage0_13[483]},
      {stage1_13[253]}
   );
   gpc1_1 gpc832 (
      {stage0_13[484]},
      {stage1_13[254]}
   );
   gpc1_1 gpc833 (
      {stage0_13[485]},
      {stage1_13[255]}
   );
   gpc1_1 gpc834 (
      {stage0_13[486]},
      {stage1_13[256]}
   );
   gpc1_1 gpc835 (
      {stage0_13[487]},
      {stage1_13[257]}
   );
   gpc1_1 gpc836 (
      {stage0_13[488]},
      {stage1_13[258]}
   );
   gpc1_1 gpc837 (
      {stage0_13[489]},
      {stage1_13[259]}
   );
   gpc1_1 gpc838 (
      {stage0_13[490]},
      {stage1_13[260]}
   );
   gpc1_1 gpc839 (
      {stage0_13[491]},
      {stage1_13[261]}
   );
   gpc1_1 gpc840 (
      {stage0_13[492]},
      {stage1_13[262]}
   );
   gpc1_1 gpc841 (
      {stage0_13[493]},
      {stage1_13[263]}
   );
   gpc1_1 gpc842 (
      {stage0_13[494]},
      {stage1_13[264]}
   );
   gpc1_1 gpc843 (
      {stage0_13[495]},
      {stage1_13[265]}
   );
   gpc1_1 gpc844 (
      {stage0_13[496]},
      {stage1_13[266]}
   );
   gpc1_1 gpc845 (
      {stage0_13[497]},
      {stage1_13[267]}
   );
   gpc1_1 gpc846 (
      {stage0_13[498]},
      {stage1_13[268]}
   );
   gpc1_1 gpc847 (
      {stage0_13[499]},
      {stage1_13[269]}
   );
   gpc1_1 gpc848 (
      {stage0_13[500]},
      {stage1_13[270]}
   );
   gpc1_1 gpc849 (
      {stage0_13[501]},
      {stage1_13[271]}
   );
   gpc1_1 gpc850 (
      {stage0_13[502]},
      {stage1_13[272]}
   );
   gpc1_1 gpc851 (
      {stage0_13[503]},
      {stage1_13[273]}
   );
   gpc1_1 gpc852 (
      {stage0_13[504]},
      {stage1_13[274]}
   );
   gpc1_1 gpc853 (
      {stage0_13[505]},
      {stage1_13[275]}
   );
   gpc1_1 gpc854 (
      {stage0_13[506]},
      {stage1_13[276]}
   );
   gpc1_1 gpc855 (
      {stage0_13[507]},
      {stage1_13[277]}
   );
   gpc1_1 gpc856 (
      {stage0_13[508]},
      {stage1_13[278]}
   );
   gpc1_1 gpc857 (
      {stage0_13[509]},
      {stage1_13[279]}
   );
   gpc1_1 gpc858 (
      {stage0_13[510]},
      {stage1_13[280]}
   );
   gpc1_1 gpc859 (
      {stage0_13[511]},
      {stage1_13[281]}
   );
   gpc1_1 gpc860 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc861 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc862 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc863 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc864 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc865 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc866 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc867 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc868 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc869 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc870 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc871 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc872 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc873 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc874 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc875 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc876 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc877 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc878 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc879 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc880 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc881 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc882 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc883 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc884 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc885 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc886 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc887 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc888 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc889 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc890 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc891 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc892 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc893 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc894 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc895 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc896 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc897 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc898 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc899 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc900 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc901 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc902 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc903 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc904 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc905 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc906 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc907 (
      {stage0_14[486]},
      {stage1_14[219]}
   );
   gpc1_1 gpc908 (
      {stage0_14[487]},
      {stage1_14[220]}
   );
   gpc1_1 gpc909 (
      {stage0_14[488]},
      {stage1_14[221]}
   );
   gpc1_1 gpc910 (
      {stage0_14[489]},
      {stage1_14[222]}
   );
   gpc1_1 gpc911 (
      {stage0_14[490]},
      {stage1_14[223]}
   );
   gpc1_1 gpc912 (
      {stage0_14[491]},
      {stage1_14[224]}
   );
   gpc1_1 gpc913 (
      {stage0_14[492]},
      {stage1_14[225]}
   );
   gpc1_1 gpc914 (
      {stage0_14[493]},
      {stage1_14[226]}
   );
   gpc1_1 gpc915 (
      {stage0_14[494]},
      {stage1_14[227]}
   );
   gpc1_1 gpc916 (
      {stage0_14[495]},
      {stage1_14[228]}
   );
   gpc1_1 gpc917 (
      {stage0_14[496]},
      {stage1_14[229]}
   );
   gpc1_1 gpc918 (
      {stage0_14[497]},
      {stage1_14[230]}
   );
   gpc1_1 gpc919 (
      {stage0_14[498]},
      {stage1_14[231]}
   );
   gpc1_1 gpc920 (
      {stage0_14[499]},
      {stage1_14[232]}
   );
   gpc1_1 gpc921 (
      {stage0_14[500]},
      {stage1_14[233]}
   );
   gpc1_1 gpc922 (
      {stage0_14[501]},
      {stage1_14[234]}
   );
   gpc1_1 gpc923 (
      {stage0_14[502]},
      {stage1_14[235]}
   );
   gpc1_1 gpc924 (
      {stage0_14[503]},
      {stage1_14[236]}
   );
   gpc1_1 gpc925 (
      {stage0_14[504]},
      {stage1_14[237]}
   );
   gpc1_1 gpc926 (
      {stage0_14[505]},
      {stage1_14[238]}
   );
   gpc1_1 gpc927 (
      {stage0_14[506]},
      {stage1_14[239]}
   );
   gpc1_1 gpc928 (
      {stage0_14[507]},
      {stage1_14[240]}
   );
   gpc1_1 gpc929 (
      {stage0_14[508]},
      {stage1_14[241]}
   );
   gpc1_1 gpc930 (
      {stage0_14[509]},
      {stage1_14[242]}
   );
   gpc1_1 gpc931 (
      {stage0_14[510]},
      {stage1_14[243]}
   );
   gpc1_1 gpc932 (
      {stage0_14[511]},
      {stage1_14[244]}
   );
   gpc1_1 gpc933 (
      {stage0_15[384]},
      {stage1_15[144]}
   );
   gpc1_1 gpc934 (
      {stage0_15[385]},
      {stage1_15[145]}
   );
   gpc1_1 gpc935 (
      {stage0_15[386]},
      {stage1_15[146]}
   );
   gpc1_1 gpc936 (
      {stage0_15[387]},
      {stage1_15[147]}
   );
   gpc1_1 gpc937 (
      {stage0_15[388]},
      {stage1_15[148]}
   );
   gpc1_1 gpc938 (
      {stage0_15[389]},
      {stage1_15[149]}
   );
   gpc1_1 gpc939 (
      {stage0_15[390]},
      {stage1_15[150]}
   );
   gpc1_1 gpc940 (
      {stage0_15[391]},
      {stage1_15[151]}
   );
   gpc1_1 gpc941 (
      {stage0_15[392]},
      {stage1_15[152]}
   );
   gpc1_1 gpc942 (
      {stage0_15[393]},
      {stage1_15[153]}
   );
   gpc1_1 gpc943 (
      {stage0_15[394]},
      {stage1_15[154]}
   );
   gpc1_1 gpc944 (
      {stage0_15[395]},
      {stage1_15[155]}
   );
   gpc1_1 gpc945 (
      {stage0_15[396]},
      {stage1_15[156]}
   );
   gpc1_1 gpc946 (
      {stage0_15[397]},
      {stage1_15[157]}
   );
   gpc1_1 gpc947 (
      {stage0_15[398]},
      {stage1_15[158]}
   );
   gpc1_1 gpc948 (
      {stage0_15[399]},
      {stage1_15[159]}
   );
   gpc1_1 gpc949 (
      {stage0_15[400]},
      {stage1_15[160]}
   );
   gpc1_1 gpc950 (
      {stage0_15[401]},
      {stage1_15[161]}
   );
   gpc1_1 gpc951 (
      {stage0_15[402]},
      {stage1_15[162]}
   );
   gpc1_1 gpc952 (
      {stage0_15[403]},
      {stage1_15[163]}
   );
   gpc1_1 gpc953 (
      {stage0_15[404]},
      {stage1_15[164]}
   );
   gpc1_1 gpc954 (
      {stage0_15[405]},
      {stage1_15[165]}
   );
   gpc1_1 gpc955 (
      {stage0_15[406]},
      {stage1_15[166]}
   );
   gpc1_1 gpc956 (
      {stage0_15[407]},
      {stage1_15[167]}
   );
   gpc1_1 gpc957 (
      {stage0_15[408]},
      {stage1_15[168]}
   );
   gpc1_1 gpc958 (
      {stage0_15[409]},
      {stage1_15[169]}
   );
   gpc1_1 gpc959 (
      {stage0_15[410]},
      {stage1_15[170]}
   );
   gpc1_1 gpc960 (
      {stage0_15[411]},
      {stage1_15[171]}
   );
   gpc1_1 gpc961 (
      {stage0_15[412]},
      {stage1_15[172]}
   );
   gpc1_1 gpc962 (
      {stage0_15[413]},
      {stage1_15[173]}
   );
   gpc1_1 gpc963 (
      {stage0_15[414]},
      {stage1_15[174]}
   );
   gpc1_1 gpc964 (
      {stage0_15[415]},
      {stage1_15[175]}
   );
   gpc1_1 gpc965 (
      {stage0_15[416]},
      {stage1_15[176]}
   );
   gpc1_1 gpc966 (
      {stage0_15[417]},
      {stage1_15[177]}
   );
   gpc1_1 gpc967 (
      {stage0_15[418]},
      {stage1_15[178]}
   );
   gpc1_1 gpc968 (
      {stage0_15[419]},
      {stage1_15[179]}
   );
   gpc1_1 gpc969 (
      {stage0_15[420]},
      {stage1_15[180]}
   );
   gpc1_1 gpc970 (
      {stage0_15[421]},
      {stage1_15[181]}
   );
   gpc1_1 gpc971 (
      {stage0_15[422]},
      {stage1_15[182]}
   );
   gpc1_1 gpc972 (
      {stage0_15[423]},
      {stage1_15[183]}
   );
   gpc1_1 gpc973 (
      {stage0_15[424]},
      {stage1_15[184]}
   );
   gpc1_1 gpc974 (
      {stage0_15[425]},
      {stage1_15[185]}
   );
   gpc1_1 gpc975 (
      {stage0_15[426]},
      {stage1_15[186]}
   );
   gpc1_1 gpc976 (
      {stage0_15[427]},
      {stage1_15[187]}
   );
   gpc1_1 gpc977 (
      {stage0_15[428]},
      {stage1_15[188]}
   );
   gpc1_1 gpc978 (
      {stage0_15[429]},
      {stage1_15[189]}
   );
   gpc1_1 gpc979 (
      {stage0_15[430]},
      {stage1_15[190]}
   );
   gpc1_1 gpc980 (
      {stage0_15[431]},
      {stage1_15[191]}
   );
   gpc1_1 gpc981 (
      {stage0_15[432]},
      {stage1_15[192]}
   );
   gpc1_1 gpc982 (
      {stage0_15[433]},
      {stage1_15[193]}
   );
   gpc1_1 gpc983 (
      {stage0_15[434]},
      {stage1_15[194]}
   );
   gpc1_1 gpc984 (
      {stage0_15[435]},
      {stage1_15[195]}
   );
   gpc1_1 gpc985 (
      {stage0_15[436]},
      {stage1_15[196]}
   );
   gpc1_1 gpc986 (
      {stage0_15[437]},
      {stage1_15[197]}
   );
   gpc1_1 gpc987 (
      {stage0_15[438]},
      {stage1_15[198]}
   );
   gpc1_1 gpc988 (
      {stage0_15[439]},
      {stage1_15[199]}
   );
   gpc1_1 gpc989 (
      {stage0_15[440]},
      {stage1_15[200]}
   );
   gpc1_1 gpc990 (
      {stage0_15[441]},
      {stage1_15[201]}
   );
   gpc1_1 gpc991 (
      {stage0_15[442]},
      {stage1_15[202]}
   );
   gpc1_1 gpc992 (
      {stage0_15[443]},
      {stage1_15[203]}
   );
   gpc1_1 gpc993 (
      {stage0_15[444]},
      {stage1_15[204]}
   );
   gpc1_1 gpc994 (
      {stage0_15[445]},
      {stage1_15[205]}
   );
   gpc1_1 gpc995 (
      {stage0_15[446]},
      {stage1_15[206]}
   );
   gpc1_1 gpc996 (
      {stage0_15[447]},
      {stage1_15[207]}
   );
   gpc1_1 gpc997 (
      {stage0_15[448]},
      {stage1_15[208]}
   );
   gpc1_1 gpc998 (
      {stage0_15[449]},
      {stage1_15[209]}
   );
   gpc1_1 gpc999 (
      {stage0_15[450]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[451]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[452]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[453]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[454]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[455]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[456]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[457]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1007 (
      {stage0_15[458]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1008 (
      {stage0_15[459]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1009 (
      {stage0_15[460]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1010 (
      {stage0_15[461]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1011 (
      {stage0_15[462]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1012 (
      {stage0_15[463]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1013 (
      {stage0_15[464]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1014 (
      {stage0_15[465]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1015 (
      {stage0_15[466]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1016 (
      {stage0_15[467]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1017 (
      {stage0_15[468]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1018 (
      {stage0_15[469]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1019 (
      {stage0_15[470]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1020 (
      {stage0_15[471]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1021 (
      {stage0_15[472]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1022 (
      {stage0_15[473]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1023 (
      {stage0_15[474]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1024 (
      {stage0_15[475]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1025 (
      {stage0_15[476]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1026 (
      {stage0_15[477]},
      {stage1_15[237]}
   );
   gpc1_1 gpc1027 (
      {stage0_15[478]},
      {stage1_15[238]}
   );
   gpc1_1 gpc1028 (
      {stage0_15[479]},
      {stage1_15[239]}
   );
   gpc1_1 gpc1029 (
      {stage0_15[480]},
      {stage1_15[240]}
   );
   gpc1_1 gpc1030 (
      {stage0_15[481]},
      {stage1_15[241]}
   );
   gpc1_1 gpc1031 (
      {stage0_15[482]},
      {stage1_15[242]}
   );
   gpc1_1 gpc1032 (
      {stage0_15[483]},
      {stage1_15[243]}
   );
   gpc1_1 gpc1033 (
      {stage0_15[484]},
      {stage1_15[244]}
   );
   gpc1_1 gpc1034 (
      {stage0_15[485]},
      {stage1_15[245]}
   );
   gpc1_1 gpc1035 (
      {stage0_15[486]},
      {stage1_15[246]}
   );
   gpc1_1 gpc1036 (
      {stage0_15[487]},
      {stage1_15[247]}
   );
   gpc1_1 gpc1037 (
      {stage0_15[488]},
      {stage1_15[248]}
   );
   gpc1_1 gpc1038 (
      {stage0_15[489]},
      {stage1_15[249]}
   );
   gpc1_1 gpc1039 (
      {stage0_15[490]},
      {stage1_15[250]}
   );
   gpc1_1 gpc1040 (
      {stage0_15[491]},
      {stage1_15[251]}
   );
   gpc1_1 gpc1041 (
      {stage0_15[492]},
      {stage1_15[252]}
   );
   gpc1_1 gpc1042 (
      {stage0_15[493]},
      {stage1_15[253]}
   );
   gpc1_1 gpc1043 (
      {stage0_15[494]},
      {stage1_15[254]}
   );
   gpc1_1 gpc1044 (
      {stage0_15[495]},
      {stage1_15[255]}
   );
   gpc1_1 gpc1045 (
      {stage0_15[496]},
      {stage1_15[256]}
   );
   gpc1_1 gpc1046 (
      {stage0_15[497]},
      {stage1_15[257]}
   );
   gpc1_1 gpc1047 (
      {stage0_15[498]},
      {stage1_15[258]}
   );
   gpc1_1 gpc1048 (
      {stage0_15[499]},
      {stage1_15[259]}
   );
   gpc1_1 gpc1049 (
      {stage0_15[500]},
      {stage1_15[260]}
   );
   gpc1_1 gpc1050 (
      {stage0_15[501]},
      {stage1_15[261]}
   );
   gpc1_1 gpc1051 (
      {stage0_15[502]},
      {stage1_15[262]}
   );
   gpc1_1 gpc1052 (
      {stage0_15[503]},
      {stage1_15[263]}
   );
   gpc1_1 gpc1053 (
      {stage0_15[504]},
      {stage1_15[264]}
   );
   gpc1_1 gpc1054 (
      {stage0_15[505]},
      {stage1_15[265]}
   );
   gpc1_1 gpc1055 (
      {stage0_15[506]},
      {stage1_15[266]}
   );
   gpc1_1 gpc1056 (
      {stage0_15[507]},
      {stage1_15[267]}
   );
   gpc1_1 gpc1057 (
      {stage0_15[508]},
      {stage1_15[268]}
   );
   gpc1_1 gpc1058 (
      {stage0_15[509]},
      {stage1_15[269]}
   );
   gpc1_1 gpc1059 (
      {stage0_15[510]},
      {stage1_15[270]}
   );
   gpc1_1 gpc1060 (
      {stage0_15[511]},
      {stage1_15[271]}
   );
   gpc1163_5 gpc1061 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1062 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1063 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1064 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1065 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1066 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1067 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1068 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1069 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1070 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1071 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1072 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1073 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1074 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1075 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1076 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1077 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1078 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1079 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1080 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1081 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1082 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc615_5 gpc1083 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100]},
      {stage1_1[72]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1084 (
      {stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc1085 (
      {stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc1086 (
      {stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc1087 (
      {stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc1088 (
      {stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc1089 (
      {stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1090 (
      {stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1091 (
      {stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1092 (
      {stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1093 (
      {stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1094 (
      {stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1095 (
      {stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1096 (
      {stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc1097 (
      {stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc1098 (
      {stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc1099 (
      {stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc1100 (
      {stage1_1[169], stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc1101 (
      {stage1_1[175], stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], 1'b0},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc615_5 gpc1102 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[120]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1103 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[121]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1104 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[122]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1105 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[123]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc1106 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[124]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc1107 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[125]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc1108 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[126]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc1109 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[127]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc1110 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[128]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc1111 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[129]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc1112 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[130]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc1113 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[131]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc1114 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[132]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc1115 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[133]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[31],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc1116 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[134]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[32],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc1117 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[135]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[33],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc1118 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[136]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[34],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc1119 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[137]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[35],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc1120 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[138]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[36],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc615_5 gpc1121 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[114]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[19],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1122 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[115]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[20],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1123 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[116]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[21],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1124 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[117]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[22],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1125 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[118]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[23],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1126 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[119]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[24],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1127 (
      {stage1_3[169], stage1_3[170], stage1_3[171], stage1_3[172], stage1_3[173]},
      {stage1_4[120]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[25],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1128 (
      {stage1_3[174], stage1_3[175], stage1_3[176], stage1_3[177], stage1_3[178]},
      {stage1_4[121]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[26],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1129 (
      {stage1_3[179], stage1_3[180], stage1_3[181], stage1_3[182], stage1_3[183]},
      {stage1_4[122]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[27],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1130 (
      {stage1_3[184], stage1_3[185], stage1_3[186], stage1_3[187], stage1_3[188]},
      {stage1_4[123]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[28],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1131 (
      {stage1_3[189], stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193]},
      {stage1_4[124]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[29],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1132 (
      {stage1_3[194], stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198]},
      {stage1_4[125]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[30],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1133 (
      {stage1_3[199], stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203]},
      {stage1_4[126]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[31],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1134 (
      {stage1_3[204], stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208]},
      {stage1_4[127]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[32],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1135 (
      {stage1_3[209], stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213]},
      {stage1_4[128]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[33],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1136 (
      {stage1_3[214], stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218]},
      {stage1_4[129]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[34],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc606_5 gpc1137 (
      {stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[16],stage2_6[35],stage2_5[53],stage2_4[76]}
   );
   gpc606_5 gpc1138 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[17],stage2_6[36],stage2_5[54],stage2_4[77]}
   );
   gpc606_5 gpc1139 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[18],stage2_6[37],stage2_5[55],stage2_4[78]}
   );
   gpc606_5 gpc1140 (
      {stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[19],stage2_6[38],stage2_5[56],stage2_4[79]}
   );
   gpc606_5 gpc1141 (
      {stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[20],stage2_6[39],stage2_5[57],stage2_4[80]}
   );
   gpc606_5 gpc1142 (
      {stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[21],stage2_6[40],stage2_5[58],stage2_4[81]}
   );
   gpc606_5 gpc1143 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[22],stage2_6[41],stage2_5[59],stage2_4[82]}
   );
   gpc606_5 gpc1144 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[23],stage2_6[42],stage2_5[60],stage2_4[83]}
   );
   gpc606_5 gpc1145 (
      {stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[24],stage2_6[43],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc1146 (
      {stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[25],stage2_6[44],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc1147 (
      {stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[26],stage2_6[45],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc1148 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[27],stage2_6[46],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc1149 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206], stage1_4[207]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[28],stage2_6[47],stage2_5[65],stage2_4[88]}
   );
   gpc606_5 gpc1150 (
      {stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211], stage1_4[212], stage1_4[213]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[29],stage2_6[48],stage2_5[66],stage2_4[89]}
   );
   gpc606_5 gpc1151 (
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[14],stage2_7[30],stage2_6[49],stage2_5[67]}
   );
   gpc606_5 gpc1152 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[15],stage2_7[31],stage2_6[50],stage2_5[68]}
   );
   gpc606_5 gpc1153 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[16],stage2_7[32],stage2_6[51],stage2_5[69]}
   );
   gpc606_5 gpc1154 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[17],stage2_7[33],stage2_6[52],stage2_5[70]}
   );
   gpc606_5 gpc1155 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[18],stage2_7[34],stage2_6[53],stage2_5[71]}
   );
   gpc606_5 gpc1156 (
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[19],stage2_7[35],stage2_6[54],stage2_5[72]}
   );
   gpc606_5 gpc1157 (
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[20],stage2_7[36],stage2_6[55],stage2_5[73]}
   );
   gpc606_5 gpc1158 (
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[21],stage2_7[37],stage2_6[56],stage2_5[74]}
   );
   gpc606_5 gpc1159 (
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[22],stage2_7[38],stage2_6[57],stage2_5[75]}
   );
   gpc606_5 gpc1160 (
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[23],stage2_7[39],stage2_6[58],stage2_5[76]}
   );
   gpc606_5 gpc1161 (
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[24],stage2_7[40],stage2_6[59],stage2_5[77]}
   );
   gpc606_5 gpc1162 (
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[25],stage2_7[41],stage2_6[60],stage2_5[78]}
   );
   gpc606_5 gpc1163 (
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[26],stage2_7[42],stage2_6[61],stage2_5[79]}
   );
   gpc606_5 gpc1164 (
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[27],stage2_7[43],stage2_6[62],stage2_5[80]}
   );
   gpc606_5 gpc1165 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[28],stage2_7[44],stage2_6[63],stage2_5[81]}
   );
   gpc606_5 gpc1166 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[29],stage2_7[45],stage2_6[64],stage2_5[82]}
   );
   gpc606_5 gpc1167 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[30],stage2_7[46],stage2_6[65],stage2_5[83]}
   );
   gpc606_5 gpc1168 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[31],stage2_7[47],stage2_6[66],stage2_5[84]}
   );
   gpc606_5 gpc1169 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[32],stage2_7[48],stage2_6[67],stage2_5[85]}
   );
   gpc606_5 gpc1170 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[19],stage2_8[33],stage2_7[49],stage2_6[68]}
   );
   gpc606_5 gpc1171 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[20],stage2_8[34],stage2_7[50],stage2_6[69]}
   );
   gpc606_5 gpc1172 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[21],stage2_8[35],stage2_7[51],stage2_6[70]}
   );
   gpc606_5 gpc1173 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[22],stage2_8[36],stage2_7[52],stage2_6[71]}
   );
   gpc606_5 gpc1174 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[23],stage2_8[37],stage2_7[53],stage2_6[72]}
   );
   gpc606_5 gpc1175 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[24],stage2_8[38],stage2_7[54],stage2_6[73]}
   );
   gpc606_5 gpc1176 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[25],stage2_8[39],stage2_7[55],stage2_6[74]}
   );
   gpc606_5 gpc1177 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[26],stage2_8[40],stage2_7[56],stage2_6[75]}
   );
   gpc606_5 gpc1178 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[27],stage2_8[41],stage2_7[57],stage2_6[76]}
   );
   gpc606_5 gpc1179 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[28],stage2_8[42],stage2_7[58],stage2_6[77]}
   );
   gpc606_5 gpc1180 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[29],stage2_8[43],stage2_7[59],stage2_6[78]}
   );
   gpc606_5 gpc1181 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[30],stage2_8[44],stage2_7[60],stage2_6[79]}
   );
   gpc606_5 gpc1182 (
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[31],stage2_8[45],stage2_7[61],stage2_6[80]}
   );
   gpc606_5 gpc1183 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[32],stage2_8[46],stage2_7[62],stage2_6[81]}
   );
   gpc606_5 gpc1184 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[33],stage2_8[47],stage2_7[63],stage2_6[82]}
   );
   gpc615_5 gpc1185 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178]},
      {stage1_7[114]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[34],stage2_8[48],stage2_7[64],stage2_6[83]}
   );
   gpc615_5 gpc1186 (
      {stage1_6[179], stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183]},
      {stage1_7[115]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[35],stage2_8[49],stage2_7[65],stage2_6[84]}
   );
   gpc615_5 gpc1187 (
      {stage1_6[184], stage1_6[185], stage1_6[186], stage1_6[187], stage1_6[188]},
      {stage1_7[116]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[36],stage2_8[50],stage2_7[66],stage2_6[85]}
   );
   gpc615_5 gpc1188 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[108]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[18],stage2_9[37],stage2_8[51],stage2_7[67]}
   );
   gpc615_5 gpc1189 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[109]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[19],stage2_9[38],stage2_8[52],stage2_7[68]}
   );
   gpc615_5 gpc1190 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[110]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[20],stage2_9[39],stage2_8[53],stage2_7[69]}
   );
   gpc615_5 gpc1191 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[111]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[21],stage2_9[40],stage2_8[54],stage2_7[70]}
   );
   gpc615_5 gpc1192 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[112]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[22],stage2_9[41],stage2_8[55],stage2_7[71]}
   );
   gpc615_5 gpc1193 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[113]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[23],stage2_9[42],stage2_8[56],stage2_7[72]}
   );
   gpc615_5 gpc1194 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[114]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[24],stage2_9[43],stage2_8[57],stage2_7[73]}
   );
   gpc615_5 gpc1195 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[115]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[25],stage2_9[44],stage2_8[58],stage2_7[74]}
   );
   gpc615_5 gpc1196 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[116]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[26],stage2_9[45],stage2_8[59],stage2_7[75]}
   );
   gpc615_5 gpc1197 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[117]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[27],stage2_9[46],stage2_8[60],stage2_7[76]}
   );
   gpc615_5 gpc1198 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[118]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[28],stage2_9[47],stage2_8[61],stage2_7[77]}
   );
   gpc615_5 gpc1199 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[119]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[29],stage2_9[48],stage2_8[62],stage2_7[78]}
   );
   gpc615_5 gpc1200 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[120]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[30],stage2_9[49],stage2_8[63],stage2_7[79]}
   );
   gpc615_5 gpc1201 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[121]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[31],stage2_9[50],stage2_8[64],stage2_7[80]}
   );
   gpc615_5 gpc1202 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[122]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[32],stage2_9[51],stage2_8[65],stage2_7[81]}
   );
   gpc615_5 gpc1203 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[123]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[33],stage2_9[52],stage2_8[66],stage2_7[82]}
   );
   gpc615_5 gpc1204 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[124]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[34],stage2_9[53],stage2_8[67],stage2_7[83]}
   );
   gpc615_5 gpc1205 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[125]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[35],stage2_9[54],stage2_8[68],stage2_7[84]}
   );
   gpc606_5 gpc1206 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[18],stage2_10[36],stage2_9[55],stage2_8[69]}
   );
   gpc606_5 gpc1207 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[19],stage2_10[37],stage2_9[56],stage2_8[70]}
   );
   gpc615_5 gpc1208 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142]},
      {stage1_9[108]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[20],stage2_10[38],stage2_9[57],stage2_8[71]}
   );
   gpc615_5 gpc1209 (
      {stage1_8[143], stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147]},
      {stage1_9[109]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[21],stage2_10[39],stage2_9[58],stage2_8[72]}
   );
   gpc615_5 gpc1210 (
      {stage1_8[148], stage1_8[149], stage1_8[150], stage1_8[151], stage1_8[152]},
      {stage1_9[110]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[22],stage2_10[40],stage2_9[59],stage2_8[73]}
   );
   gpc615_5 gpc1211 (
      {stage1_8[153], stage1_8[154], stage1_8[155], stage1_8[156], stage1_8[157]},
      {stage1_9[111]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[23],stage2_10[41],stage2_9[60],stage2_8[74]}
   );
   gpc615_5 gpc1212 (
      {stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161], stage1_8[162]},
      {stage1_9[112]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[24],stage2_10[42],stage2_9[61],stage2_8[75]}
   );
   gpc615_5 gpc1213 (
      {stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_9[113]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[25],stage2_10[43],stage2_9[62],stage2_8[76]}
   );
   gpc615_5 gpc1214 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172]},
      {stage1_9[114]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[26],stage2_10[44],stage2_9[63],stage2_8[77]}
   );
   gpc615_5 gpc1215 (
      {stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_9[115]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[27],stage2_10[45],stage2_9[64],stage2_8[78]}
   );
   gpc615_5 gpc1216 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_9[116]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[28],stage2_10[46],stage2_9[65],stage2_8[79]}
   );
   gpc615_5 gpc1217 (
      {stage1_8[183], stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187]},
      {stage1_9[117]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[29],stage2_10[47],stage2_9[66],stage2_8[80]}
   );
   gpc615_5 gpc1218 (
      {stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_9[118]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[30],stage2_10[48],stage2_9[67],stage2_8[81]}
   );
   gpc615_5 gpc1219 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197]},
      {stage1_9[119]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[31],stage2_10[49],stage2_9[68],stage2_8[82]}
   );
   gpc615_5 gpc1220 (
      {stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202]},
      {stage1_9[120]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[32],stage2_10[50],stage2_9[69],stage2_8[83]}
   );
   gpc615_5 gpc1221 (
      {stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_9[121]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[33],stage2_10[51],stage2_9[70],stage2_8[84]}
   );
   gpc615_5 gpc1222 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212]},
      {stage1_9[122]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[34],stage2_10[52],stage2_9[71],stage2_8[85]}
   );
   gpc615_5 gpc1223 (
      {stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217]},
      {stage1_9[123]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[35],stage2_10[53],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc1224 (
      {stage1_9[124], stage1_9[125], stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[36],stage2_10[54],stage2_9[73]}
   );
   gpc606_5 gpc1225 (
      {stage1_9[130], stage1_9[131], stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[37],stage2_10[55],stage2_9[74]}
   );
   gpc606_5 gpc1226 (
      {stage1_9[136], stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[38],stage2_10[56],stage2_9[75]}
   );
   gpc606_5 gpc1227 (
      {stage1_9[142], stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[21],stage2_11[39],stage2_10[57],stage2_9[76]}
   );
   gpc606_5 gpc1228 (
      {stage1_9[148], stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[22],stage2_11[40],stage2_10[58],stage2_9[77]}
   );
   gpc606_5 gpc1229 (
      {stage1_9[154], stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[23],stage2_11[41],stage2_10[59],stage2_9[78]}
   );
   gpc606_5 gpc1230 (
      {stage1_9[160], stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[24],stage2_11[42],stage2_10[60],stage2_9[79]}
   );
   gpc606_5 gpc1231 (
      {stage1_9[166], stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[25],stage2_11[43],stage2_10[61],stage2_9[80]}
   );
   gpc606_5 gpc1232 (
      {stage1_9[172], stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[26],stage2_11[44],stage2_10[62],stage2_9[81]}
   );
   gpc606_5 gpc1233 (
      {stage1_9[178], stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[27],stage2_11[45],stage2_10[63],stage2_9[82]}
   );
   gpc606_5 gpc1234 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[28],stage2_11[46],stage2_10[64],stage2_9[83]}
   );
   gpc606_5 gpc1235 (
      {stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[29],stage2_11[47],stage2_10[65],stage2_9[84]}
   );
   gpc606_5 gpc1236 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[30],stage2_11[48],stage2_10[66],stage2_9[85]}
   );
   gpc606_5 gpc1237 (
      {stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[31],stage2_11[49],stage2_10[67],stage2_9[86]}
   );
   gpc606_5 gpc1238 (
      {stage1_9[208], stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[32],stage2_11[50],stage2_10[68],stage2_9[87]}
   );
   gpc606_5 gpc1239 (
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[15],stage2_12[33],stage2_11[51],stage2_10[69]}
   );
   gpc606_5 gpc1240 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[16],stage2_12[34],stage2_11[52],stage2_10[70]}
   );
   gpc606_5 gpc1241 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[17],stage2_12[35],stage2_11[53],stage2_10[71]}
   );
   gpc606_5 gpc1242 (
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[18],stage2_12[36],stage2_11[54],stage2_10[72]}
   );
   gpc606_5 gpc1243 (
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[19],stage2_12[37],stage2_11[55],stage2_10[73]}
   );
   gpc606_5 gpc1244 (
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[20],stage2_12[38],stage2_11[56],stage2_10[74]}
   );
   gpc606_5 gpc1245 (
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[21],stage2_12[39],stage2_11[57],stage2_10[75]}
   );
   gpc606_5 gpc1246 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[22],stage2_12[40],stage2_11[58],stage2_10[76]}
   );
   gpc606_5 gpc1247 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[23],stage2_12[41],stage2_11[59],stage2_10[77]}
   );
   gpc606_5 gpc1248 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[24],stage2_12[42],stage2_11[60],stage2_10[78]}
   );
   gpc606_5 gpc1249 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[25],stage2_12[43],stage2_11[61],stage2_10[79]}
   );
   gpc606_5 gpc1250 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[26],stage2_12[44],stage2_11[62],stage2_10[80]}
   );
   gpc606_5 gpc1251 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[27],stage2_12[45],stage2_11[63],stage2_10[81]}
   );
   gpc606_5 gpc1252 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[28],stage2_12[46],stage2_11[64],stage2_10[82]}
   );
   gpc606_5 gpc1253 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[29],stage2_12[47],stage2_11[65],stage2_10[83]}
   );
   gpc606_5 gpc1254 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[30],stage2_12[48],stage2_11[66],stage2_10[84]}
   );
   gpc606_5 gpc1255 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[31],stage2_12[49],stage2_11[67],stage2_10[85]}
   );
   gpc615_5 gpc1256 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[17],stage2_13[32],stage2_12[50],stage2_11[68]}
   );
   gpc615_5 gpc1257 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[103]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[18],stage2_13[33],stage2_12[51],stage2_11[69]}
   );
   gpc615_5 gpc1258 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[104]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[19],stage2_13[34],stage2_12[52],stage2_11[70]}
   );
   gpc615_5 gpc1259 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[105]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[20],stage2_13[35],stage2_12[53],stage2_11[71]}
   );
   gpc615_5 gpc1260 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[106]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[21],stage2_13[36],stage2_12[54],stage2_11[72]}
   );
   gpc615_5 gpc1261 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[107]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[22],stage2_13[37],stage2_12[55],stage2_11[73]}
   );
   gpc606_5 gpc1262 (
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[23],stage2_13[38],stage2_12[56]}
   );
   gpc606_5 gpc1263 (
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[24],stage2_13[39],stage2_12[57]}
   );
   gpc606_5 gpc1264 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[8],stage2_14[25],stage2_13[40],stage2_12[58]}
   );
   gpc606_5 gpc1265 (
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[9],stage2_14[26],stage2_13[41],stage2_12[59]}
   );
   gpc606_5 gpc1266 (
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[10],stage2_14[27],stage2_13[42],stage2_12[60]}
   );
   gpc606_5 gpc1267 (
      {stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[11],stage2_14[28],stage2_13[43],stage2_12[61]}
   );
   gpc606_5 gpc1268 (
      {stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[12],stage2_14[29],stage2_13[44],stage2_12[62]}
   );
   gpc606_5 gpc1269 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[13],stage2_14[30],stage2_13[45],stage2_12[63]}
   );
   gpc606_5 gpc1270 (
      {stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[14],stage2_14[31],stage2_13[46],stage2_12[64]}
   );
   gpc606_5 gpc1271 (
      {stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[15],stage2_14[32],stage2_13[47],stage2_12[65]}
   );
   gpc606_5 gpc1272 (
      {stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[16],stage2_14[33],stage2_13[48],stage2_12[66]}
   );
   gpc606_5 gpc1273 (
      {stage1_12[174], stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[17],stage2_14[34],stage2_13[49],stage2_12[67]}
   );
   gpc606_5 gpc1274 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[18],stage2_14[35],stage2_13[50],stage2_12[68]}
   );
   gpc606_5 gpc1275 (
      {stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[19],stage2_14[36],stage2_13[51],stage2_12[69]}
   );
   gpc606_5 gpc1276 (
      {stage1_12[192], stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[20],stage2_14[37],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc1277 (
      {stage1_12[198], stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[21],stage2_14[38],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc1278 (
      {stage1_12[204], stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[22],stage2_14[39],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc1279 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[17],stage2_15[23],stage2_14[40],stage2_13[55]}
   );
   gpc606_5 gpc1280 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[18],stage2_15[24],stage2_14[41],stage2_13[56]}
   );
   gpc606_5 gpc1281 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[19],stage2_15[25],stage2_14[42],stage2_13[57]}
   );
   gpc606_5 gpc1282 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[20],stage2_15[26],stage2_14[43],stage2_13[58]}
   );
   gpc606_5 gpc1283 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[21],stage2_15[27],stage2_14[44],stage2_13[59]}
   );
   gpc606_5 gpc1284 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[22],stage2_15[28],stage2_14[45],stage2_13[60]}
   );
   gpc606_5 gpc1285 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[23],stage2_15[29],stage2_14[46],stage2_13[61]}
   );
   gpc606_5 gpc1286 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[24],stage2_15[30],stage2_14[47],stage2_13[62]}
   );
   gpc606_5 gpc1287 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[25],stage2_15[31],stage2_14[48],stage2_13[63]}
   );
   gpc606_5 gpc1288 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[26],stage2_15[32],stage2_14[49],stage2_13[64]}
   );
   gpc606_5 gpc1289 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[27],stage2_15[33],stage2_14[50],stage2_13[65]}
   );
   gpc606_5 gpc1290 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[28],stage2_15[34],stage2_14[51],stage2_13[66]}
   );
   gpc606_5 gpc1291 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[29],stage2_15[35],stage2_14[52],stage2_13[67]}
   );
   gpc606_5 gpc1292 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[30],stage2_15[36],stage2_14[53],stage2_13[68]}
   );
   gpc606_5 gpc1293 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[31],stage2_15[37],stage2_14[54],stage2_13[69]}
   );
   gpc606_5 gpc1294 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[32],stage2_15[38],stage2_14[55],stage2_13[70]}
   );
   gpc615_5 gpc1295 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136]},
      {stage1_14[102]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[33],stage2_15[39],stage2_14[56],stage2_13[71]}
   );
   gpc615_5 gpc1296 (
      {stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141]},
      {stage1_14[103]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[34],stage2_15[40],stage2_14[57],stage2_13[72]}
   );
   gpc615_5 gpc1297 (
      {stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage1_14[104]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[35],stage2_15[41],stage2_14[58],stage2_13[73]}
   );
   gpc615_5 gpc1298 (
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151]},
      {stage1_14[105]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[36],stage2_15[42],stage2_14[59],stage2_13[74]}
   );
   gpc615_5 gpc1299 (
      {stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156]},
      {stage1_14[106]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[37],stage2_15[43],stage2_14[60],stage2_13[75]}
   );
   gpc615_5 gpc1300 (
      {stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_14[107]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[38],stage2_15[44],stage2_14[61],stage2_13[76]}
   );
   gpc615_5 gpc1301 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166]},
      {stage1_14[108]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage2_17[22],stage2_16[39],stage2_15[45],stage2_14[62],stage2_13[77]}
   );
   gpc615_5 gpc1302 (
      {stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171]},
      {stage1_14[109]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage2_17[23],stage2_16[40],stage2_15[46],stage2_14[63],stage2_13[78]}
   );
   gpc615_5 gpc1303 (
      {stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage1_14[110]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage2_17[24],stage2_16[41],stage2_15[47],stage2_14[64],stage2_13[79]}
   );
   gpc615_5 gpc1304 (
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181]},
      {stage1_14[111]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage2_17[25],stage2_16[42],stage2_15[48],stage2_14[65],stage2_13[80]}
   );
   gpc615_5 gpc1305 (
      {stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185], stage1_13[186]},
      {stage1_14[112]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage2_17[26],stage2_16[43],stage2_15[49],stage2_14[66],stage2_13[81]}
   );
   gpc615_5 gpc1306 (
      {stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_14[113]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage2_17[27],stage2_16[44],stage2_15[50],stage2_14[67],stage2_13[82]}
   );
   gpc615_5 gpc1307 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196]},
      {stage1_14[114]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage2_17[28],stage2_16[45],stage2_15[51],stage2_14[68],stage2_13[83]}
   );
   gpc615_5 gpc1308 (
      {stage1_13[197], stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201]},
      {stage1_14[115]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage2_17[29],stage2_16[46],stage2_15[52],stage2_14[69],stage2_13[84]}
   );
   gpc615_5 gpc1309 (
      {stage1_13[202], stage1_13[203], stage1_13[204], stage1_13[205], stage1_13[206]},
      {stage1_14[116]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage2_17[30],stage2_16[47],stage2_15[53],stage2_14[70],stage2_13[85]}
   );
   gpc615_5 gpc1310 (
      {stage1_13[207], stage1_13[208], stage1_13[209], stage1_13[210], stage1_13[211]},
      {stage1_14[117]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage2_17[31],stage2_16[48],stage2_15[54],stage2_14[71],stage2_13[86]}
   );
   gpc615_5 gpc1311 (
      {stage1_13[212], stage1_13[213], stage1_13[214], stage1_13[215], stage1_13[216]},
      {stage1_14[118]},
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196], stage1_15[197]},
      {stage2_17[32],stage2_16[49],stage2_15[55],stage2_14[72],stage2_13[87]}
   );
   gpc615_5 gpc1312 (
      {stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_14[119]},
      {stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201], stage1_15[202], stage1_15[203]},
      {stage2_17[33],stage2_16[50],stage2_15[56],stage2_14[73],stage2_13[88]}
   );
   gpc615_5 gpc1313 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226]},
      {stage1_14[120]},
      {stage1_15[204], stage1_15[205], stage1_15[206], stage1_15[207], stage1_15[208], stage1_15[209]},
      {stage2_17[34],stage2_16[51],stage2_15[57],stage2_14[74],stage2_13[89]}
   );
   gpc615_5 gpc1314 (
      {stage1_13[227], stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231]},
      {stage1_14[121]},
      {stage1_15[210], stage1_15[211], stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215]},
      {stage2_17[35],stage2_16[52],stage2_15[58],stage2_14[75],stage2_13[90]}
   );
   gpc606_5 gpc1315 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[36],stage2_16[53],stage2_15[59],stage2_14[76]}
   );
   gpc606_5 gpc1316 (
      {stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[37],stage2_16[54],stage2_15[60],stage2_14[77]}
   );
   gpc606_5 gpc1317 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[38],stage2_16[55],stage2_15[61],stage2_14[78]}
   );
   gpc606_5 gpc1318 (
      {stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[39],stage2_16[56],stage2_15[62],stage2_14[79]}
   );
   gpc606_5 gpc1319 (
      {stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[40],stage2_16[57],stage2_15[63],stage2_14[80]}
   );
   gpc606_5 gpc1320 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[41],stage2_16[58],stage2_15[64],stage2_14[81]}
   );
   gpc606_5 gpc1321 (
      {stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[42],stage2_16[59],stage2_15[65],stage2_14[82]}
   );
   gpc606_5 gpc1322 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[43],stage2_16[60],stage2_15[66],stage2_14[83]}
   );
   gpc606_5 gpc1323 (
      {stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[44],stage2_16[61],stage2_15[67],stage2_14[84]}
   );
   gpc606_5 gpc1324 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[45],stage2_16[62],stage2_15[68],stage2_14[85]}
   );
   gpc606_5 gpc1325 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186], stage1_14[187]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[46],stage2_16[63],stage2_15[69],stage2_14[86]}
   );
   gpc606_5 gpc1326 (
      {stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191], stage1_14[192], stage1_14[193]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[47],stage2_16[64],stage2_15[70],stage2_14[87]}
   );
   gpc606_5 gpc1327 (
      {stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[48],stage2_16[65],stage2_15[71],stage2_14[88]}
   );
   gpc606_5 gpc1328 (
      {stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[49],stage2_16[66],stage2_15[72],stage2_14[89]}
   );
   gpc615_5 gpc1329 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[216]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[50],stage2_16[67],stage2_15[73],stage2_14[90]}
   );
   gpc615_5 gpc1330 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[90]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[15],stage2_17[51],stage2_16[68],stage2_15[74]}
   );
   gpc615_5 gpc1331 (
      {stage1_15[222], stage1_15[223], stage1_15[224], stage1_15[225], stage1_15[226]},
      {stage1_16[91]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[16],stage2_17[52],stage2_16[69],stage2_15[75]}
   );
   gpc615_5 gpc1332 (
      {stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230], stage1_15[231]},
      {stage1_16[92]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[17],stage2_17[53],stage2_16[70],stage2_15[76]}
   );
   gpc615_5 gpc1333 (
      {stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_16[93]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[18],stage2_17[54],stage2_16[71],stage2_15[77]}
   );
   gpc615_5 gpc1334 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241]},
      {stage1_16[94]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[19],stage2_17[55],stage2_16[72],stage2_15[78]}
   );
   gpc615_5 gpc1335 (
      {stage1_15[242], stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246]},
      {stage1_16[95]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[20],stage2_17[56],stage2_16[73],stage2_15[79]}
   );
   gpc615_5 gpc1336 (
      {stage1_15[247], stage1_15[248], stage1_15[249], stage1_15[250], stage1_15[251]},
      {stage1_16[96]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[21],stage2_17[57],stage2_16[74],stage2_15[80]}
   );
   gpc615_5 gpc1337 (
      {stage1_15[252], stage1_15[253], stage1_15[254], stage1_15[255], stage1_15[256]},
      {stage1_16[97]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[22],stage2_17[58],stage2_16[75],stage2_15[81]}
   );
   gpc615_5 gpc1338 (
      {stage1_15[257], stage1_15[258], stage1_15[259], stage1_15[260], stage1_15[261]},
      {stage1_16[98]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[23],stage2_17[59],stage2_16[76],stage2_15[82]}
   );
   gpc615_5 gpc1339 (
      {stage1_15[262], stage1_15[263], stage1_15[264], stage1_15[265], stage1_15[266]},
      {stage1_16[99]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[24],stage2_17[60],stage2_16[77],stage2_15[83]}
   );
   gpc615_5 gpc1340 (
      {stage1_15[267], stage1_15[268], stage1_15[269], stage1_15[270], stage1_15[271]},
      {stage1_16[100]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], 1'b0, 1'b0},
      {stage2_19[10],stage2_18[25],stage2_17[61],stage2_16[78],stage2_15[84]}
   );
   gpc1_1 gpc1341 (
      {stage1_3[219]},
      {stage2_3[76]}
   );
   gpc1_1 gpc1342 (
      {stage1_3[220]},
      {stage2_3[77]}
   );
   gpc1_1 gpc1343 (
      {stage1_3[221]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1344 (
      {stage1_3[222]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1345 (
      {stage1_3[223]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1346 (
      {stage1_3[224]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1347 (
      {stage1_3[225]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1348 (
      {stage1_3[226]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1349 (
      {stage1_3[227]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1350 (
      {stage1_3[228]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1351 (
      {stage1_3[229]},
      {stage2_3[86]}
   );
   gpc1_1 gpc1352 (
      {stage1_3[230]},
      {stage2_3[87]}
   );
   gpc1_1 gpc1353 (
      {stage1_3[231]},
      {stage2_3[88]}
   );
   gpc1_1 gpc1354 (
      {stage1_3[232]},
      {stage2_3[89]}
   );
   gpc1_1 gpc1355 (
      {stage1_3[233]},
      {stage2_3[90]}
   );
   gpc1_1 gpc1356 (
      {stage1_3[234]},
      {stage2_3[91]}
   );
   gpc1_1 gpc1357 (
      {stage1_3[235]},
      {stage2_3[92]}
   );
   gpc1_1 gpc1358 (
      {stage1_3[236]},
      {stage2_3[93]}
   );
   gpc1_1 gpc1359 (
      {stage1_3[237]},
      {stage2_3[94]}
   );
   gpc1_1 gpc1360 (
      {stage1_3[238]},
      {stage2_3[95]}
   );
   gpc1_1 gpc1361 (
      {stage1_3[239]},
      {stage2_3[96]}
   );
   gpc1_1 gpc1362 (
      {stage1_3[240]},
      {stage2_3[97]}
   );
   gpc1_1 gpc1363 (
      {stage1_3[241]},
      {stage2_3[98]}
   );
   gpc1_1 gpc1364 (
      {stage1_3[242]},
      {stage2_3[99]}
   );
   gpc1_1 gpc1365 (
      {stage1_3[243]},
      {stage2_3[100]}
   );
   gpc1_1 gpc1366 (
      {stage1_3[244]},
      {stage2_3[101]}
   );
   gpc1_1 gpc1367 (
      {stage1_3[245]},
      {stage2_3[102]}
   );
   gpc1_1 gpc1368 (
      {stage1_4[214]},
      {stage2_4[90]}
   );
   gpc1_1 gpc1369 (
      {stage1_4[215]},
      {stage2_4[91]}
   );
   gpc1_1 gpc1370 (
      {stage1_4[216]},
      {stage2_4[92]}
   );
   gpc1_1 gpc1371 (
      {stage1_4[217]},
      {stage2_4[93]}
   );
   gpc1_1 gpc1372 (
      {stage1_4[218]},
      {stage2_4[94]}
   );
   gpc1_1 gpc1373 (
      {stage1_4[219]},
      {stage2_4[95]}
   );
   gpc1_1 gpc1374 (
      {stage1_4[220]},
      {stage2_4[96]}
   );
   gpc1_1 gpc1375 (
      {stage1_4[221]},
      {stage2_4[97]}
   );
   gpc1_1 gpc1376 (
      {stage1_4[222]},
      {stage2_4[98]}
   );
   gpc1_1 gpc1377 (
      {stage1_4[223]},
      {stage2_4[99]}
   );
   gpc1_1 gpc1378 (
      {stage1_4[224]},
      {stage2_4[100]}
   );
   gpc1_1 gpc1379 (
      {stage1_4[225]},
      {stage2_4[101]}
   );
   gpc1_1 gpc1380 (
      {stage1_4[226]},
      {stage2_4[102]}
   );
   gpc1_1 gpc1381 (
      {stage1_4[227]},
      {stage2_4[103]}
   );
   gpc1_1 gpc1382 (
      {stage1_4[228]},
      {stage2_4[104]}
   );
   gpc1_1 gpc1383 (
      {stage1_4[229]},
      {stage2_4[105]}
   );
   gpc1_1 gpc1384 (
      {stage1_4[230]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1385 (
      {stage1_4[231]},
      {stage2_4[107]}
   );
   gpc1_1 gpc1386 (
      {stage1_4[232]},
      {stage2_4[108]}
   );
   gpc1_1 gpc1387 (
      {stage1_4[233]},
      {stage2_4[109]}
   );
   gpc1_1 gpc1388 (
      {stage1_4[234]},
      {stage2_4[110]}
   );
   gpc1_1 gpc1389 (
      {stage1_4[235]},
      {stage2_4[111]}
   );
   gpc1_1 gpc1390 (
      {stage1_4[236]},
      {stage2_4[112]}
   );
   gpc1_1 gpc1391 (
      {stage1_4[237]},
      {stage2_4[113]}
   );
   gpc1_1 gpc1392 (
      {stage1_4[238]},
      {stage2_4[114]}
   );
   gpc1_1 gpc1393 (
      {stage1_4[239]},
      {stage2_4[115]}
   );
   gpc1_1 gpc1394 (
      {stage1_4[240]},
      {stage2_4[116]}
   );
   gpc1_1 gpc1395 (
      {stage1_5[210]},
      {stage2_5[86]}
   );
   gpc1_1 gpc1396 (
      {stage1_5[211]},
      {stage2_5[87]}
   );
   gpc1_1 gpc1397 (
      {stage1_5[212]},
      {stage2_5[88]}
   );
   gpc1_1 gpc1398 (
      {stage1_5[213]},
      {stage2_5[89]}
   );
   gpc1_1 gpc1399 (
      {stage1_5[214]},
      {stage2_5[90]}
   );
   gpc1_1 gpc1400 (
      {stage1_5[215]},
      {stage2_5[91]}
   );
   gpc1_1 gpc1401 (
      {stage1_5[216]},
      {stage2_5[92]}
   );
   gpc1_1 gpc1402 (
      {stage1_5[217]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1403 (
      {stage1_6[189]},
      {stage2_6[86]}
   );
   gpc1_1 gpc1404 (
      {stage1_6[190]},
      {stage2_6[87]}
   );
   gpc1_1 gpc1405 (
      {stage1_6[191]},
      {stage2_6[88]}
   );
   gpc1_1 gpc1406 (
      {stage1_6[192]},
      {stage2_6[89]}
   );
   gpc1_1 gpc1407 (
      {stage1_6[193]},
      {stage2_6[90]}
   );
   gpc1_1 gpc1408 (
      {stage1_6[194]},
      {stage2_6[91]}
   );
   gpc1_1 gpc1409 (
      {stage1_6[195]},
      {stage2_6[92]}
   );
   gpc1_1 gpc1410 (
      {stage1_6[196]},
      {stage2_6[93]}
   );
   gpc1_1 gpc1411 (
      {stage1_6[197]},
      {stage2_6[94]}
   );
   gpc1_1 gpc1412 (
      {stage1_6[198]},
      {stage2_6[95]}
   );
   gpc1_1 gpc1413 (
      {stage1_6[199]},
      {stage2_6[96]}
   );
   gpc1_1 gpc1414 (
      {stage1_6[200]},
      {stage2_6[97]}
   );
   gpc1_1 gpc1415 (
      {stage1_6[201]},
      {stage2_6[98]}
   );
   gpc1_1 gpc1416 (
      {stage1_6[202]},
      {stage2_6[99]}
   );
   gpc1_1 gpc1417 (
      {stage1_6[203]},
      {stage2_6[100]}
   );
   gpc1_1 gpc1418 (
      {stage1_6[204]},
      {stage2_6[101]}
   );
   gpc1_1 gpc1419 (
      {stage1_6[205]},
      {stage2_6[102]}
   );
   gpc1_1 gpc1420 (
      {stage1_6[206]},
      {stage2_6[103]}
   );
   gpc1_1 gpc1421 (
      {stage1_9[214]},
      {stage2_9[88]}
   );
   gpc1_1 gpc1422 (
      {stage1_9[215]},
      {stage2_9[89]}
   );
   gpc1_1 gpc1423 (
      {stage1_9[216]},
      {stage2_9[90]}
   );
   gpc1_1 gpc1424 (
      {stage1_9[217]},
      {stage2_9[91]}
   );
   gpc1_1 gpc1425 (
      {stage1_9[218]},
      {stage2_9[92]}
   );
   gpc1_1 gpc1426 (
      {stage1_9[219]},
      {stage2_9[93]}
   );
   gpc1_1 gpc1427 (
      {stage1_9[220]},
      {stage2_9[94]}
   );
   gpc1_1 gpc1428 (
      {stage1_9[221]},
      {stage2_9[95]}
   );
   gpc1_1 gpc1429 (
      {stage1_9[222]},
      {stage2_9[96]}
   );
   gpc1_1 gpc1430 (
      {stage1_9[223]},
      {stage2_9[97]}
   );
   gpc1_1 gpc1431 (
      {stage1_9[224]},
      {stage2_9[98]}
   );
   gpc1_1 gpc1432 (
      {stage1_9[225]},
      {stage2_9[99]}
   );
   gpc1_1 gpc1433 (
      {stage1_9[226]},
      {stage2_9[100]}
   );
   gpc1_1 gpc1434 (
      {stage1_9[227]},
      {stage2_9[101]}
   );
   gpc1_1 gpc1435 (
      {stage1_9[228]},
      {stage2_9[102]}
   );
   gpc1_1 gpc1436 (
      {stage1_9[229]},
      {stage2_9[103]}
   );
   gpc1_1 gpc1437 (
      {stage1_9[230]},
      {stage2_9[104]}
   );
   gpc1_1 gpc1438 (
      {stage1_9[231]},
      {stage2_9[105]}
   );
   gpc1_1 gpc1439 (
      {stage1_9[232]},
      {stage2_9[106]}
   );
   gpc1_1 gpc1440 (
      {stage1_9[233]},
      {stage2_9[107]}
   );
   gpc1_1 gpc1441 (
      {stage1_9[234]},
      {stage2_9[108]}
   );
   gpc1_1 gpc1442 (
      {stage1_9[235]},
      {stage2_9[109]}
   );
   gpc1_1 gpc1443 (
      {stage1_9[236]},
      {stage2_9[110]}
   );
   gpc1_1 gpc1444 (
      {stage1_9[237]},
      {stage2_9[111]}
   );
   gpc1_1 gpc1445 (
      {stage1_9[238]},
      {stage2_9[112]}
   );
   gpc1_1 gpc1446 (
      {stage1_9[239]},
      {stage2_9[113]}
   );
   gpc1_1 gpc1447 (
      {stage1_9[240]},
      {stage2_9[114]}
   );
   gpc1_1 gpc1448 (
      {stage1_9[241]},
      {stage2_9[115]}
   );
   gpc1_1 gpc1449 (
      {stage1_9[242]},
      {stage2_9[116]}
   );
   gpc1_1 gpc1450 (
      {stage1_9[243]},
      {stage2_9[117]}
   );
   gpc1_1 gpc1451 (
      {stage1_9[244]},
      {stage2_9[118]}
   );
   gpc1_1 gpc1452 (
      {stage1_9[245]},
      {stage2_9[119]}
   );
   gpc1_1 gpc1453 (
      {stage1_9[246]},
      {stage2_9[120]}
   );
   gpc1_1 gpc1454 (
      {stage1_9[247]},
      {stage2_9[121]}
   );
   gpc1_1 gpc1455 (
      {stage1_9[248]},
      {stage2_9[122]}
   );
   gpc1_1 gpc1456 (
      {stage1_9[249]},
      {stage2_9[123]}
   );
   gpc1_1 gpc1457 (
      {stage1_9[250]},
      {stage2_9[124]}
   );
   gpc1_1 gpc1458 (
      {stage1_9[251]},
      {stage2_9[125]}
   );
   gpc1_1 gpc1459 (
      {stage1_9[252]},
      {stage2_9[126]}
   );
   gpc1_1 gpc1460 (
      {stage1_9[253]},
      {stage2_9[127]}
   );
   gpc1_1 gpc1461 (
      {stage1_9[254]},
      {stage2_9[128]}
   );
   gpc1_1 gpc1462 (
      {stage1_9[255]},
      {stage2_9[129]}
   );
   gpc1_1 gpc1463 (
      {stage1_9[256]},
      {stage2_9[130]}
   );
   gpc1_1 gpc1464 (
      {stage1_9[257]},
      {stage2_9[131]}
   );
   gpc1_1 gpc1465 (
      {stage1_9[258]},
      {stage2_9[132]}
   );
   gpc1_1 gpc1466 (
      {stage1_9[259]},
      {stage2_9[133]}
   );
   gpc1_1 gpc1467 (
      {stage1_9[260]},
      {stage2_9[134]}
   );
   gpc1_1 gpc1468 (
      {stage1_9[261]},
      {stage2_9[135]}
   );
   gpc1_1 gpc1469 (
      {stage1_9[262]},
      {stage2_9[136]}
   );
   gpc1_1 gpc1470 (
      {stage1_9[263]},
      {stage2_9[137]}
   );
   gpc1_1 gpc1471 (
      {stage1_11[120]},
      {stage2_11[74]}
   );
   gpc1_1 gpc1472 (
      {stage1_11[121]},
      {stage2_11[75]}
   );
   gpc1_1 gpc1473 (
      {stage1_11[122]},
      {stage2_11[76]}
   );
   gpc1_1 gpc1474 (
      {stage1_11[123]},
      {stage2_11[77]}
   );
   gpc1_1 gpc1475 (
      {stage1_11[124]},
      {stage2_11[78]}
   );
   gpc1_1 gpc1476 (
      {stage1_11[125]},
      {stage2_11[79]}
   );
   gpc1_1 gpc1477 (
      {stage1_11[126]},
      {stage2_11[80]}
   );
   gpc1_1 gpc1478 (
      {stage1_11[127]},
      {stage2_11[81]}
   );
   gpc1_1 gpc1479 (
      {stage1_11[128]},
      {stage2_11[82]}
   );
   gpc1_1 gpc1480 (
      {stage1_11[129]},
      {stage2_11[83]}
   );
   gpc1_1 gpc1481 (
      {stage1_11[130]},
      {stage2_11[84]}
   );
   gpc1_1 gpc1482 (
      {stage1_11[131]},
      {stage2_11[85]}
   );
   gpc1_1 gpc1483 (
      {stage1_11[132]},
      {stage2_11[86]}
   );
   gpc1_1 gpc1484 (
      {stage1_11[133]},
      {stage2_11[87]}
   );
   gpc1_1 gpc1485 (
      {stage1_11[134]},
      {stage2_11[88]}
   );
   gpc1_1 gpc1486 (
      {stage1_11[135]},
      {stage2_11[89]}
   );
   gpc1_1 gpc1487 (
      {stage1_11[136]},
      {stage2_11[90]}
   );
   gpc1_1 gpc1488 (
      {stage1_11[137]},
      {stage2_11[91]}
   );
   gpc1_1 gpc1489 (
      {stage1_11[138]},
      {stage2_11[92]}
   );
   gpc1_1 gpc1490 (
      {stage1_11[139]},
      {stage2_11[93]}
   );
   gpc1_1 gpc1491 (
      {stage1_11[140]},
      {stage2_11[94]}
   );
   gpc1_1 gpc1492 (
      {stage1_11[141]},
      {stage2_11[95]}
   );
   gpc1_1 gpc1493 (
      {stage1_11[142]},
      {stage2_11[96]}
   );
   gpc1_1 gpc1494 (
      {stage1_11[143]},
      {stage2_11[97]}
   );
   gpc1_1 gpc1495 (
      {stage1_11[144]},
      {stage2_11[98]}
   );
   gpc1_1 gpc1496 (
      {stage1_11[145]},
      {stage2_11[99]}
   );
   gpc1_1 gpc1497 (
      {stage1_11[146]},
      {stage2_11[100]}
   );
   gpc1_1 gpc1498 (
      {stage1_11[147]},
      {stage2_11[101]}
   );
   gpc1_1 gpc1499 (
      {stage1_11[148]},
      {stage2_11[102]}
   );
   gpc1_1 gpc1500 (
      {stage1_11[149]},
      {stage2_11[103]}
   );
   gpc1_1 gpc1501 (
      {stage1_11[150]},
      {stage2_11[104]}
   );
   gpc1_1 gpc1502 (
      {stage1_11[151]},
      {stage2_11[105]}
   );
   gpc1_1 gpc1503 (
      {stage1_11[152]},
      {stage2_11[106]}
   );
   gpc1_1 gpc1504 (
      {stage1_11[153]},
      {stage2_11[107]}
   );
   gpc1_1 gpc1505 (
      {stage1_11[154]},
      {stage2_11[108]}
   );
   gpc1_1 gpc1506 (
      {stage1_11[155]},
      {stage2_11[109]}
   );
   gpc1_1 gpc1507 (
      {stage1_11[156]},
      {stage2_11[110]}
   );
   gpc1_1 gpc1508 (
      {stage1_11[157]},
      {stage2_11[111]}
   );
   gpc1_1 gpc1509 (
      {stage1_11[158]},
      {stage2_11[112]}
   );
   gpc1_1 gpc1510 (
      {stage1_11[159]},
      {stage2_11[113]}
   );
   gpc1_1 gpc1511 (
      {stage1_11[160]},
      {stage2_11[114]}
   );
   gpc1_1 gpc1512 (
      {stage1_11[161]},
      {stage2_11[115]}
   );
   gpc1_1 gpc1513 (
      {stage1_11[162]},
      {stage2_11[116]}
   );
   gpc1_1 gpc1514 (
      {stage1_11[163]},
      {stage2_11[117]}
   );
   gpc1_1 gpc1515 (
      {stage1_11[164]},
      {stage2_11[118]}
   );
   gpc1_1 gpc1516 (
      {stage1_11[165]},
      {stage2_11[119]}
   );
   gpc1_1 gpc1517 (
      {stage1_11[166]},
      {stage2_11[120]}
   );
   gpc1_1 gpc1518 (
      {stage1_11[167]},
      {stage2_11[121]}
   );
   gpc1_1 gpc1519 (
      {stage1_11[168]},
      {stage2_11[122]}
   );
   gpc1_1 gpc1520 (
      {stage1_11[169]},
      {stage2_11[123]}
   );
   gpc1_1 gpc1521 (
      {stage1_11[170]},
      {stage2_11[124]}
   );
   gpc1_1 gpc1522 (
      {stage1_11[171]},
      {stage2_11[125]}
   );
   gpc1_1 gpc1523 (
      {stage1_11[172]},
      {stage2_11[126]}
   );
   gpc1_1 gpc1524 (
      {stage1_11[173]},
      {stage2_11[127]}
   );
   gpc1_1 gpc1525 (
      {stage1_11[174]},
      {stage2_11[128]}
   );
   gpc1_1 gpc1526 (
      {stage1_11[175]},
      {stage2_11[129]}
   );
   gpc1_1 gpc1527 (
      {stage1_11[176]},
      {stage2_11[130]}
   );
   gpc1_1 gpc1528 (
      {stage1_11[177]},
      {stage2_11[131]}
   );
   gpc1_1 gpc1529 (
      {stage1_11[178]},
      {stage2_11[132]}
   );
   gpc1_1 gpc1530 (
      {stage1_11[179]},
      {stage2_11[133]}
   );
   gpc1_1 gpc1531 (
      {stage1_11[180]},
      {stage2_11[134]}
   );
   gpc1_1 gpc1532 (
      {stage1_11[181]},
      {stage2_11[135]}
   );
   gpc1_1 gpc1533 (
      {stage1_11[182]},
      {stage2_11[136]}
   );
   gpc1_1 gpc1534 (
      {stage1_11[183]},
      {stage2_11[137]}
   );
   gpc1_1 gpc1535 (
      {stage1_11[184]},
      {stage2_11[138]}
   );
   gpc1_1 gpc1536 (
      {stage1_11[185]},
      {stage2_11[139]}
   );
   gpc1_1 gpc1537 (
      {stage1_11[186]},
      {stage2_11[140]}
   );
   gpc1_1 gpc1538 (
      {stage1_11[187]},
      {stage2_11[141]}
   );
   gpc1_1 gpc1539 (
      {stage1_11[188]},
      {stage2_11[142]}
   );
   gpc1_1 gpc1540 (
      {stage1_11[189]},
      {stage2_11[143]}
   );
   gpc1_1 gpc1541 (
      {stage1_12[210]},
      {stage2_12[73]}
   );
   gpc1_1 gpc1542 (
      {stage1_12[211]},
      {stage2_12[74]}
   );
   gpc1_1 gpc1543 (
      {stage1_12[212]},
      {stage2_12[75]}
   );
   gpc1_1 gpc1544 (
      {stage1_12[213]},
      {stage2_12[76]}
   );
   gpc1_1 gpc1545 (
      {stage1_12[214]},
      {stage2_12[77]}
   );
   gpc1_1 gpc1546 (
      {stage1_12[215]},
      {stage2_12[78]}
   );
   gpc1_1 gpc1547 (
      {stage1_12[216]},
      {stage2_12[79]}
   );
   gpc1_1 gpc1548 (
      {stage1_12[217]},
      {stage2_12[80]}
   );
   gpc1_1 gpc1549 (
      {stage1_12[218]},
      {stage2_12[81]}
   );
   gpc1_1 gpc1550 (
      {stage1_12[219]},
      {stage2_12[82]}
   );
   gpc1_1 gpc1551 (
      {stage1_12[220]},
      {stage2_12[83]}
   );
   gpc1_1 gpc1552 (
      {stage1_12[221]},
      {stage2_12[84]}
   );
   gpc1_1 gpc1553 (
      {stage1_13[232]},
      {stage2_13[91]}
   );
   gpc1_1 gpc1554 (
      {stage1_13[233]},
      {stage2_13[92]}
   );
   gpc1_1 gpc1555 (
      {stage1_13[234]},
      {stage2_13[93]}
   );
   gpc1_1 gpc1556 (
      {stage1_13[235]},
      {stage2_13[94]}
   );
   gpc1_1 gpc1557 (
      {stage1_13[236]},
      {stage2_13[95]}
   );
   gpc1_1 gpc1558 (
      {stage1_13[237]},
      {stage2_13[96]}
   );
   gpc1_1 gpc1559 (
      {stage1_13[238]},
      {stage2_13[97]}
   );
   gpc1_1 gpc1560 (
      {stage1_13[239]},
      {stage2_13[98]}
   );
   gpc1_1 gpc1561 (
      {stage1_13[240]},
      {stage2_13[99]}
   );
   gpc1_1 gpc1562 (
      {stage1_13[241]},
      {stage2_13[100]}
   );
   gpc1_1 gpc1563 (
      {stage1_13[242]},
      {stage2_13[101]}
   );
   gpc1_1 gpc1564 (
      {stage1_13[243]},
      {stage2_13[102]}
   );
   gpc1_1 gpc1565 (
      {stage1_13[244]},
      {stage2_13[103]}
   );
   gpc1_1 gpc1566 (
      {stage1_13[245]},
      {stage2_13[104]}
   );
   gpc1_1 gpc1567 (
      {stage1_13[246]},
      {stage2_13[105]}
   );
   gpc1_1 gpc1568 (
      {stage1_13[247]},
      {stage2_13[106]}
   );
   gpc1_1 gpc1569 (
      {stage1_13[248]},
      {stage2_13[107]}
   );
   gpc1_1 gpc1570 (
      {stage1_13[249]},
      {stage2_13[108]}
   );
   gpc1_1 gpc1571 (
      {stage1_13[250]},
      {stage2_13[109]}
   );
   gpc1_1 gpc1572 (
      {stage1_13[251]},
      {stage2_13[110]}
   );
   gpc1_1 gpc1573 (
      {stage1_13[252]},
      {stage2_13[111]}
   );
   gpc1_1 gpc1574 (
      {stage1_13[253]},
      {stage2_13[112]}
   );
   gpc1_1 gpc1575 (
      {stage1_13[254]},
      {stage2_13[113]}
   );
   gpc1_1 gpc1576 (
      {stage1_13[255]},
      {stage2_13[114]}
   );
   gpc1_1 gpc1577 (
      {stage1_13[256]},
      {stage2_13[115]}
   );
   gpc1_1 gpc1578 (
      {stage1_13[257]},
      {stage2_13[116]}
   );
   gpc1_1 gpc1579 (
      {stage1_13[258]},
      {stage2_13[117]}
   );
   gpc1_1 gpc1580 (
      {stage1_13[259]},
      {stage2_13[118]}
   );
   gpc1_1 gpc1581 (
      {stage1_13[260]},
      {stage2_13[119]}
   );
   gpc1_1 gpc1582 (
      {stage1_13[261]},
      {stage2_13[120]}
   );
   gpc1_1 gpc1583 (
      {stage1_13[262]},
      {stage2_13[121]}
   );
   gpc1_1 gpc1584 (
      {stage1_13[263]},
      {stage2_13[122]}
   );
   gpc1_1 gpc1585 (
      {stage1_13[264]},
      {stage2_13[123]}
   );
   gpc1_1 gpc1586 (
      {stage1_13[265]},
      {stage2_13[124]}
   );
   gpc1_1 gpc1587 (
      {stage1_13[266]},
      {stage2_13[125]}
   );
   gpc1_1 gpc1588 (
      {stage1_13[267]},
      {stage2_13[126]}
   );
   gpc1_1 gpc1589 (
      {stage1_13[268]},
      {stage2_13[127]}
   );
   gpc1_1 gpc1590 (
      {stage1_13[269]},
      {stage2_13[128]}
   );
   gpc1_1 gpc1591 (
      {stage1_13[270]},
      {stage2_13[129]}
   );
   gpc1_1 gpc1592 (
      {stage1_13[271]},
      {stage2_13[130]}
   );
   gpc1_1 gpc1593 (
      {stage1_13[272]},
      {stage2_13[131]}
   );
   gpc1_1 gpc1594 (
      {stage1_13[273]},
      {stage2_13[132]}
   );
   gpc1_1 gpc1595 (
      {stage1_13[274]},
      {stage2_13[133]}
   );
   gpc1_1 gpc1596 (
      {stage1_13[275]},
      {stage2_13[134]}
   );
   gpc1_1 gpc1597 (
      {stage1_13[276]},
      {stage2_13[135]}
   );
   gpc1_1 gpc1598 (
      {stage1_13[277]},
      {stage2_13[136]}
   );
   gpc1_1 gpc1599 (
      {stage1_13[278]},
      {stage2_13[137]}
   );
   gpc1_1 gpc1600 (
      {stage1_13[279]},
      {stage2_13[138]}
   );
   gpc1_1 gpc1601 (
      {stage1_13[280]},
      {stage2_13[139]}
   );
   gpc1_1 gpc1602 (
      {stage1_13[281]},
      {stage2_13[140]}
   );
   gpc1_1 gpc1603 (
      {stage1_14[211]},
      {stage2_14[91]}
   );
   gpc1_1 gpc1604 (
      {stage1_14[212]},
      {stage2_14[92]}
   );
   gpc1_1 gpc1605 (
      {stage1_14[213]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1606 (
      {stage1_14[214]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1607 (
      {stage1_14[215]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1608 (
      {stage1_14[216]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1609 (
      {stage1_14[217]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1610 (
      {stage1_14[218]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1611 (
      {stage1_14[219]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1612 (
      {stage1_14[220]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1613 (
      {stage1_14[221]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1614 (
      {stage1_14[222]},
      {stage2_14[102]}
   );
   gpc1_1 gpc1615 (
      {stage1_14[223]},
      {stage2_14[103]}
   );
   gpc1_1 gpc1616 (
      {stage1_14[224]},
      {stage2_14[104]}
   );
   gpc1_1 gpc1617 (
      {stage1_14[225]},
      {stage2_14[105]}
   );
   gpc1_1 gpc1618 (
      {stage1_14[226]},
      {stage2_14[106]}
   );
   gpc1_1 gpc1619 (
      {stage1_14[227]},
      {stage2_14[107]}
   );
   gpc1_1 gpc1620 (
      {stage1_14[228]},
      {stage2_14[108]}
   );
   gpc1_1 gpc1621 (
      {stage1_14[229]},
      {stage2_14[109]}
   );
   gpc1_1 gpc1622 (
      {stage1_14[230]},
      {stage2_14[110]}
   );
   gpc1_1 gpc1623 (
      {stage1_14[231]},
      {stage2_14[111]}
   );
   gpc1_1 gpc1624 (
      {stage1_14[232]},
      {stage2_14[112]}
   );
   gpc1_1 gpc1625 (
      {stage1_14[233]},
      {stage2_14[113]}
   );
   gpc1_1 gpc1626 (
      {stage1_14[234]},
      {stage2_14[114]}
   );
   gpc1_1 gpc1627 (
      {stage1_14[235]},
      {stage2_14[115]}
   );
   gpc1_1 gpc1628 (
      {stage1_14[236]},
      {stage2_14[116]}
   );
   gpc1_1 gpc1629 (
      {stage1_14[237]},
      {stage2_14[117]}
   );
   gpc1_1 gpc1630 (
      {stage1_14[238]},
      {stage2_14[118]}
   );
   gpc1_1 gpc1631 (
      {stage1_14[239]},
      {stage2_14[119]}
   );
   gpc1_1 gpc1632 (
      {stage1_14[240]},
      {stage2_14[120]}
   );
   gpc1_1 gpc1633 (
      {stage1_14[241]},
      {stage2_14[121]}
   );
   gpc1_1 gpc1634 (
      {stage1_14[242]},
      {stage2_14[122]}
   );
   gpc1_1 gpc1635 (
      {stage1_14[243]},
      {stage2_14[123]}
   );
   gpc1_1 gpc1636 (
      {stage1_14[244]},
      {stage2_14[124]}
   );
   gpc1_1 gpc1637 (
      {stage1_16[101]},
      {stage2_16[79]}
   );
   gpc1_1 gpc1638 (
      {stage1_16[102]},
      {stage2_16[80]}
   );
   gpc1_1 gpc1639 (
      {stage1_16[103]},
      {stage2_16[81]}
   );
   gpc1_1 gpc1640 (
      {stage1_16[104]},
      {stage2_16[82]}
   );
   gpc1_1 gpc1641 (
      {stage1_16[105]},
      {stage2_16[83]}
   );
   gpc1_1 gpc1642 (
      {stage1_16[106]},
      {stage2_16[84]}
   );
   gpc1_1 gpc1643 (
      {stage1_16[107]},
      {stage2_16[85]}
   );
   gpc1_1 gpc1644 (
      {stage1_16[108]},
      {stage2_16[86]}
   );
   gpc1_1 gpc1645 (
      {stage1_16[109]},
      {stage2_16[87]}
   );
   gpc1_1 gpc1646 (
      {stage1_16[110]},
      {stage2_16[88]}
   );
   gpc1_1 gpc1647 (
      {stage1_16[111]},
      {stage2_16[89]}
   );
   gpc1_1 gpc1648 (
      {stage1_16[112]},
      {stage2_16[90]}
   );
   gpc1_1 gpc1649 (
      {stage1_16[113]},
      {stage2_16[91]}
   );
   gpc1_1 gpc1650 (
      {stage1_16[114]},
      {stage2_16[92]}
   );
   gpc1_1 gpc1651 (
      {stage1_16[115]},
      {stage2_16[93]}
   );
   gpc1_1 gpc1652 (
      {stage1_16[116]},
      {stage2_16[94]}
   );
   gpc1_1 gpc1653 (
      {stage1_16[117]},
      {stage2_16[95]}
   );
   gpc1_1 gpc1654 (
      {stage1_16[118]},
      {stage2_16[96]}
   );
   gpc1_1 gpc1655 (
      {stage1_16[119]},
      {stage2_16[97]}
   );
   gpc1_1 gpc1656 (
      {stage1_16[120]},
      {stage2_16[98]}
   );
   gpc1_1 gpc1657 (
      {stage1_16[121]},
      {stage2_16[99]}
   );
   gpc1_1 gpc1658 (
      {stage1_16[122]},
      {stage2_16[100]}
   );
   gpc1_1 gpc1659 (
      {stage1_16[123]},
      {stage2_16[101]}
   );
   gpc1_1 gpc1660 (
      {stage1_16[124]},
      {stage2_16[102]}
   );
   gpc1_1 gpc1661 (
      {stage1_16[125]},
      {stage2_16[103]}
   );
   gpc1_1 gpc1662 (
      {stage1_16[126]},
      {stage2_16[104]}
   );
   gpc606_5 gpc1663 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc1664 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_1[0]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc1665 (
      {stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15]},
      {stage2_1[1]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc1666 (
      {stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[2]},
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1667 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc1668 (
      {stage2_1[9], stage2_1[10], stage2_1[11], stage2_1[12], stage2_1[13], stage2_1[14]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc1669 (
      {stage2_1[15], stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1670 (
      {stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24], stage2_1[25], stage2_1[26]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1671 (
      {stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30], stage2_1[31], stage2_1[32]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1672 (
      {stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36], stage2_1[37], stage2_1[38]},
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1673 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc1674 (
      {stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[36]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc1675 (
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38], stage2_2[39]},
      {stage2_3[37]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc1676 (
      {stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_3[38]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc1677 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49]},
      {stage2_3[39]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1678 (
      {stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage2_3[40]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1679 (
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59]},
      {stage2_3[41]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc606_5 gpc1680 (
      {stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc1681 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52]},
      {stage2_4[42]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc1682 (
      {stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57]},
      {stage2_4[43]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1683 (
      {stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62]},
      {stage2_4[44]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1684 (
      {stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67]},
      {stage2_4[45]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1685 (
      {stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage2_4[46]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1686 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[47]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc1687 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[48]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc1688 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[49]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc1689 (
      {stage2_3[88], stage2_3[89], stage2_3[90], stage2_3[91], stage2_3[92]},
      {stage2_4[50]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc1690 (
      {stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96], stage2_3[97]},
      {stage2_4[51]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc1691 (
      {stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102]},
      {stage2_4[52]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc1692 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc1693 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc1694 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[14],stage3_6[21],stage3_5[27],stage3_4[31]}
   );
   gpc606_5 gpc1695 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[15],stage3_6[22],stage3_5[28],stage3_4[32]}
   );
   gpc606_5 gpc1696 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[16],stage3_6[23],stage3_5[29],stage3_4[33]}
   );
   gpc606_5 gpc1697 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[17],stage3_6[24],stage3_5[30],stage3_4[34]}
   );
   gpc606_5 gpc1698 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[18],stage3_6[25],stage3_5[31],stage3_4[35]}
   );
   gpc606_5 gpc1699 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[19],stage3_6[26],stage3_5[32],stage3_4[36]}
   );
   gpc606_5 gpc1700 (
      {stage2_4[101], stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[20],stage3_6[27],stage3_5[33],stage3_4[37]}
   );
   gpc615_5 gpc1701 (
      {stage2_4[107], stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111]},
      {stage2_5[72]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[21],stage3_6[28],stage3_5[34],stage3_4[38]}
   );
   gpc615_5 gpc1702 (
      {stage2_4[112], stage2_4[113], stage2_4[114], stage2_4[115], stage2_4[116]},
      {stage2_5[73]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[22],stage3_6[29],stage3_5[35],stage3_4[39]}
   );
   gpc615_5 gpc1703 (
      {stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77], stage2_5[78]},
      {stage2_6[66]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[11],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc615_5 gpc1704 (
      {stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_6[67]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[12],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1705 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[13],stage3_7[25],stage3_6[32]}
   );
   gpc606_5 gpc1706 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78], stage2_6[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[14],stage3_7[26],stage3_6[33]}
   );
   gpc606_5 gpc1707 (
      {stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83], stage2_6[84], stage2_6[85]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[15],stage3_7[27],stage3_6[34]}
   );
   gpc606_5 gpc1708 (
      {stage2_6[86], stage2_6[87], stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[5],stage3_8[16],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc1709 (
      {stage2_6[92], stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[6],stage3_8[17],stage3_7[29],stage3_6[36]}
   );
   gpc606_5 gpc1710 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102], stage2_6[103]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[7],stage3_8[18],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1711 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[8],stage3_8[19],stage3_7[31]}
   );
   gpc615_5 gpc1712 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[9],stage3_8[20],stage3_7[32]}
   );
   gpc615_5 gpc1713 (
      {stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[10],stage3_8[21],stage3_7[33]}
   );
   gpc615_5 gpc1714 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[11],stage3_8[22],stage3_7[34]}
   );
   gpc615_5 gpc1715 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[40]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[10],stage3_9[12],stage3_8[23],stage3_7[35]}
   );
   gpc615_5 gpc1716 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[41]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[11],stage3_9[13],stage3_8[24],stage3_7[36]}
   );
   gpc615_5 gpc1717 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[42]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[12],stage3_9[14],stage3_8[25],stage3_7[37]}
   );
   gpc615_5 gpc1718 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[43]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[13],stage3_9[15],stage3_8[26],stage3_7[38]}
   );
   gpc615_5 gpc1719 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[44]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[14],stage3_9[16],stage3_8[27],stage3_7[39]}
   );
   gpc615_5 gpc1720 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[45]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[15],stage3_9[17],stage3_8[28],stage3_7[40]}
   );
   gpc615_5 gpc1721 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[46]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[16],stage3_9[18],stage3_8[29],stage3_7[41]}
   );
   gpc615_5 gpc1722 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[47]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[17],stage3_9[19],stage3_8[30],stage3_7[42]}
   );
   gpc615_5 gpc1723 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[48]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[18],stage3_9[20],stage3_8[31],stage3_7[43]}
   );
   gpc615_5 gpc1724 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[49]},
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage3_11[13],stage3_10[19],stage3_9[21],stage3_8[32],stage3_7[44]}
   );
   gpc615_5 gpc1725 (
      {stage2_7[82], stage2_7[83], stage2_7[84], 1'b0, 1'b0},
      {stage2_8[50]},
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage3_11[14],stage3_10[20],stage3_9[22],stage3_8[33],stage3_7[45]}
   );
   gpc606_5 gpc1726 (
      {stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[15],stage3_10[21],stage3_9[23],stage3_8[34]}
   );
   gpc615_5 gpc1727 (
      {stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61]},
      {stage2_9[90]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[16],stage3_10[22],stage3_9[24],stage3_8[35]}
   );
   gpc615_5 gpc1728 (
      {stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65], stage2_8[66]},
      {stage2_9[91]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[17],stage3_10[23],stage3_9[25],stage3_8[36]}
   );
   gpc615_5 gpc1729 (
      {stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_9[92]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[18],stage3_10[24],stage3_9[26],stage3_8[37]}
   );
   gpc615_5 gpc1730 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_9[93]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[19],stage3_10[25],stage3_9[27],stage3_8[38]}
   );
   gpc615_5 gpc1731 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_9[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[20],stage3_10[26],stage3_9[28],stage3_8[39]}
   );
   gpc615_5 gpc1732 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86]},
      {stage2_9[95]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[21],stage3_10[27],stage3_9[29],stage3_8[40]}
   );
   gpc606_5 gpc1733 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[22],stage3_10[28],stage3_9[30]}
   );
   gpc606_5 gpc1734 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[8],stage3_11[23],stage3_10[29],stage3_9[31]}
   );
   gpc606_5 gpc1735 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[9],stage3_11[24],stage3_10[30],stage3_9[32]}
   );
   gpc606_5 gpc1736 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[10],stage3_11[25],stage3_10[31],stage3_9[33]}
   );
   gpc615_5 gpc1737 (
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[11],stage3_11[26],stage3_10[32]}
   );
   gpc615_5 gpc1738 (
      {stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51]},
      {stage2_11[25]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[5],stage3_12[12],stage3_11[27],stage3_10[33]}
   );
   gpc615_5 gpc1739 (
      {stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_11[26]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[6],stage3_12[13],stage3_11[28],stage3_10[34]}
   );
   gpc606_5 gpc1740 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[7],stage3_12[14],stage3_11[29]}
   );
   gpc606_5 gpc1741 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[8],stage3_12[15],stage3_11[30]}
   );
   gpc606_5 gpc1742 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[9],stage3_12[16],stage3_11[31]}
   );
   gpc606_5 gpc1743 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[10],stage3_12[17],stage3_11[32]}
   );
   gpc606_5 gpc1744 (
      {stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[11],stage3_12[18],stage3_11[33]}
   );
   gpc606_5 gpc1745 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[12],stage3_12[19],stage3_11[34]}
   );
   gpc606_5 gpc1746 (
      {stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[9],stage3_13[13],stage3_12[20],stage3_11[35]}
   );
   gpc606_5 gpc1747 (
      {stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[10],stage3_13[14],stage3_12[21],stage3_11[36]}
   );
   gpc606_5 gpc1748 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[11],stage3_13[15],stage3_12[22],stage3_11[37]}
   );
   gpc606_5 gpc1749 (
      {stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[12],stage3_13[16],stage3_12[23],stage3_11[38]}
   );
   gpc606_5 gpc1750 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91], stage2_11[92]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[13],stage3_13[17],stage3_12[24],stage3_11[39]}
   );
   gpc606_5 gpc1751 (
      {stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[14],stage3_13[18],stage3_12[25],stage3_11[40]}
   );
   gpc606_5 gpc1752 (
      {stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[15],stage3_13[19],stage3_12[26],stage3_11[41]}
   );
   gpc606_5 gpc1753 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109], stage2_11[110]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[16],stage3_13[20],stage3_12[27],stage3_11[42]}
   );
   gpc606_5 gpc1754 (
      {stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114], stage2_11[115], stage2_11[116]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[17],stage3_13[21],stage3_12[28],stage3_11[43]}
   );
   gpc606_5 gpc1755 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121], stage2_11[122]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[18],stage3_13[22],stage3_12[29],stage3_11[44]}
   );
   gpc606_5 gpc1756 (
      {stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126], stage2_11[127], stage2_11[128]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[19],stage3_13[23],stage3_12[30],stage3_11[45]}
   );
   gpc606_5 gpc1757 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[17],stage3_14[20],stage3_13[24],stage3_12[31]}
   );
   gpc606_5 gpc1758 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[18],stage3_14[21],stage3_13[25],stage3_12[32]}
   );
   gpc606_5 gpc1759 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[19],stage3_14[22],stage3_13[26],stage3_12[33]}
   );
   gpc606_5 gpc1760 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[20],stage3_14[23],stage3_13[27],stage3_12[34]}
   );
   gpc606_5 gpc1761 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[21],stage3_14[24],stage3_13[28],stage3_12[35]}
   );
   gpc606_5 gpc1762 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[22],stage3_14[25],stage3_13[29],stage3_12[36]}
   );
   gpc606_5 gpc1763 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[23],stage3_14[26],stage3_13[30],stage3_12[37]}
   );
   gpc606_5 gpc1764 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[24],stage3_14[27],stage3_13[31],stage3_12[38]}
   );
   gpc606_5 gpc1765 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[25],stage3_14[28],stage3_13[32],stage3_12[39]}
   );
   gpc606_5 gpc1766 (
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[9],stage3_15[26],stage3_14[29],stage3_13[33]}
   );
   gpc606_5 gpc1767 (
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[10],stage3_15[27],stage3_14[30],stage3_13[34]}
   );
   gpc606_5 gpc1768 (
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[11],stage3_15[28],stage3_14[31],stage3_13[35]}
   );
   gpc606_5 gpc1769 (
      {stage2_13[120], stage2_13[121], stage2_13[122], stage2_13[123], stage2_13[124], stage2_13[125]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[12],stage3_15[29],stage3_14[32],stage3_13[36]}
   );
   gpc606_5 gpc1770 (
      {stage2_13[126], stage2_13[127], stage2_13[128], stage2_13[129], stage2_13[130], stage2_13[131]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[13],stage3_15[30],stage3_14[33],stage3_13[37]}
   );
   gpc606_5 gpc1771 (
      {stage2_13[132], stage2_13[133], stage2_13[134], stage2_13[135], stage2_13[136], stage2_13[137]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[14],stage3_15[31],stage3_14[34],stage3_13[38]}
   );
   gpc606_5 gpc1772 (
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[15],stage3_15[32],stage3_14[35]}
   );
   gpc606_5 gpc1773 (
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[16],stage3_15[33],stage3_14[36]}
   );
   gpc606_5 gpc1774 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[17],stage3_15[34],stage3_14[37]}
   );
   gpc606_5 gpc1775 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[18],stage3_15[35],stage3_14[38]}
   );
   gpc606_5 gpc1776 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[19],stage3_15[36],stage3_14[39]}
   );
   gpc606_5 gpc1777 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[20],stage3_15[37],stage3_14[40]}
   );
   gpc606_5 gpc1778 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[21],stage3_15[38],stage3_14[41]}
   );
   gpc606_5 gpc1779 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[13],stage3_16[22],stage3_15[39],stage3_14[42]}
   );
   gpc615_5 gpc1780 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106]},
      {stage2_15[36]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[14],stage3_16[23],stage3_15[40],stage3_14[43]}
   );
   gpc615_5 gpc1781 (
      {stage2_14[107], stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111]},
      {stage2_15[37]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[15],stage3_16[24],stage3_15[41],stage3_14[44]}
   );
   gpc615_5 gpc1782 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[16],stage3_16[25],stage3_15[42]}
   );
   gpc615_5 gpc1783 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[17],stage3_16[26],stage3_15[43]}
   );
   gpc615_5 gpc1784 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[18],stage3_16[27],stage3_15[44]}
   );
   gpc615_5 gpc1785 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[19],stage3_16[28],stage3_15[45]}
   );
   gpc615_5 gpc1786 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[20],stage3_16[29],stage3_15[46]}
   );
   gpc615_5 gpc1787 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[21],stage3_16[30],stage3_15[47]}
   );
   gpc615_5 gpc1788 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[22],stage3_16[31],stage3_15[48]}
   );
   gpc615_5 gpc1789 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[23],stage3_16[32],stage3_15[49]}
   );
   gpc606_5 gpc1790 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[18],stage3_17[24],stage3_16[33]}
   );
   gpc606_5 gpc1791 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[9],stage3_18[19],stage3_17[25],stage3_16[34]}
   );
   gpc606_5 gpc1792 (
      {stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83], stage2_16[84], stage2_16[85]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[10],stage3_18[20],stage3_17[26],stage3_16[35]}
   );
   gpc606_5 gpc1793 (
      {stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89], stage2_16[90], stage2_16[91]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[11],stage3_18[21],stage3_17[27],stage3_16[36]}
   );
   gpc606_5 gpc1794 (
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[4],stage3_19[12],stage3_18[22],stage3_17[28]}
   );
   gpc606_5 gpc1795 (
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], 1'b0},
      {stage3_21[1],stage3_20[5],stage3_19[13],stage3_18[23],stage3_17[29]}
   );
   gpc1_1 gpc1796 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1797 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1798 (
      {stage2_1[39]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1799 (
      {stage2_1[40]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1800 (
      {stage2_5[84]},
      {stage3_5[38]}
   );
   gpc1_1 gpc1801 (
      {stage2_5[85]},
      {stage3_5[39]}
   );
   gpc1_1 gpc1802 (
      {stage2_5[86]},
      {stage3_5[40]}
   );
   gpc1_1 gpc1803 (
      {stage2_5[87]},
      {stage3_5[41]}
   );
   gpc1_1 gpc1804 (
      {stage2_5[88]},
      {stage3_5[42]}
   );
   gpc1_1 gpc1805 (
      {stage2_5[89]},
      {stage3_5[43]}
   );
   gpc1_1 gpc1806 (
      {stage2_5[90]},
      {stage3_5[44]}
   );
   gpc1_1 gpc1807 (
      {stage2_5[91]},
      {stage3_5[45]}
   );
   gpc1_1 gpc1808 (
      {stage2_5[92]},
      {stage3_5[46]}
   );
   gpc1_1 gpc1809 (
      {stage2_5[93]},
      {stage3_5[47]}
   );
   gpc1_1 gpc1810 (
      {stage2_9[120]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_9[121]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_9[122]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_9[123]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_9[124]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_9[125]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_9[126]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1817 (
      {stage2_9[127]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1818 (
      {stage2_9[128]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1819 (
      {stage2_9[129]},
      {stage3_9[43]}
   );
   gpc1_1 gpc1820 (
      {stage2_9[130]},
      {stage3_9[44]}
   );
   gpc1_1 gpc1821 (
      {stage2_9[131]},
      {stage3_9[45]}
   );
   gpc1_1 gpc1822 (
      {stage2_9[132]},
      {stage3_9[46]}
   );
   gpc1_1 gpc1823 (
      {stage2_9[133]},
      {stage3_9[47]}
   );
   gpc1_1 gpc1824 (
      {stage2_9[134]},
      {stage3_9[48]}
   );
   gpc1_1 gpc1825 (
      {stage2_9[135]},
      {stage3_9[49]}
   );
   gpc1_1 gpc1826 (
      {stage2_9[136]},
      {stage3_9[50]}
   );
   gpc1_1 gpc1827 (
      {stage2_9[137]},
      {stage3_9[51]}
   );
   gpc1_1 gpc1828 (
      {stage2_10[57]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1829 (
      {stage2_10[58]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1830 (
      {stage2_10[59]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1831 (
      {stage2_10[60]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1832 (
      {stage2_10[61]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1833 (
      {stage2_10[62]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1834 (
      {stage2_10[63]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1835 (
      {stage2_10[64]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1836 (
      {stage2_10[65]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1837 (
      {stage2_10[66]},
      {stage3_10[44]}
   );
   gpc1_1 gpc1838 (
      {stage2_10[67]},
      {stage3_10[45]}
   );
   gpc1_1 gpc1839 (
      {stage2_10[68]},
      {stage3_10[46]}
   );
   gpc1_1 gpc1840 (
      {stage2_10[69]},
      {stage3_10[47]}
   );
   gpc1_1 gpc1841 (
      {stage2_10[70]},
      {stage3_10[48]}
   );
   gpc1_1 gpc1842 (
      {stage2_10[71]},
      {stage3_10[49]}
   );
   gpc1_1 gpc1843 (
      {stage2_10[72]},
      {stage3_10[50]}
   );
   gpc1_1 gpc1844 (
      {stage2_10[73]},
      {stage3_10[51]}
   );
   gpc1_1 gpc1845 (
      {stage2_10[74]},
      {stage3_10[52]}
   );
   gpc1_1 gpc1846 (
      {stage2_10[75]},
      {stage3_10[53]}
   );
   gpc1_1 gpc1847 (
      {stage2_10[76]},
      {stage3_10[54]}
   );
   gpc1_1 gpc1848 (
      {stage2_10[77]},
      {stage3_10[55]}
   );
   gpc1_1 gpc1849 (
      {stage2_10[78]},
      {stage3_10[56]}
   );
   gpc1_1 gpc1850 (
      {stage2_10[79]},
      {stage3_10[57]}
   );
   gpc1_1 gpc1851 (
      {stage2_10[80]},
      {stage3_10[58]}
   );
   gpc1_1 gpc1852 (
      {stage2_10[81]},
      {stage3_10[59]}
   );
   gpc1_1 gpc1853 (
      {stage2_10[82]},
      {stage3_10[60]}
   );
   gpc1_1 gpc1854 (
      {stage2_10[83]},
      {stage3_10[61]}
   );
   gpc1_1 gpc1855 (
      {stage2_10[84]},
      {stage3_10[62]}
   );
   gpc1_1 gpc1856 (
      {stage2_10[85]},
      {stage3_10[63]}
   );
   gpc1_1 gpc1857 (
      {stage2_11[129]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1858 (
      {stage2_11[130]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1859 (
      {stage2_11[131]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1860 (
      {stage2_11[132]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1861 (
      {stage2_11[133]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1862 (
      {stage2_11[134]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1863 (
      {stage2_11[135]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1864 (
      {stage2_11[136]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1865 (
      {stage2_11[137]},
      {stage3_11[54]}
   );
   gpc1_1 gpc1866 (
      {stage2_11[138]},
      {stage3_11[55]}
   );
   gpc1_1 gpc1867 (
      {stage2_11[139]},
      {stage3_11[56]}
   );
   gpc1_1 gpc1868 (
      {stage2_11[140]},
      {stage3_11[57]}
   );
   gpc1_1 gpc1869 (
      {stage2_11[141]},
      {stage3_11[58]}
   );
   gpc1_1 gpc1870 (
      {stage2_11[142]},
      {stage3_11[59]}
   );
   gpc1_1 gpc1871 (
      {stage2_11[143]},
      {stage3_11[60]}
   );
   gpc1_1 gpc1872 (
      {stage2_12[72]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1873 (
      {stage2_12[73]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1874 (
      {stage2_12[74]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1875 (
      {stage2_12[75]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1876 (
      {stage2_12[76]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1877 (
      {stage2_12[77]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1878 (
      {stage2_12[78]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1879 (
      {stage2_12[79]},
      {stage3_12[47]}
   );
   gpc1_1 gpc1880 (
      {stage2_12[80]},
      {stage3_12[48]}
   );
   gpc1_1 gpc1881 (
      {stage2_12[81]},
      {stage3_12[49]}
   );
   gpc1_1 gpc1882 (
      {stage2_12[82]},
      {stage3_12[50]}
   );
   gpc1_1 gpc1883 (
      {stage2_12[83]},
      {stage3_12[51]}
   );
   gpc1_1 gpc1884 (
      {stage2_12[84]},
      {stage3_12[52]}
   );
   gpc1_1 gpc1885 (
      {stage2_13[138]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1886 (
      {stage2_13[139]},
      {stage3_13[40]}
   );
   gpc1_1 gpc1887 (
      {stage2_13[140]},
      {stage3_13[41]}
   );
   gpc1_1 gpc1888 (
      {stage2_14[112]},
      {stage3_14[45]}
   );
   gpc1_1 gpc1889 (
      {stage2_14[113]},
      {stage3_14[46]}
   );
   gpc1_1 gpc1890 (
      {stage2_14[114]},
      {stage3_14[47]}
   );
   gpc1_1 gpc1891 (
      {stage2_14[115]},
      {stage3_14[48]}
   );
   gpc1_1 gpc1892 (
      {stage2_14[116]},
      {stage3_14[49]}
   );
   gpc1_1 gpc1893 (
      {stage2_14[117]},
      {stage3_14[50]}
   );
   gpc1_1 gpc1894 (
      {stage2_14[118]},
      {stage3_14[51]}
   );
   gpc1_1 gpc1895 (
      {stage2_14[119]},
      {stage3_14[52]}
   );
   gpc1_1 gpc1896 (
      {stage2_14[120]},
      {stage3_14[53]}
   );
   gpc1_1 gpc1897 (
      {stage2_14[121]},
      {stage3_14[54]}
   );
   gpc1_1 gpc1898 (
      {stage2_14[122]},
      {stage3_14[55]}
   );
   gpc1_1 gpc1899 (
      {stage2_14[123]},
      {stage3_14[56]}
   );
   gpc1_1 gpc1900 (
      {stage2_14[124]},
      {stage3_14[57]}
   );
   gpc1_1 gpc1901 (
      {stage2_15[78]},
      {stage3_15[50]}
   );
   gpc1_1 gpc1902 (
      {stage2_15[79]},
      {stage3_15[51]}
   );
   gpc1_1 gpc1903 (
      {stage2_15[80]},
      {stage3_15[52]}
   );
   gpc1_1 gpc1904 (
      {stage2_15[81]},
      {stage3_15[53]}
   );
   gpc1_1 gpc1905 (
      {stage2_15[82]},
      {stage3_15[54]}
   );
   gpc1_1 gpc1906 (
      {stage2_15[83]},
      {stage3_15[55]}
   );
   gpc1_1 gpc1907 (
      {stage2_15[84]},
      {stage3_15[56]}
   );
   gpc1_1 gpc1908 (
      {stage2_16[92]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1909 (
      {stage2_16[93]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1910 (
      {stage2_16[94]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1911 (
      {stage2_16[95]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1912 (
      {stage2_16[96]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1913 (
      {stage2_16[97]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1914 (
      {stage2_16[98]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1915 (
      {stage2_16[99]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1916 (
      {stage2_16[100]},
      {stage3_16[45]}
   );
   gpc1_1 gpc1917 (
      {stage2_16[101]},
      {stage3_16[46]}
   );
   gpc1_1 gpc1918 (
      {stage2_16[102]},
      {stage3_16[47]}
   );
   gpc1_1 gpc1919 (
      {stage2_16[103]},
      {stage3_16[48]}
   );
   gpc1_1 gpc1920 (
      {stage2_16[104]},
      {stage3_16[49]}
   );
   gpc1_1 gpc1921 (
      {stage2_17[60]},
      {stage3_17[30]}
   );
   gpc1_1 gpc1922 (
      {stage2_17[61]},
      {stage3_17[31]}
   );
   gpc1_1 gpc1923 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1924 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc606_5 gpc1925 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc1926 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1927 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[12]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc615_5 gpc1928 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[13]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc615_5 gpc1929 (
      {stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17], stage3_3[18]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc1930 (
      {stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5]}
   );
   gpc606_5 gpc1931 (
      {stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[4],stage4_5[6],stage4_4[6]}
   );
   gpc615_5 gpc1932 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16]},
      {stage3_6[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[5],stage4_5[7]}
   );
   gpc615_5 gpc1933 (
      {stage3_5[17], stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21]},
      {stage3_6[7]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[6],stage4_5[8]}
   );
   gpc615_5 gpc1934 (
      {stage3_5[22], stage3_5[23], stage3_5[24], stage3_5[25], stage3_5[26]},
      {stage3_6[8]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[7],stage4_5[9]}
   );
   gpc615_5 gpc1935 (
      {stage3_5[27], stage3_5[28], stage3_5[29], stage3_5[30], stage3_5[31]},
      {stage3_6[9]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc1936 (
      {stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35], stage3_5[36]},
      {stage3_6[10]},
      {stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage4_9[4],stage4_8[5],stage4_7[7],stage4_6[9],stage4_5[11]}
   );
   gpc615_5 gpc1937 (
      {stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[11]},
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35]},
      {stage4_9[5],stage4_8[6],stage4_7[8],stage4_6[10],stage4_5[12]}
   );
   gpc615_5 gpc1938 (
      {stage3_5[42], stage3_5[43], stage3_5[44], stage3_5[45], stage3_5[46]},
      {stage3_6[12]},
      {stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41]},
      {stage4_9[6],stage4_8[7],stage4_7[9],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc1939 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[7],stage4_8[8],stage4_7[10],stage4_6[12]}
   );
   gpc606_5 gpc1940 (
      {stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[8],stage4_8[9],stage4_7[11],stage4_6[13]}
   );
   gpc606_5 gpc1941 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29], stage3_6[30]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[9],stage4_8[10],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1942 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[10],stage4_8[11]}
   );
   gpc615_5 gpc1943 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[11],stage4_8[12]}
   );
   gpc606_5 gpc1944 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[12]}
   );
   gpc615_5 gpc1945 (
      {stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12]},
      {stage3_10[12]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[13]}
   );
   gpc615_5 gpc1946 (
      {stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_10[13]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[4],stage4_10[7],stage4_9[14]}
   );
   gpc615_5 gpc1947 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22]},
      {stage3_10[14]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[5],stage4_11[5],stage4_10[8],stage4_9[15]}
   );
   gpc615_5 gpc1948 (
      {stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[6],stage4_11[6],stage4_10[9],stage4_9[16]}
   );
   gpc615_5 gpc1949 (
      {stage3_9[28], stage3_9[29], stage3_9[30], stage3_9[31], stage3_9[32]},
      {stage3_10[16]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[7],stage4_11[7],stage4_10[10],stage4_9[17]}
   );
   gpc615_5 gpc1950 (
      {stage3_9[33], stage3_9[34], stage3_9[35], stage3_9[36], stage3_9[37]},
      {stage3_10[17]},
      {stage3_11[36], stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage4_13[6],stage4_12[8],stage4_11[8],stage4_10[11],stage4_9[18]}
   );
   gpc615_5 gpc1951 (
      {stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41], stage3_9[42]},
      {stage3_10[18]},
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage4_13[7],stage4_12[9],stage4_11[9],stage4_10[12],stage4_9[19]}
   );
   gpc615_5 gpc1952 (
      {stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_10[19]},
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52], stage3_11[53]},
      {stage4_13[8],stage4_12[10],stage4_11[10],stage4_10[13],stage4_9[20]}
   );
   gpc606_5 gpc1953 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[9],stage4_12[11],stage4_11[11],stage4_10[14]}
   );
   gpc606_5 gpc1954 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[10],stage4_12[12],stage4_11[12],stage4_10[15]}
   );
   gpc606_5 gpc1955 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[11],stage4_12[13],stage4_11[13],stage4_10[16]}
   );
   gpc606_5 gpc1956 (
      {stage3_10[38], stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[12],stage4_12[14],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1957 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[4],stage4_13[13],stage4_12[15]}
   );
   gpc606_5 gpc1958 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[5],stage4_13[14],stage4_12[16]}
   );
   gpc606_5 gpc1959 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[2],stage4_14[6],stage4_13[15],stage4_12[17]}
   );
   gpc606_5 gpc1960 (
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[3],stage4_14[7],stage4_13[16],stage4_12[18]}
   );
   gpc1163_5 gpc1961 (
      {stage3_13[0], stage3_13[1], stage3_13[2]},
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[0]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[4],stage4_15[4],stage4_14[8],stage4_13[17]}
   );
   gpc1163_5 gpc1962 (
      {stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[30], stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[1]},
      {stage3_16[1]},
      {stage4_17[1],stage4_16[5],stage4_15[5],stage4_14[9],stage4_13[18]}
   );
   gpc1163_5 gpc1963 (
      {stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[36], stage3_14[37], stage3_14[38], stage3_14[39], stage3_14[40], stage3_14[41]},
      {stage3_15[2]},
      {stage3_16[2]},
      {stage4_17[2],stage4_16[6],stage4_15[6],stage4_14[10],stage4_13[19]}
   );
   gpc1163_5 gpc1964 (
      {stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_14[42], stage3_14[43], stage3_14[44], stage3_14[45], stage3_14[46], stage3_14[47]},
      {stage3_15[3]},
      {stage3_16[3]},
      {stage4_17[3],stage4_16[7],stage4_15[7],stage4_14[11],stage4_13[20]}
   );
   gpc606_5 gpc1965 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[4],stage4_16[8],stage4_15[8],stage4_14[12],stage4_13[21]}
   );
   gpc606_5 gpc1966 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[5],stage4_16[9],stage4_15[9],stage4_14[13],stage4_13[22]}
   );
   gpc606_5 gpc1967 (
      {stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29]},
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage4_17[6],stage4_16[10],stage4_15[10],stage4_14[14],stage4_13[23]}
   );
   gpc606_5 gpc1968 (
      {stage3_13[30], stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35]},
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27]},
      {stage4_17[7],stage4_16[11],stage4_15[11],stage4_14[15],stage4_13[24]}
   );
   gpc606_5 gpc1969 (
      {stage3_13[36], stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41]},
      {stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33]},
      {stage4_17[8],stage4_16[12],stage4_15[12],stage4_14[16],stage4_13[25]}
   );
   gpc615_5 gpc1970 (
      {stage3_14[48], stage3_14[49], stage3_14[50], stage3_14[51], stage3_14[52]},
      {stage3_15[34]},
      {stage3_16[4], stage3_16[5], stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9]},
      {stage4_18[0],stage4_17[9],stage4_16[13],stage4_15[13],stage4_14[17]}
   );
   gpc615_5 gpc1971 (
      {stage3_14[53], stage3_14[54], stage3_14[55], stage3_14[56], stage3_14[57]},
      {stage3_15[35]},
      {stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage4_18[1],stage4_17[10],stage4_16[14],stage4_15[14],stage4_14[18]}
   );
   gpc606_5 gpc1972 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40], stage3_15[41]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[2],stage4_17[11],stage4_16[15],stage4_15[15]}
   );
   gpc606_5 gpc1973 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46], stage3_15[47]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[3],stage4_17[12],stage4_16[16],stage4_15[16]}
   );
   gpc615_5 gpc1974 (
      {stage3_15[48], stage3_15[49], stage3_15[50], stage3_15[51], stage3_15[52]},
      {stage3_16[16]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[4],stage4_17[13],stage4_16[17],stage4_15[17]}
   );
   gpc606_5 gpc1975 (
      {stage3_16[17], stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[5],stage4_17[14],stage4_16[18]}
   );
   gpc606_5 gpc1976 (
      {stage3_16[23], stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[6],stage4_17[15],stage4_16[19]}
   );
   gpc606_5 gpc1977 (
      {stage3_16[29], stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34]},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[5],stage4_18[7],stage4_17[16],stage4_16[20]}
   );
   gpc606_5 gpc1978 (
      {stage3_16[35], stage3_16[36], stage3_16[37], stage3_16[38], stage3_16[39], stage3_16[40]},
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23]},
      {stage4_20[3],stage4_19[6],stage4_18[8],stage4_17[17],stage4_16[21]}
   );
   gpc606_5 gpc1979 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[7],stage4_18[9],stage4_17[18]}
   );
   gpc606_5 gpc1980 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[8],stage4_18[10],stage4_17[19]}
   );
   gpc1_1 gpc1981 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1982 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1983 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1984 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1985 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1986 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1987 (
      {stage3_2[10]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1988 (
      {stage3_2[11]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1989 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1990 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1991 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1992 (
      {stage3_2[15]},
      {stage4_2[9]}
   );
   gpc1_1 gpc1993 (
      {stage3_2[16]},
      {stage4_2[10]}
   );
   gpc1_1 gpc1994 (
      {stage3_3[24]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1995 (
      {stage3_3[25]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1996 (
      {stage3_3[26]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1997 (
      {stage3_3[27]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1998 (
      {stage3_3[28]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1999 (
      {stage3_4[20]},
      {stage4_4[7]}
   );
   gpc1_1 gpc2000 (
      {stage3_4[21]},
      {stage4_4[8]}
   );
   gpc1_1 gpc2001 (
      {stage3_4[22]},
      {stage4_4[9]}
   );
   gpc1_1 gpc2002 (
      {stage3_4[23]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2003 (
      {stage3_4[24]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2004 (
      {stage3_4[25]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2005 (
      {stage3_4[26]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2006 (
      {stage3_4[27]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2007 (
      {stage3_4[28]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2008 (
      {stage3_4[29]},
      {stage4_4[16]}
   );
   gpc1_1 gpc2009 (
      {stage3_4[30]},
      {stage4_4[17]}
   );
   gpc1_1 gpc2010 (
      {stage3_4[31]},
      {stage4_4[18]}
   );
   gpc1_1 gpc2011 (
      {stage3_4[32]},
      {stage4_4[19]}
   );
   gpc1_1 gpc2012 (
      {stage3_4[33]},
      {stage4_4[20]}
   );
   gpc1_1 gpc2013 (
      {stage3_4[34]},
      {stage4_4[21]}
   );
   gpc1_1 gpc2014 (
      {stage3_4[35]},
      {stage4_4[22]}
   );
   gpc1_1 gpc2015 (
      {stage3_4[36]},
      {stage4_4[23]}
   );
   gpc1_1 gpc2016 (
      {stage3_4[37]},
      {stage4_4[24]}
   );
   gpc1_1 gpc2017 (
      {stage3_4[38]},
      {stage4_4[25]}
   );
   gpc1_1 gpc2018 (
      {stage3_4[39]},
      {stage4_4[26]}
   );
   gpc1_1 gpc2019 (
      {stage3_5[47]},
      {stage4_5[14]}
   );
   gpc1_1 gpc2020 (
      {stage3_6[31]},
      {stage4_6[15]}
   );
   gpc1_1 gpc2021 (
      {stage3_6[32]},
      {stage4_6[16]}
   );
   gpc1_1 gpc2022 (
      {stage3_6[33]},
      {stage4_6[17]}
   );
   gpc1_1 gpc2023 (
      {stage3_6[34]},
      {stage4_6[18]}
   );
   gpc1_1 gpc2024 (
      {stage3_6[35]},
      {stage4_6[19]}
   );
   gpc1_1 gpc2025 (
      {stage3_6[36]},
      {stage4_6[20]}
   );
   gpc1_1 gpc2026 (
      {stage3_6[37]},
      {stage4_6[21]}
   );
   gpc1_1 gpc2027 (
      {stage3_7[42]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2028 (
      {stage3_7[43]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2029 (
      {stage3_7[44]},
      {stage4_7[15]}
   );
   gpc1_1 gpc2030 (
      {stage3_7[45]},
      {stage4_7[16]}
   );
   gpc1_1 gpc2031 (
      {stage3_8[28]},
      {stage4_8[13]}
   );
   gpc1_1 gpc2032 (
      {stage3_8[29]},
      {stage4_8[14]}
   );
   gpc1_1 gpc2033 (
      {stage3_8[30]},
      {stage4_8[15]}
   );
   gpc1_1 gpc2034 (
      {stage3_8[31]},
      {stage4_8[16]}
   );
   gpc1_1 gpc2035 (
      {stage3_8[32]},
      {stage4_8[17]}
   );
   gpc1_1 gpc2036 (
      {stage3_8[33]},
      {stage4_8[18]}
   );
   gpc1_1 gpc2037 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc2038 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc2039 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc2040 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc2041 (
      {stage3_8[38]},
      {stage4_8[23]}
   );
   gpc1_1 gpc2042 (
      {stage3_8[39]},
      {stage4_8[24]}
   );
   gpc1_1 gpc2043 (
      {stage3_8[40]},
      {stage4_8[25]}
   );
   gpc1_1 gpc2044 (
      {stage3_9[48]},
      {stage4_9[21]}
   );
   gpc1_1 gpc2045 (
      {stage3_9[49]},
      {stage4_9[22]}
   );
   gpc1_1 gpc2046 (
      {stage3_9[50]},
      {stage4_9[23]}
   );
   gpc1_1 gpc2047 (
      {stage3_9[51]},
      {stage4_9[24]}
   );
   gpc1_1 gpc2048 (
      {stage3_10[44]},
      {stage4_10[18]}
   );
   gpc1_1 gpc2049 (
      {stage3_10[45]},
      {stage4_10[19]}
   );
   gpc1_1 gpc2050 (
      {stage3_10[46]},
      {stage4_10[20]}
   );
   gpc1_1 gpc2051 (
      {stage3_10[47]},
      {stage4_10[21]}
   );
   gpc1_1 gpc2052 (
      {stage3_10[48]},
      {stage4_10[22]}
   );
   gpc1_1 gpc2053 (
      {stage3_10[49]},
      {stage4_10[23]}
   );
   gpc1_1 gpc2054 (
      {stage3_10[50]},
      {stage4_10[24]}
   );
   gpc1_1 gpc2055 (
      {stage3_10[51]},
      {stage4_10[25]}
   );
   gpc1_1 gpc2056 (
      {stage3_10[52]},
      {stage4_10[26]}
   );
   gpc1_1 gpc2057 (
      {stage3_10[53]},
      {stage4_10[27]}
   );
   gpc1_1 gpc2058 (
      {stage3_10[54]},
      {stage4_10[28]}
   );
   gpc1_1 gpc2059 (
      {stage3_10[55]},
      {stage4_10[29]}
   );
   gpc1_1 gpc2060 (
      {stage3_10[56]},
      {stage4_10[30]}
   );
   gpc1_1 gpc2061 (
      {stage3_10[57]},
      {stage4_10[31]}
   );
   gpc1_1 gpc2062 (
      {stage3_10[58]},
      {stage4_10[32]}
   );
   gpc1_1 gpc2063 (
      {stage3_10[59]},
      {stage4_10[33]}
   );
   gpc1_1 gpc2064 (
      {stage3_10[60]},
      {stage4_10[34]}
   );
   gpc1_1 gpc2065 (
      {stage3_10[61]},
      {stage4_10[35]}
   );
   gpc1_1 gpc2066 (
      {stage3_10[62]},
      {stage4_10[36]}
   );
   gpc1_1 gpc2067 (
      {stage3_10[63]},
      {stage4_10[37]}
   );
   gpc1_1 gpc2068 (
      {stage3_11[54]},
      {stage4_11[15]}
   );
   gpc1_1 gpc2069 (
      {stage3_11[55]},
      {stage4_11[16]}
   );
   gpc1_1 gpc2070 (
      {stage3_11[56]},
      {stage4_11[17]}
   );
   gpc1_1 gpc2071 (
      {stage3_11[57]},
      {stage4_11[18]}
   );
   gpc1_1 gpc2072 (
      {stage3_11[58]},
      {stage4_11[19]}
   );
   gpc1_1 gpc2073 (
      {stage3_11[59]},
      {stage4_11[20]}
   );
   gpc1_1 gpc2074 (
      {stage3_11[60]},
      {stage4_11[21]}
   );
   gpc1_1 gpc2075 (
      {stage3_12[48]},
      {stage4_12[19]}
   );
   gpc1_1 gpc2076 (
      {stage3_12[49]},
      {stage4_12[20]}
   );
   gpc1_1 gpc2077 (
      {stage3_12[50]},
      {stage4_12[21]}
   );
   gpc1_1 gpc2078 (
      {stage3_12[51]},
      {stage4_12[22]}
   );
   gpc1_1 gpc2079 (
      {stage3_12[52]},
      {stage4_12[23]}
   );
   gpc1_1 gpc2080 (
      {stage3_15[53]},
      {stage4_15[18]}
   );
   gpc1_1 gpc2081 (
      {stage3_15[54]},
      {stage4_15[19]}
   );
   gpc1_1 gpc2082 (
      {stage3_15[55]},
      {stage4_15[20]}
   );
   gpc1_1 gpc2083 (
      {stage3_15[56]},
      {stage4_15[21]}
   );
   gpc1_1 gpc2084 (
      {stage3_16[41]},
      {stage4_16[22]}
   );
   gpc1_1 gpc2085 (
      {stage3_16[42]},
      {stage4_16[23]}
   );
   gpc1_1 gpc2086 (
      {stage3_16[43]},
      {stage4_16[24]}
   );
   gpc1_1 gpc2087 (
      {stage3_16[44]},
      {stage4_16[25]}
   );
   gpc1_1 gpc2088 (
      {stage3_16[45]},
      {stage4_16[26]}
   );
   gpc1_1 gpc2089 (
      {stage3_16[46]},
      {stage4_16[27]}
   );
   gpc1_1 gpc2090 (
      {stage3_16[47]},
      {stage4_16[28]}
   );
   gpc1_1 gpc2091 (
      {stage3_16[48]},
      {stage4_16[29]}
   );
   gpc1_1 gpc2092 (
      {stage3_16[49]},
      {stage4_16[30]}
   );
   gpc1_1 gpc2093 (
      {stage3_17[30]},
      {stage4_17[20]}
   );
   gpc1_1 gpc2094 (
      {stage3_17[31]},
      {stage4_17[21]}
   );
   gpc1_1 gpc2095 (
      {stage3_18[24]},
      {stage4_18[11]}
   );
   gpc1_1 gpc2096 (
      {stage3_18[25]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2097 (
      {stage3_19[12]},
      {stage4_19[9]}
   );
   gpc1_1 gpc2098 (
      {stage3_19[13]},
      {stage4_19[10]}
   );
   gpc1_1 gpc2099 (
      {stage3_20[0]},
      {stage4_20[6]}
   );
   gpc1_1 gpc2100 (
      {stage3_20[1]},
      {stage4_20[7]}
   );
   gpc1_1 gpc2101 (
      {stage3_20[2]},
      {stage4_20[8]}
   );
   gpc1_1 gpc2102 (
      {stage3_20[3]},
      {stage4_20[9]}
   );
   gpc1_1 gpc2103 (
      {stage3_20[4]},
      {stage4_20[10]}
   );
   gpc1_1 gpc2104 (
      {stage3_20[5]},
      {stage4_20[11]}
   );
   gpc1_1 gpc2105 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc1_1 gpc2106 (
      {stage3_21[1]},
      {stage4_21[3]}
   );
   gpc615_5 gpc2107 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc606_5 gpc2108 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1406_5 gpc2109 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc606_5 gpc2110 (
      {stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16], stage4_4[17]},
      {stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9]},
      {stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc606_5 gpc2111 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc615_5 gpc2112 (
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[3],stage5_7[4]}
   );
   gpc615_5 gpc2113 (
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[2],stage5_8[4],stage5_7[5]}
   );
   gpc1163_5 gpc2114 (
      {stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17]},
      {stage4_10[0]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[3],stage5_8[5]}
   );
   gpc1163_5 gpc2115 (
      {stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_9[18], stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23]},
      {stage4_10[1]},
      {stage4_11[1]},
      {stage5_12[1],stage5_11[3],stage5_10[3],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc2116 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12], stage4_8[13]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[2],stage5_11[4],stage5_10[4],stage5_9[5],stage5_8[7]}
   );
   gpc606_5 gpc2117 (
      {stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17], stage4_8[18], stage4_8[19]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[3],stage5_11[5],stage5_10[5],stage5_9[6],stage5_8[8]}
   );
   gpc606_5 gpc2118 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19]},
      {stage5_12[4],stage5_11[6],stage5_10[6],stage5_9[7],stage5_8[9]}
   );
   gpc606_5 gpc2119 (
      {stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24], stage4_10[25]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[5],stage5_11[7],stage5_10[7]}
   );
   gpc606_5 gpc2120 (
      {stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30], stage4_10[31]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[1],stage5_12[6],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc2121 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[12]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc2122 (
      {stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage4_12[13]},
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[8],stage5_11[10]}
   );
   gpc615_5 gpc2123 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16]},
      {stage4_12[14]},
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[9],stage5_11[11]}
   );
   gpc615_5 gpc2124 (
      {stage4_11[17], stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21]},
      {stage4_12[15]},
      {stage4_13[18], stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[10],stage5_11[12]}
   );
   gpc606_5 gpc2125 (
      {stage4_12[16], stage4_12[17], stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[11]}
   );
   gpc615_5 gpc2126 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc2127 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc2128 (
      {stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage4_16[12]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7]}
   );
   gpc615_5 gpc2129 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[13]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8]}
   );
   gpc615_5 gpc2130 (
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16]},
      {stage4_16[14]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc606_5 gpc2131 (
      {stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18], stage4_16[19], stage4_16[20]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[3],stage5_18[5],stage5_17[5],stage5_16[6]}
   );
   gpc606_5 gpc2132 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], 1'b0, 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[4],stage5_18[6],stage5_17[6]}
   );
   gpc606_5 gpc2133 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[5],stage5_18[7]}
   );
   gpc1343_5 gpc2134 (
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {1'b0},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[6]}
   );
   gpc1_1 gpc2135 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc2136 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc2137 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc2138 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc2139 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc2140 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc2141 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2142 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2143 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2144 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2145 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2146 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2147 (
      {stage4_2[9]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2148 (
      {stage4_2[10]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2149 (
      {stage4_3[7]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2150 (
      {stage4_3[8]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2151 (
      {stage4_3[9]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2152 (
      {stage4_3[10]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2153 (
      {stage4_4[18]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2154 (
      {stage4_4[19]},
      {stage5_4[5]}
   );
   gpc1_1 gpc2155 (
      {stage4_4[20]},
      {stage5_4[6]}
   );
   gpc1_1 gpc2156 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc2157 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc2158 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc2159 (
      {stage4_4[24]},
      {stage5_4[10]}
   );
   gpc1_1 gpc2160 (
      {stage4_4[25]},
      {stage5_4[11]}
   );
   gpc1_1 gpc2161 (
      {stage4_4[26]},
      {stage5_4[12]}
   );
   gpc1_1 gpc2162 (
      {stage4_5[12]},
      {stage5_5[5]}
   );
   gpc1_1 gpc2163 (
      {stage4_5[13]},
      {stage5_5[6]}
   );
   gpc1_1 gpc2164 (
      {stage4_5[14]},
      {stage5_5[7]}
   );
   gpc1_1 gpc2165 (
      {stage4_6[10]},
      {stage5_6[5]}
   );
   gpc1_1 gpc2166 (
      {stage4_6[11]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2167 (
      {stage4_6[12]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2168 (
      {stage4_6[13]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2169 (
      {stage4_6[14]},
      {stage5_6[9]}
   );
   gpc1_1 gpc2170 (
      {stage4_6[15]},
      {stage5_6[10]}
   );
   gpc1_1 gpc2171 (
      {stage4_6[16]},
      {stage5_6[11]}
   );
   gpc1_1 gpc2172 (
      {stage4_6[17]},
      {stage5_6[12]}
   );
   gpc1_1 gpc2173 (
      {stage4_6[18]},
      {stage5_6[13]}
   );
   gpc1_1 gpc2174 (
      {stage4_6[19]},
      {stage5_6[14]}
   );
   gpc1_1 gpc2175 (
      {stage4_6[20]},
      {stage5_6[15]}
   );
   gpc1_1 gpc2176 (
      {stage4_6[21]},
      {stage5_6[16]}
   );
   gpc1_1 gpc2177 (
      {stage4_9[24]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2178 (
      {stage4_10[32]},
      {stage5_10[9]}
   );
   gpc1_1 gpc2179 (
      {stage4_10[33]},
      {stage5_10[10]}
   );
   gpc1_1 gpc2180 (
      {stage4_10[34]},
      {stage5_10[11]}
   );
   gpc1_1 gpc2181 (
      {stage4_10[35]},
      {stage5_10[12]}
   );
   gpc1_1 gpc2182 (
      {stage4_10[36]},
      {stage5_10[13]}
   );
   gpc1_1 gpc2183 (
      {stage4_10[37]},
      {stage5_10[14]}
   );
   gpc1_1 gpc2184 (
      {stage4_12[22]},
      {stage5_12[12]}
   );
   gpc1_1 gpc2185 (
      {stage4_12[23]},
      {stage5_12[13]}
   );
   gpc1_1 gpc2186 (
      {stage4_13[24]},
      {stage5_13[7]}
   );
   gpc1_1 gpc2187 (
      {stage4_13[25]},
      {stage5_13[8]}
   );
   gpc1_1 gpc2188 (
      {stage4_14[16]},
      {stage5_14[9]}
   );
   gpc1_1 gpc2189 (
      {stage4_14[17]},
      {stage5_14[10]}
   );
   gpc1_1 gpc2190 (
      {stage4_14[18]},
      {stage5_14[11]}
   );
   gpc1_1 gpc2191 (
      {stage4_15[17]},
      {stage5_15[10]}
   );
   gpc1_1 gpc2192 (
      {stage4_15[18]},
      {stage5_15[11]}
   );
   gpc1_1 gpc2193 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc2194 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc2195 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc2196 (
      {stage4_16[21]},
      {stage5_16[7]}
   );
   gpc1_1 gpc2197 (
      {stage4_16[22]},
      {stage5_16[8]}
   );
   gpc1_1 gpc2198 (
      {stage4_16[23]},
      {stage5_16[9]}
   );
   gpc1_1 gpc2199 (
      {stage4_16[24]},
      {stage5_16[10]}
   );
   gpc1_1 gpc2200 (
      {stage4_16[25]},
      {stage5_16[11]}
   );
   gpc1_1 gpc2201 (
      {stage4_16[26]},
      {stage5_16[12]}
   );
   gpc1_1 gpc2202 (
      {stage4_16[27]},
      {stage5_16[13]}
   );
   gpc1_1 gpc2203 (
      {stage4_16[28]},
      {stage5_16[14]}
   );
   gpc1_1 gpc2204 (
      {stage4_16[29]},
      {stage5_16[15]}
   );
   gpc1_1 gpc2205 (
      {stage4_16[30]},
      {stage5_16[16]}
   );
   gpc1_1 gpc2206 (
      {stage4_18[12]},
      {stage5_18[8]}
   );
   gpc1_1 gpc2207 (
      {stage4_19[9]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2208 (
      {stage4_19[10]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2209 (
      {stage4_20[10]},
      {stage5_20[4]}
   );
   gpc1_1 gpc2210 (
      {stage4_20[11]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2211 (
      {stage4_21[3]},
      {stage5_21[3]}
   );
   gpc1163_5 gpc2212 (
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[0]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc207_4 gpc2213 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[0],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc7_3 gpc2214 (
      {stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5], stage5_5[6], stage5_5[7]},
      {stage6_7[1],stage6_6[2],stage6_5[2]}
   );
   gpc1325_5 gpc2215 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[3]}
   );
   gpc1325_5 gpc2216 (
      {stage5_6[7], stage5_6[8], stage5_6[9], stage5_6[10], stage5_6[11]},
      {stage5_7[2], stage5_7[3]},
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[4]}
   );
   gpc1325_5 gpc2217 (
      {stage5_6[12], stage5_6[13], stage5_6[14], stage5_6[15], stage5_6[16]},
      {stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7], stage5_8[8]},
      {stage5_9[2]},
      {stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[5]}
   );
   gpc1163_5 gpc2218 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[3]}
   );
   gpc1163_5 gpc2219 (
      {stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage5_11[6], stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11]},
      {stage5_12[1]},
      {stage5_13[1]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[1],stage6_10[4]}
   );
   gpc615_5 gpc2220 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10]},
      {stage5_11[12]},
      {stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7]},
      {stage6_14[2],stage6_13[2],stage6_12[2],stage6_11[2],stage6_10[5]}
   );
   gpc2116_5 gpc2221 (
      {stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {stage5_13[2]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[3]}
   );
   gpc623_5 gpc2222 (
      {stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[1], stage5_14[2]},
      {stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc1423_5 gpc2223 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5]}
   );
   gpc615_5 gpc2224 (
      {stage5_14[6], stage5_14[7], stage5_14[8], stage5_14[9], stage5_14[10]},
      {stage5_15[10]},
      {stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], stage5_16[8], stage5_16[9]},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[3],stage6_14[6]}
   );
   gpc606_5 gpc2225 (
      {stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14], stage5_16[15]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[3],stage6_16[4]}
   );
   gpc606_5 gpc2226 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[1],stage6_19[1],stage6_18[3],stage6_17[4]}
   );
   gpc1_1 gpc2227 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc2228 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2229 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2230 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2231 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2232 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2233 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc2234 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2235 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc2236 (
      {stage5_2[4]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2237 (
      {stage5_2[5]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2238 (
      {stage5_2[6]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2239 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2240 (
      {stage5_4[9]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2241 (
      {stage5_4[10]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2242 (
      {stage5_4[11]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2243 (
      {stage5_4[12]},
      {stage6_4[6]}
   );
   gpc1_1 gpc2244 (
      {stage5_8[9]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2245 (
      {stage5_9[3]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2246 (
      {stage5_9[4]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2247 (
      {stage5_9[5]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2248 (
      {stage5_9[6]},
      {stage6_9[6]}
   );
   gpc1_1 gpc2249 (
      {stage5_9[7]},
      {stage6_9[7]}
   );
   gpc1_1 gpc2250 (
      {stage5_9[8]},
      {stage6_9[8]}
   );
   gpc1_1 gpc2251 (
      {stage5_10[11]},
      {stage6_10[6]}
   );
   gpc1_1 gpc2252 (
      {stage5_10[12]},
      {stage6_10[7]}
   );
   gpc1_1 gpc2253 (
      {stage5_10[13]},
      {stage6_10[8]}
   );
   gpc1_1 gpc2254 (
      {stage5_10[14]},
      {stage6_10[9]}
   );
   gpc1_1 gpc2255 (
      {stage5_13[6]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2256 (
      {stage5_13[7]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2257 (
      {stage5_13[8]},
      {stage6_13[7]}
   );
   gpc1_1 gpc2258 (
      {stage5_14[11]},
      {stage6_14[7]}
   );
   gpc1_1 gpc2259 (
      {stage5_15[11]},
      {stage6_15[4]}
   );
   gpc1_1 gpc2260 (
      {stage5_15[12]},
      {stage6_15[5]}
   );
   gpc1_1 gpc2261 (
      {stage5_15[13]},
      {stage6_15[6]}
   );
   gpc1_1 gpc2262 (
      {stage5_15[14]},
      {stage6_15[7]}
   );
   gpc1_1 gpc2263 (
      {stage5_16[16]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2264 (
      {stage5_18[6]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2265 (
      {stage5_18[7]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2266 (
      {stage5_18[8]},
      {stage6_18[6]}
   );
   gpc1_1 gpc2267 (
      {stage5_19[6]},
      {stage6_19[2]}
   );
   gpc1_1 gpc2268 (
      {stage5_19[7]},
      {stage6_19[3]}
   );
   gpc1_1 gpc2269 (
      {stage5_19[8]},
      {stage6_19[4]}
   );
   gpc1_1 gpc2270 (
      {stage5_20[0]},
      {stage6_20[2]}
   );
   gpc1_1 gpc2271 (
      {stage5_20[1]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2272 (
      {stage5_20[2]},
      {stage6_20[4]}
   );
   gpc1_1 gpc2273 (
      {stage5_20[3]},
      {stage6_20[5]}
   );
   gpc1_1 gpc2274 (
      {stage5_20[4]},
      {stage6_20[6]}
   );
   gpc1_1 gpc2275 (
      {stage5_20[5]},
      {stage6_20[7]}
   );
   gpc1_1 gpc2276 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc2277 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc2278 (
      {stage5_21[2]},
      {stage6_21[3]}
   );
   gpc1_1 gpc2279 (
      {stage5_21[3]},
      {stage6_21[4]}
   );
   gpc1_1 gpc2280 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
   gpc1_1 gpc2281 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc2282 (
      {stage5_23[0]},
      {stage6_23[0]}
   );
   gpc1406_5 gpc2283 (
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[0]}
   );
   gpc117_4 gpc2284 (
      {stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5], stage6_9[6], stage6_9[7]},
      {stage6_10[0]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc1415_5 gpc2285 (
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[2]}
   );
   gpc606_5 gpc2286 (
      {stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc606_5 gpc2287 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[1],stage7_16[1],stage7_15[1],stage7_14[2]}
   );
   gpc606_5 gpc2288 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc1406_5 gpc2289 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc1_1 gpc2290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc2291 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2292 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc2293 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc2294 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc2295 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc2296 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc2297 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2298 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc2299 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc2300 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc2301 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc2302 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc2303 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc2304 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc2305 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc2306 (
      {stage6_4[2]},
      {stage7_4[2]}
   );
   gpc1_1 gpc2307 (
      {stage6_4[3]},
      {stage7_4[3]}
   );
   gpc1_1 gpc2308 (
      {stage6_4[4]},
      {stage7_4[4]}
   );
   gpc1_1 gpc2309 (
      {stage6_4[5]},
      {stage7_4[5]}
   );
   gpc1_1 gpc2310 (
      {stage6_4[6]},
      {stage7_4[6]}
   );
   gpc1_1 gpc2311 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc2312 (
      {stage6_5[1]},
      {stage7_5[1]}
   );
   gpc1_1 gpc2313 (
      {stage6_5[2]},
      {stage7_5[2]}
   );
   gpc1_1 gpc2314 (
      {stage6_7[0]},
      {stage7_7[1]}
   );
   gpc1_1 gpc2315 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc2316 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc2317 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc2318 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc2319 (
      {stage6_9[8]},
      {stage7_9[2]}
   );
   gpc1_1 gpc2320 (
      {stage6_10[6]},
      {stage7_10[3]}
   );
   gpc1_1 gpc2321 (
      {stage6_10[7]},
      {stage7_10[4]}
   );
   gpc1_1 gpc2322 (
      {stage6_10[8]},
      {stage7_10[5]}
   );
   gpc1_1 gpc2323 (
      {stage6_10[9]},
      {stage7_10[6]}
   );
   gpc1_1 gpc2324 (
      {stage6_11[2]},
      {stage7_11[2]}
   );
   gpc1_1 gpc2325 (
      {stage6_13[7]},
      {stage7_13[2]}
   );
   gpc1_1 gpc2326 (
      {stage6_14[6]},
      {stage7_14[3]}
   );
   gpc1_1 gpc2327 (
      {stage6_14[7]},
      {stage7_14[4]}
   );
   gpc1_1 gpc2328 (
      {stage6_15[6]},
      {stage7_15[2]}
   );
   gpc1_1 gpc2329 (
      {stage6_15[7]},
      {stage7_15[3]}
   );
   gpc1_1 gpc2330 (
      {stage6_17[0]},
      {stage7_17[2]}
   );
   gpc1_1 gpc2331 (
      {stage6_17[1]},
      {stage7_17[3]}
   );
   gpc1_1 gpc2332 (
      {stage6_17[2]},
      {stage7_17[4]}
   );
   gpc1_1 gpc2333 (
      {stage6_17[3]},
      {stage7_17[5]}
   );
   gpc1_1 gpc2334 (
      {stage6_17[4]},
      {stage7_17[6]}
   );
   gpc1_1 gpc2335 (
      {stage6_18[6]},
      {stage7_18[2]}
   );
   gpc1_1 gpc2336 (
      {stage6_20[6]},
      {stage7_20[2]}
   );
   gpc1_1 gpc2337 (
      {stage6_20[7]},
      {stage7_20[3]}
   );
   gpc1_1 gpc2338 (
      {stage6_21[4]},
      {stage7_21[2]}
   );
   gpc1_1 gpc2339 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc2340 (
      {stage6_23[0]},
      {stage7_23[1]}
   );
   gpc615_5 gpc2341 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc7_3 gpc2342 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc615_5 gpc2343 (
      {stage7_5[0], stage7_5[1], stage7_5[2], 1'b0, 1'b0},
      {stage7_6[0]},
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5]},
      {stage8_9[0],stage8_8[0],stage8_7[0],stage8_6[1],stage8_5[1]}
   );
   gpc23_3 gpc2344 (
      {stage7_9[0], stage7_9[1], stage7_9[2]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc135_4 gpc2345 (
      {stage7_10[2], stage7_10[3], stage7_10[4], stage7_10[5], stage7_10[6]},
      {stage7_11[0], stage7_11[1], stage7_11[2]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1]}
   );
   gpc1343_5 gpc2346 (
      {stage7_13[0], stage7_13[1], stage7_13[2]},
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3]},
      {stage7_15[0], stage7_15[1], stage7_15[2]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc7_3 gpc2347 (
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3], stage7_17[4], stage7_17[5], stage7_17[6]},
      {stage8_19[0],stage8_18[0],stage8_17[1]}
   );
   gpc1325_5 gpc2348 (
      {stage7_18[0], stage7_18[1], stage7_18[2], 1'b0, 1'b0},
      {stage7_19[0], stage7_19[1]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1],stage8_18[1]}
   );
   gpc1163_5 gpc2349 (
      {stage7_21[1], stage7_21[2], 1'b0},
      {stage7_22[0], stage7_22[1], stage7_22[2], 1'b0, 1'b0, 1'b0},
      {stage7_23[0]},
      {1'b0},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1]}
   );
   gpc1_1 gpc2350 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc2351 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc2352 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc2353 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc2354 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc2355 (
      {stage7_14[4]},
      {stage8_14[1]}
   );
   gpc1_1 gpc2356 (
      {stage7_15[3]},
      {stage8_15[1]}
   );
   gpc1_1 gpc2357 (
      {stage7_16[1]},
      {stage8_16[1]}
   );
   gpc1_1 gpc2358 (
      {stage7_20[3]},
      {stage8_20[1]}
   );
   gpc1_1 gpc2359 (
      {stage7_23[1]},
      {stage8_23[1]}
   );
endmodule
module rowadder2_1_25(input [24:0] src0, input [24:0] src1, output [25:0] dst0);
    wire [24:0] gene;
    wire [24:0] prop;
    wire [27:0] out;
    wire [27:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[24:24]}),
        .S({3'h0, prop[24:24]})
    );
    assign dst0 = {carryout[24], out[24:0]};
endmodule


module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor2_1_512_16 compressor2_1_512_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9b3efca63c51239e96acb4cc372b3030f8ef75adc0c2cd4f1d9456a0795c079cae4e548cc6fbd8bec4b914689bc86fce47a3978c0d4070c3b33657207bdcf58f2049c6fbb90e2a230a04d9f74031c0ab85293e0dac4b87de8f6787d2c280cb0dac1cf11daadc9a1ccb6f5643996612d8a4cdb14ec76b0ac011824df14b4d15bd5918930cd6555dd590a964aef7b4168b07c72e57852cffc063c629114723e9746516f43395f1e5aa6067e4ff93462a5f64dce94a320ed26cfe0cd62bce081da246b96051da647c2895c8a9042b332b7cf14cae8cecdc47df806388f5a8764785a8a01ee0e7d01047aa87f8d0d62421f7fc0a21173a777d5f417da79a294934df19f2e3b134db0bb343badb7d4e766de02d90a4bc37003522f769891d4802e16854206e2a503cee76b28b6092fe9e8e65f9db16048130faeea28e4da879f9d69347717ec7998377d1ad3742901af6e783f439f0eafe4d9772dadd73bb44e106517c9239a5c9a7de92af20a7929fcfcf6aaa0fd597f3284938d663e0149054948c47e8e439746ed1a9589b982c783a1e419a249134f991c51450ede8548c23bf5b2397525478eb7351a2045db8619f687ceb82f0b24539465c1279fb83a4037915692fb3cfc49ca111c45bd81ad972dca4438f00f1252f7cf324b3ea4bfdcced54465448296df4aa825024140547555c6cd75aac5e2774556c48c723fcfad8ef451ea28305c7a4d99e6dab90d74d9693bb1768c97490f149654f3315d8647f5d2ac38bbbd670f6b9ff43c4921b2f374f98eb75c85a47a27b01ccdece969f48676fed8fdbd92054cb8abb9be4544099dac3bbfafe6e38924aecd1a006163782230b4ad827e8b605fe1828485dda67b27f7f0fa3808d76e5a2620bf48f8aeda9c2b3bc110affeea66969ab65cdef03236547ce84889c9d9e32d18c4abc605c36368bc811d9023fec6ff7de37efc0712b69a849e9a97f0dd58614e8e49c2237e67c3b5211e3b51f84ff15e5bb808a022d486e39914bb4ee69fa545d1c3a6f2813421582a9cccdb3839ac076017cf1c57cb68880ba10d22a9744d9ba88f42ec2c0dba0e0a6b1165e35852d1865037bebb2e392c0300699d6783c9bbe798c62a3e56dabd65694764131252a449bac58f970ecf6fb8cc8dbc3ac196d2cc1f01394230da22ced11a80070999bfd82ad282de5f82c18944a9c6a82b9948000c02c103137805988d1a8eb310a3e961781e78abd65277a8edb0433a53eebba0b4d38ee74da21a899847b29fa5dd68f7366f2a65edd2159d37c6eabb6bc6a2681c32076d19108b8c298da35052a8d752d72f6eacc2bddc10ef36e805c0d558ac35ca3e603d8f816f002ba3627a1380b6d9a9f05c86c1f4d9c58f30c85305497ce9d4272468c53f0cb3185112fb6b357de3b7ad44716fd51b24d08eb09eda12296ba8907a0cf2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe88152dee5c1606a9720890c53406ace8d5eeacf16499e3c3b536922d3375dbd7508c9b2d8eddd354b536e38230dd9068328ec74e2cf4156c5c591570f8e05d18bc19a09e3742fe4b917d1b60322f012229060cce062a5dba25a66d170430c9422eaa2fc6876119039bb0f2b6240e5b4a684e05c5278615370eb96b3d6b4135d5c893f78e0f99b33d29ace7f398d49f3492472f826c64774870c31f131ac869efe3b8e3d2b74f337bb9dcc1993915cf72193f26854097d97f26c87b6186bc452567a95f434917748841ae5d7c949e9f3bddefebb648494484ca661a3fec744da32b879e4c1d6a818ab094d88d48add03d6bc4e3740d84d43e246f89d5eee6ba61f3748b31a74e8611afa1c5f0b85195d3eb5ca6c18dfa49900b507e34ae7c89893db031c0f6ef847442bdff2eae99d0e7aaa8212771fe7006ce22a7d0f0b06843622b503b43052a994ce7c366f846c5886d05ccbc7938708aeada527bffb57cfa208921fd7f04bf309cb0b2c4f3b6a4812eb538418e73ff2e50f19206813f6d04f8b7b7799b85b9f2268a8dfa316f95a8d2c93c333cc7ca4cf51ce8af2de4290ce9a878340946712320565857dad4bbf055b97dd0262d54243435fab8b4a5f9048054950ea508d98f6dec4259fbf4696779bee0bb6125a910d8f02e8895d0717e8aecad510a9dd007b70c56b31c24b7493b8eba8b4add2bd66e32ee518893cf4657948b7a88178bce0f573a97fd5038679f3c71e98a41c39ea1996fdb4b759c222cb2af2bd09a514b9986c5e1abbf1afaaae33393be4c51ce9674b2bf596a7322e42591add9e5acc8702cca68885d3c347dc688a39d57d9d812f1307ea9fc5fe626446f8586e5ed8a460f2cdb45e90e4341f999bee03b36e5b8d74d2eba92370a510949d8158a1968966d416e149de6134524c5542b8acc5c242c897b87b8132a41f8033423f8d652d8dba29a2893ace57594482965aef8812115e8b7609b334a51353a70d6affbac4bc339077c6d9bff0ccaefb039167e5ecc23f204510e09db575ed86669a0248a14e612843d401dff0412d2d274a210c14e469733fa6052ac84e7d8bd5baa1304fdccd2ba4f50f58c58b324e1d00736c32f46a6d2a1ed86719cdffeb353501486773c2155eaeeaa7a979521db52372faef9eac90f12c2ff7c68428dc567b22a144cd956cc6163862e10a0331163bfffd48808475c2147c72de983d68c71293c269fb174e25d5daf48c645ef7ee6ffbe2667d69c687b652169f8691d474477661f994a49b4fa7f9c0cabe1c16d1cfb9f35815705f4e895cd9ed5e372c6ad8fa52fe3dfe1a07cccbca2db0da3611f08cf1a25dfa6336b29d4187c3a9d29df01cf5997458c842cea1ab68b491de5994b5f873c618dea8d05d3a1ad96805e65e6edbf71956e3bceb7a84df1cd99c106904fd78ae34488897fc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc3109cb2a48acf770b6228810785bca168f4ce7c1bcd61f22b5f2cf719dd8eaaea50289240d3aa509009b42aef8511ed10c2a89dc14be7037800361e3be17dad18a5318d9b5bcc5db0e0f19db5e4e77191a844f199b1c4ac72bb18fd4978b432a7198357365bf51ccaf6cf72be6f9a19355affbeddd84a2908096aae3e280fd17686c71099c927030adb2e78f7f891d0db55c1ec3738ba808498b11262f78245bbc3ca1369a5e3ca5b8e58d4669a645ed74ada5c9dfc80f8e19910608dc82bba11ade0b96320c1f78c7c507c616acfbb38414add15545b0f6e4e5230caf252da023e028989ef1290a31dd052e6c3efa6dc7667fa8ddbb07f712aadf7ad57f8eec4f328615d9688d11c8905482bdf0c8a05b5911452547dc85c51fc749ec45f8e77cc4ebbe0228054f19e9f8f117f7d25ea4f3e315415a89094034664ac36dc9c7a02fdba65dbd48af58bedf6a7e46470c45f42263601794e929a6f8470207b846c081dfdb1610e24bd52c78dc27174333af5ad8eaddbaec1080b2f20505d21e40e0ad36f312d21e80308d44bd19577c6377874a181cf08f57ee2012cf3151c29e9a6861cf59fd60aee1487c11a6a371a5bbd444b5c1359e1de831aa567dd391e4fde4be6ea866dce835a1adfac02de00e9b78151a500bc9df0cadc405f409dbd328efab516b14774c4ce9a575c3f1766ba7ce336adbf3a75b5401fa7d32a728a444ae1378c013c99ea67752d769241eb31f70cf9f6b02f6c909915dbf2e037017ce8701910b39579c6aecc220fa4d1af06a80d68dcf8aaec081abf45e17093d77e169624841993071765010dd813f08c4ab591f2b8202592be79afcf65db0e1b06f4328783d90069713fb56e9dc2c2a07f1936a803992126f427f5861009f155d69e6cb236731cab6cdc73e42a043e25bc0f60e07f6789631bc58090e808c3015429abc5605e3ffd86813fc9c44710b74e186f15d304dceb77077d8e3c5819f6bac36fbe7f2fd24a117648f8fed7c6d78f3db4b5f2ad251376dd55c7e9fc2106340ad6836bd67af3c809a4393dd44e8120f4d742274ac02e786bff4d2141fd5d0dbc8c79c13a338e49da0edaaa62730b01441771d1ec6604660f6090229107e2e1a2d644185c9c605f050da30a7b630343d89a9e334120545c64936c12c808b33784c28f9bd8ae0737d544451fbb5a1f337d2cbf0381def18be569c167a7713aaea00ca0b4a2049304257715a32f769ecdb5a77c73608bc14d95c30eb47bfc9543ac5696b371715fd66b99f953d85789bd068693b7715f8649891ae0cfdfa22d535bc65129f7b0683bde0aa36ef40a2edaf4d1e36d86cb9a0117bede3aea72616d50cd036a94d8278e49a94a5d2902f66306eea5cb470e04e93cbb51e61510e56774a6cab43a89fb281836f4f7f080c813477a513b447c44c292d8f528f1dab5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3087da866f84b2046aa1c19c4e64aec816867b713eba29b2d5474c37447ee6eef210cf4507423de01c2dd8d4a8d6afb154f24d88ae5012b395cb26c2d6cf6d6f0c0b77ea7674d737a804d7d491c143f2e4af98ea5e81c93e125e1059ac928f895d67da70c6f38e6c6eb8f477339f48544c9393789be019e399691594c5de28e78d5210d2ed9c15257dfef5e535b534f85f6a375ece0d54fcab495edbeaba20c1860796ff3331085a098b0275d2bba48c40ddae26536d3c10c858bf9da446923768e9ec585a52834d0ae4bfe7b6be1fc1a909205688aae6f421f40c549e6b9f535d3854e2ae4fe3d123d2c0acaa3b7f11094a30d8b6730f4dd5fbfcdc2fdb6c046bfe3968b5c7a6c67b3a7f0bbd696243de2a8fd942a783cd7e6edc5aa81ae033fc0325461cec50a319e2de718343c75840655c090b976da66aef0a6032f4a7cb99d0ca589064f99a8380ae323097fd0a8e5ad9d7f197e3b519c2a2c52530a87724b7be992b428bf97bca3e4b950193c545befbfb7344f9fda717ec39d4460e67a253a38a56ce8eb58d476a3c1f170593c31666dc2256fa818491ffa370fa693090ec13c01c2019804b26afcc38658b93c131de381320eeb99fafef04fd55acc64311919328e31c3ae23a4ca960bd2d9092d2844425085490a0952f0b32ecc772714f65af05b2d1b1c3c6da79817f830258a930c6c608ca3d79f361491cd5dd5c19a8afeea9e4ec8dab9355d5fb1cfdc9732c3eca336edd83db968b58a1277cbb7f43e381c6ac308af06a784f6518455f681b47f049ac16129f5082e1916d8506ef3850407b997c7c02916de9962ca4a8a6ff9cb9738df502ac363921b9da8ed336c9b3d4202ede545b8fa2e8bc7b62213337b13cdbedc43b445f2211e7f24ffb831fb541f2d1c8bb7748aca96c60206418a7c8e0e7ef2872b90aa413b0f25cfaa96129b2258de90a9debd97d2b3c76c2b7fd2c7880c90e65c7052e2c3d95722d66a3394b85603edd1f55314bdb5832323d9d9d13cae381f5361e6ab624d7b0d0a2b0aa97e499663a6b42534eaa8fda3d88cc14ce84bc01938cf1689380b4c2949a9f0b0a8247b7cb2a0b59b5abfe761c5de474271504d55a01aae51ef3e432828efdb4309f9cd57c08a2b38d460e7e2c0af09ddea2de664e0eb34293da78eca0e8ec5cd4940c1500301dc496ea2abd343122b2d78baf6ed98a960d64b1fd9b4e28d7bfe2b72648cc259ec8f2f2fbd4f6d1b675625c71a36d39f0fe3b313af2a6e6f1ada9abb036ae105494397103b309d5664a4e8cecc8e56e19c14d034572f00c128694b55f80fa7638a129ec21e4787a8589d48d5210a1d4e57db389a95a97a2f20ecffcd4f1f42fc5a057bd30781826debde7f5c1ca333a903b6039f1c369b3324c4e164e2f37183780a2388f63d3e47f9d25565bdf21d235f165a3ed3cfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4050cf953a67326a11b0c514677cd51b6d0e27167ca48958916c0e85312100fe22b2b9d0db51cc5d0f270aa42f4e5b3cdde7a83ca82395aaf98d6cd00b31de7e00a39ad11bcd494fd469e05424e61b85e91141e46ef2fce6dd91d091af52b752abaccda4480b332cc418a65d6340b86fb8391658636cad3b52ca71bae55f585a02c425dba8ea1e844be83d1c1d2ec44796220dbb726c551be9b1c9977d54a821860efe6b0d3623617f4d77adcfd72ba6abe746fdc2142a7981eb9fc1ab51c8a331deb93eee611f90674e5c47c43cc8033b81722a0e9b55cd76f215d44723f2eba9074c0fd019f5dfbec785e3ee057de0c8149ec97cd81e090c9c0c25799aa30f0b75dd71439ca61dcd75177025fe11f99909d5746181462e85fa2699d909387111d1016decefbaf154dd05206995fd873deede4ad173a7b8a33fe33dd0001c34f4a6f00a11b501d687fdc27c84b8924d8020a3dc2a968639a2e82ec410a9ea8dd264ebbb74ebd6dc3384ed1e0ca7251c6a8561cc7f26441c3d86143bab842f2a41aba0bdfdb8fa32c312808ea1d06d3f3bf095d6cfbe22b23030ada792dbdd7940df767ea09fe26348f4d2683479d3f1860139231577baa3df6e61f8e843e06ae234d9cd1d5fa133e2d909bb27f46e2c10177a92df01f3b7780a7f5da93c167b1904db775da7bd80c49f7abc55dfa3adf3e618af409313c0a0ceef65293732e013c3b84fdca7ff67e110501824dddd811280083df564158073e2e19c7bcf501afb5847e601da70df6cd818673e00a639bbc2c72dfcca66ffa36d93431b9870e798c88d5bd97d627c293acc8eab7a22a0b10203b54b316f2071a9b87c4612b44274d40e5587306596fb2cd172ceacec11b2924e9794bc5ae2d7912dccb1050625f5856d09ee89328be68baad8e4ebf3c91c213404198b0481bd49462383c08a025f2c3b61f3137804ef985a87e4c6739f68e3c1d14f49e9084faece1acf2111dd4828ecf282fe192e766bbe5a037715c64762b758ecf6a2ea0bc7d92671d0bbb8b42925d075ec114c09151145b78290a4ec2ec3e2657715b7251865b9f4fe1d40339132008b1566f236798eeeba5c6c296d51d214da1ab78eadbe7d265ca4bef33ea662bd29343d3a7f2fecf32ec968472121f904de3fe15967be780ff4243dcd79a5b97f332bd2287110e477ef5f7c19a6f1acb49f41cf3679a627eb4ecb866c028e00a4a2f85db45aea1c745cea4a86bf12ddaa947724772981de52713e3e9a6ba9a18ec40236349057c519c260ef2eddb5f93af524e75d0ee8bd402e76601f7d1d8664f034880a866cdbd35708d9e18aed580b8332c69968f6da733862f52743b302b5637a2699a33934fd6d87a2f4f4dbf42ee52898ee68276be691705f09c487fda12387a7f1edc4f713e8e847561548851153ee482a80267bb01eede8c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7ca0356f242e9e8f0f4ed004019011dcf0ffbe445f64d344a9acc3ca1cfe7d3643b3b1db08a2e5d4177e37d01d43cadf6c727f9eb9a8fbfbc284efb9799f67a219d3396117c84ce153b91fa945dcdb59c66940181f70dfd51b08138aad0d3f0a145b5e94a95d8471fa285bc861522caa8ff4b1689b63e2622b35d966e44bef9c62946c12f2593da30007914b3261ab39fa4404fc29059798aa7d0ac54b083f5ae2beaaca95aadd13f0373e1d5a5331d6316c77cd3002503f4135111bee344e3536f0812b8fd97cdfda5352346dc41a1bb9e2e7fb40acee5bab73d4aa5a318c7eec042e7a9e60e02b72edf1f0e8ce3ee87fd453350387d2cfbc39d814b42ac668751bf0e73f79fb3e52df7e1cd081f05c5ce1678199116bc20c3ed3dc6b3884759d20ce6a154b4790f833281c5eb55e2d42c77815333a5115b4c48f45987d9ad31b4bdd448b5c27a08c32fc3f775508a8970f7d73cd7a054fc6da7a989b1f3cb3f9165ff9789adbfc03ba9007e3c3010327715a8a21b3d577369066cafb2c2d666e8be32f4acf4d9d927ff301e179253f30d79f490b1cd29c90730046caeac0f21ac5a325049f727e8f74af3aab7cce8958531292f92a30892d27917de6ac1728f1154f1d4415f8ad1778350b7b32d52713cc3535cde50ec63d1dbd17d9ea890dbd4dde1c469cbde126a07b076a9fbf179b730cc2404fc4b643e3e2a54a6ad674483f921d206b42b8b2c86ddb18693fab69320ecd023c51ee94c5f79f349f002d9facbcd149c3bfe872771a14ddfce38d7c9ab5d7970da9fdd4b2f123e94dd9c767d471c00b5a9c9907faf0479fc8663c125c45819ac484155055a4147b4833b7f08ff94b3471eb9d2ee0329f17fdfb19cf189e2663bd02706ffbe0587c3b929389e32dab399bfcb8c4fb99a44dbbf04b416e9b053e30a9508a85cabef6a5c80d402a16c01be544e6689721c4829f23510aef1a5ab7f0171fc8b7bc3df3f8f5cc579c04f670344f0eb9956255612d2cf8c3bf73f5da56d9c7c417cbdde975819646a0336b1bf4c04ecf9c391c29f5a3b65c3ae027398f6c2a6a55baa573f74c858efe34c57e1361502819aefaedfeee1979c53ff116122fa71c92732883ed98a2342b43f4c2858f33cc8207d1926db9f2eaa4e87624427a06ab48f2a4e9003a765c9a5e525819ba534a7476ed0f296024846be92cd951adb866ef6bbe9c5e7ab6ebf356fed4ec1a0fad25186c9314ccb996128f80d8b7bd614e6fc7130fa99771e27d5a8ac9e7de0b20359ee1600f4367a75241d82143fb3dc408a8f1d413edf5c5e063cda82acecb82ee1d3459c35ee43fb204c5a27778205e0aebaf137f10ac0cc2c3ac9983f0da1c924870cce53e12cbc1f2316643775c11d209b9233c724c76b175d25622a1124022790008c682df707128add3565a1c295f7679311a876f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hec2ec72bbfc7a2ff7cc210d8c129c6106f19601cb234ca9dfa3d41606c2aa2dd20dbc5dfe38867ac472288d196a7580bad27f2da4ab1e4f533ad457ed72e02f0982f2c55d5569507df8e6467a487fb106534f034d7c5c68d12ca022c6e0d7157c0bc4d04a4f797b69baeef585fabc9990f76a790e6d0230e6c5979ba7a860a3c6bd480b4869b09158aec09061ca5076b6a736a24129c6ea066fff11090cf90580e0c1670d5b081f2a9cd160d2181f8d6584ad558186653a7741bc7e248fb1cf51e43ac7873b0edda7fba30df599c125351d53614592f8d277f00e3a9abba473911f8232a55061515ab78e095ed34c3322a8669fcb12e8a9809b5852e0a72eb918136698e45cf3b12d8d0755dce31762d390c2ac329580d083f3f6caf78f9e1374ee0a239a7d8b1f28db847fe26b89f1ffdfab9e6eeed76ccb3fb1873fba36306d2a7487d2b3b6ba201a69880b2882fa2c3561884f5ca71e5099c18eef3b5e562b10e3fb77c5fde7e0cdcaa9009e2d3b0a09f3e474a57a02cc3e9dea97eb82351ad35d961d5c49a6f71696913bde80ff13ee290faa032584432e10abde6ad4f5916b13d63889e56b7ef96a2b1359d07dea47425fbc1d7fbbabbaf9d80fb9540322e2fae187be88cbcd1bb5e077d855928c742c2cd776e49f7cc43ff24c73cce3f57d0f9af3d01bedd6a617bc1f95b91fbf8508866b0442e500943375a05223559384cead6bb08a2194e02a25b193a8d6225fc20aec6c5835d35f038ca9bfb3656d36ab03eaf71d52b5504f0b110fc25ab375ceb522338ccc3ccec9883b96a9eef062c7a35fe6eefe6f869167a2303473946c4889f97fab0762264198f09540f39022ff8bf32b6d7d6c832024e74c7c863a6999a44dab2d097d7dc8cbc14a55858d2410951f40d322c733866a79cfeb577ca5edfb5de1afbc442bc1ebdef501aeb12d94843b1f9169966006bcfb4d1c78cba52ed541d0d471d97dec52ea07adff61b00c0ddeec75e2f18cf5db48feebdc882fa3886dfcd1e82387ed9f63b2f9d91d2f250c6ad705e9db0f5e9406ccb4f8d3ac52abfdb8d41ac8844789b06ff11b992eb701df22517c846997a64f0520ca6e39329cf5e1fc2527d736543373799811b63587c915acc32ba89be14e21dcacf15b75ab8a6b09e2d02a25632faf3f7f5b9685d30a1da0a84ede8a1f8d744581870ef35bd252bb0c415ffda6530c86128da13229693d317ea6eae2db55e6cbedc7ce83227f89b5d1b4600200b71f6242a3dfe1e71c1347ac8b4ac692771c622b9156c9d06ab69e7facdb7289b2611ee8a013a3e3d13e9936944b5c1992d4e15a5fe2aadec24b767062c60ffddf69d76de5498d3e807e923fe4450b6a0d10e08463102607ce77a31ad057417e51e74b67c23a1a36077d8cbf0483472d98035d89f7ad460e958bcccd04b8c18c4ff9efc2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h234d9118d48f54feb4ed51a5a55e2c4dba1cb1efedd8a15533c25fcc519b487e09cf16554c39bfd4caf10a40d08f69287c8a1ec3af7424122e0e002225d0827e46a502fcf432d13e82abcbf8b6a14da2f81733a5966c61c7661d78db75417051e9e9c92221938f4ef30af5d3d7b2832683a0773670e58b6db20d3422f7be43dbc6881ad39b69e377c5d02303a09c8340abf1f2455e0ffeebeb21d85fd83f52ad97fdc65c54362f44d5e19f75ff70eb2cbda31f5a81dd64944b792fedfe6deaa0775509be6cd3ac78b97d444aec2589e633980862c35de29166ef04cfefee3996d8cb31e55922841c23a114a07843cf00b1f6251970c6d0ccecfd175bf26ba7a1bfb3cf79d42597728221edaf0e6c1b8cd7f317a21d69ed7ecccec8567868cb28fbd3ca546c70a7afb204739fb64a8e435aa6628506327f039995c8bcb2128d49cb07ec766e93fb717df300b151838465d2b44233a9066db4a71d4e6860485ef55a1c74080b64e5e9b5f8a2fdbf0adb4e3125cf11c7acc30eabb58c002a9328ad15a9c0dcc3795204a6c4afb026fe4bd55606ab1d9d0e801f340aa2b0f81c12a2956bab93dffcb445e783a09f2c64cc20df14138a5cae4d82a600370d8abb6fe2fbd641865ab072791325611bf7bf7ad7e33dc53991721a8413dd9b3bdbba5f598ba1ac13c7397f41d7cea7dcf86fd3a91fe30090b084e6d643d5e7e49f0fe31a7b94179c7800978466656587c9496cb9e3eed740e4ce58abc414b7b1eb065bbd81cbde5e3b7ef97f89b1934fb7522b262e2843ef9717e685ddcd3f8f087978b456f39bb604a622686bca9c695bbb1b9f3740e5079e2527f2513d1176f0623c108ceabf9eba6b33703e0b5029c926f8057ef842a65e61f83eab2af6c801722b8064dbba2ca7fa8c5acb1fe5d3202e820c7e1105b1cbc6b759d5ed45fc0ce49159ca500f2523f1b06553d8a8d74339bbee89b491ddb1af424d49600bc74d32e4ce0001b123bf7eaefbf70e05f8341e5248dc5311994265f02fe8cc5a22ff11aa661a94c7d867d48342d974d45bc300a437d3ad289b8ed63eb86dd6a3bc977b3c992b7efdb45630841b4181286979bb51b9de8b7a3b34213eaaa158fef307ccb6688b237486fa266240e8141b7eab4b9b75f5177ea8218105d8bb83bbd168dbbc4c8190b8ca1adc7813279aaed3ceb5e2a495f6994d36935c8ee667e0769805acfe3b26aae1452882b6b306746604c0e0ab4739a21cd6bab449aa7ef1307d5df0d643ce332af9a6a1bfd24bbccaadadc4913d86287ccdccd8446a9c475a50ed0ba1f5a82d84de3cfa8f92091740992fd4b9a81bf40b15e50f14a7350a93f7d5df3e2c9ab8c6b373cb58a36bb8226a94e3bd10bef37a36748690e1e9a227a6e2391fb2ff5b567f113f27998a589b26c9d6e2e477bf5c3fa22f1af40773bceb60c2bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heec35e1fd7b280b2cf35e17a90fe5e0fe7d944543cd89d02dcb25c2e10946b9d2801acae52664d956f8fe69abfde1feb59950330b2913020cf78eebe63ac1dcb56920acd00c3531ecf94afb90f78ff54c62edc5c222c4259bcf868cbd3d27e2529c5d5eecab9e4c6ca7237e9619a2ea11b6edb5e0fef9a8ec20edc82aea7ed3fc8c7d8a052a1fd2754b30a1787a9eb968458275438a5de014e67294a1a38af43209c1a1f0a67c7d0032b5e9d8843098c08b318f08301a36bafad53deafb1b3e6c88153e696aabc8c084bdd4adc66bde5394881599edf4fc285a95e5fa846932afd6a55a3483d72058d5d09d6e2b614c3699286766d68b8c03e7928fafec0ebfd5303b31805781b5ccc44e85c3a3574e2a6af1c73a4aba18bfa6b6ba905c53b24f686aa1d23483adfcad09fabd3ef8bec55669783ca3278496e5a7d2b1367f55b9e6d52a041fa7a1d1bb95ea02646ad0dbbefd66f2fc8ccfe6e1e2889b7a48aa1273baa2cf4aaa1bca4c4fb73d24bab74a5e3682e05edaad21e850e10ccd6beadab71fc7b3446cf823cbf6cdcdc1a695e1ed7d129b55140eea543bb54c463ada1d84ad44bdf433f0cae942d84eff7cbfbd32ed354cf888ca068dd34aad66f73c9c4ac27718de3eb7844079b3d7da7c4d2f923a8ac2c076ee09bdabe54207a4309c176114ea32e2c3c9b54578a82eff1a73a9af20b315b3e4c716e3e5f36853fc8ab5533019c40db11964642f1429430579360ce21f6292ff5717fadd4e57554b031777892a8eaca5fcfb9c258f564d234a30a8985d713a8abb3828b5ae6c5774a08b3c208d2225f634ced2a60ffef3a982cb13b8a7d57dedd11b9cd1e0dd43fa47809fb1f26bde33c965edfbd2ef4256a90ed2a87a5199282671dee2e21b292071e057cf43b2475a35afc6b453c2e7d412968e8881c64dab8d41fecf5f0d71a8368856a7901255d3c15e2013ec70015f496e4893c5b35fbd29fbedf1c46ef9ef77002e8f3037616057107b6965c7e91b8d2cb5af34b32c11a21fd7b2ba22c76385eb421be7f2aa396cc1547108b2750a82ac7a54626082e5caacabdb5115b840fbd28c1c4caceb73c8576b54cc5f4619dbd58af852dda286fdcc582bc43abb12df2ef4c1d15cab3e8ca30fce14aa16fdec2a31ec71741c27cbc6bf522fc567ac64b0c15708fd534e1ca24aad0a7b0935a7f3195e3a352095e21e8bd305b5bbf3abfc0c51f5deb8cf8f25796f1d129809b5a4d4f07e7ed4201b9bdfcf582d926814f87a50a8a51ea16fe90c403f3f3ed74120ac5e0c81f9f523a2de2b27cdbef7e808f3f6384e70c16da9845d0efb86b1ff5f88f68281ff48628cfad8bfe18b75d60a5c0411f5e4421377f9a0f13a82ae385357d2f7f06689cfad874577973746f30e94ac52e5995bce50a333b4ebe2c46fe3c9ebc803f852e00b64d989b8919dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6b9a1ed5ce85d60922f66223b0934bcf41ebc04ad3fb1c9228f0bb5dfc094a5b01c741b67dac0f4f166474ec062815de6fdc67c92cf560838eeed648efdaa9849c747d93a38df277c9cd7fbcb6a0755f3ffb7472aca925e0ec76105d5d05d78aa58b54e4d3990581f2b39c24e022b416df11b0c38e7157993d9655339da58f45b9064d568fb835e907103cfac34b6563c5e6eed21a22fbf4ee4267c65a992e01525e805a8fc328794abbd2b68de08de78228ded624cc3e4f912d9a4d59a12fcaa178ff1871805b225eb74fdd13320e5a839c5cc0c1e0d4237b21a594f2a64a9b4d093ce3288a502fbeab765601e1cb955ff023f126e66c36bae68cf193f82de06e286f6b477692ae369ec5edae429ea05ee6f1b16c618208c3507c8b177887d83b5c8d5bf529029efdfc52bb0cf948229e081f2cb0ed11fb37443bac4dedcd2cc62c545c2d0fcd9b75b1ba4d6d8870629afc5481869424da96d7682e7d51489b15a20bf11a9c9d92beaf79fd332815f73247c0985001797952f0f73e5142f6e428b23bbd7bdf17097bb931c23438e07897b9b3c6c622e04e9963ec6933156cd0a44964181d0f0d637ab491811d0117910b4485db70801d781dce930c2ead19e8882d6376c0a2b0a33f5b40c2901473ecaa1a23e3c22f47efd6a31d37be63108996d23ae4b0ad153ad47c4a4d1edf48a0bd3ed5378b3d937fdcbdf138f4e031ed53c11e3ca9c5b0060bf2e08ceb13a3c7c47331da98424ed5eea134349e2ef4f43e02f82ebba3f3c9be211ccdded8be09813d86632083b807bcfe82cde66802faf5b54ee13c84abcd33670a87cef7a13209e839814a72de8c2f32806214ceee694abeaa9d80c986261e68c849ca16dcfd1d919bd441858966ec7a0a067ff135ac9e943d858c7f19c8101eda3dcbfd82948a38d6e3e2a5c4a4458ef827d792c590880ddb49062c9f11eb9abd6ee03a250b289efbc8fb7cafa1d92d0b3f6419a1145fe74dc4f06ecdecc3bc981f50b1daaa04fe6066efe04af91250b91765a7635bfccb514479f9246a3e49fcb9ff8e66d21977a78de8a80ac71ba4fe231f367c3523be917986f814ab18ee309b32fb46ba473bb081b37a3f73fcce34b36ee649d62a10a7b23aa36b63b946c4a0d5886e1f19d86d6627e9939c514b600de2836f872c563065112dc545c5fe39165c3f0456730bcefeaac60c3b5ddc78907a0a484ef53cae535c51e61340c056770cc96e619d2d7d85179cc8bc89470fdec99ef0f0fe17ccd8a2527646539bda7a78e0ea56b53913a9a3af609a9129d591ea86cdbb039a3baae1b3669129d8fc54f757823763c6637a6ad1c793e52123e830a403d9d1e33f113688b741a534b5c2b6f6dac1ef437e8c4ad6a956667c3994b6e073f656c4a0f416a0995dd32ccf1d6b4833981e198df273add1dd6a7460953d269b9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha7cbe1915c4cb94fc746e474525078a92d0fb6833fd533d50b2c5358fcb08910c098af0ac294c5e5ffff170b0e8f4b9bf7c46d4b8abfd20521ad03c71d99bd337576171e167bf520ab178dd9306cd0e4c2fca64d64789beea842b85d215000ff41f876c8a3989f0145b5111113fc383344900958b3d154d48894fda9c766205b6184c588ae11a67b6fff7072c113f13a998c2f7e53be5c92c3e08b4e0d1277fadc47c6a0cb5d4b72ed104d52974b0cebef71eaefef07dc2609615a7d5653b0176a5afbbba336d38ee3d0368dd1acfa5bba29b5b6bb82791f2b445ef2d76141560c9b853e66eb05dd6a87237daa2ff2a20303896cb1024286128378ad48c9533791e58a0832d5ecf4d93a7f4364ff82fa274d6ae98e420ed5033f0bd89bbb7f4e397007668094b7592dd703f9bc5df2eb128024c1983155ad0bfc8180002ccd720259ebc072ae3c7e568d9de8913796d1c2105d96e5a1211272d3236584fdfad251da3846bf15aae78cec96158470d540fbdfe3722ccb5c5a06b8433d24f424b9ca3f701374c1491ca5ae6c033a8bd8ab8b287556bf54d5bf37dbfea1c8cae13185ad3cea57fa818ea9a96a7bb9567f2242fc5ecae26d2afe38bca5d08c99f97d4dbea07acd8540e54dc5cf94759fdbadf822621b95dd93e21bd380a92b61a9dc3e17fa397518de273305fda5c653560415c7cced4c5b9599935a217f61d1984899bb230b0ec3511a8e64305551dde4cc29299c00c33eef32e38f42ad3958678e8b2d3640bd5f02b640acdbb1cd1e59e95c8044ca92be0f90a247fb11ee57520ea8630a958e67caa3f506337240fd77392e47bf2bb091f69b695c4b816859b0435ccfaa9cc5decef8b9d565da0bf9cc0bb504bd8c42a2fe908e115d7fb04078228d1f998755cada5619419e4ffec052705e7931a1475e6d78b03eafc13da362ccf090e1b1a36c4303c22e73090dbeb0c115a1d07fd5498527f99e4d237a1204c4214d852b753fc4237c5375b697ad0ea8ab68c88c12fc913ab20ba04b74fc9758d98e19ac2a349d08225c60acdaede024e44b6452927823aa96c01e9fadc347df840b6ba1ecfce4ac2c4dd86eb9f7542d2274532ca8cd85a8a62395c1e4776730daf8473d36723d73276e2b8e101aad0ee73207da402df433faa22ff8d26cbcade5c4cc33b14d99eb6283f6cb18bc033a8714694cb55e6fd14ab8f38b9607e31738eaacf73c01aa23e72c49a08e7fe022fac5142be24811f3357c2b8f47cef4076d2c1efdc18691ab32709bb61ff215f725053513db328189fa424d00ea4c6353a6e608ce2cbe2ee8e227a98ef52b48d6763c59577092a1d291e01809bdbe606ea35095113cf87c55f0d8243c488050a7cbd207018adaf197f76ecd87f96123a3325c309ea6eb4247b8f64faa8d2624498970d8f70034efc763215aea5044451f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h89f2410a174b18399b4eccee75640c839e5d20b324b3c5f0fa6a13e9c06a2bf92d590e78285123ba23d6c589f0ae3e293b6420932c50ae34a67fa61cb751ccf90821d69af062f965943840725a05385a86074f7507100790c45d51ff2e9a8d94df6df9841d928616512a54af0fbe3f5e6b601108f0a4a0a7eae8fbc650fb60746161e9679466b614ed39c33e51b125c3bde0c0d40151f58edfbdb50da6069dfc5d785da2afc54f9e185577825991631ec37b38316bfb93823f5cbbe18bad300d6dae1134074254ea2a021d5a55af47c2e89a20c086369ff2b676abde8b320314efcce4c9f91ff260f9e4433f7c321e409cdc9376fba4d9e6f4028f2bd88f9aeb94bb8ed53315db485e791343055d1c3d349546e1feda2370f55c0a256da6262070e832ecb5291a72b9e39b9b12b549f1ee92fb8be2170c53211ba9b348194dad04a50e661f348518d21cee471c82799492250f60d4ae72f5d67517871c106f4d6a0cb680886d4abbf8b1a777f3fa9c6aee2aa5a2c0f418000726ff461727940095adb8d5cb9f26cd985252346aef7646b9d884669a41960d436c31442ca4784bf04c075ae6c88a7ddcbbd860008a7f0dcfbd29d36c05c49b5be4ea8ff55b81642425932f3c7f6a84a70a205b949064f9448be053adb732ced644af5f087dd4c787b50cbbafb8739f7268fe12731ad2410641247404ff8a63abd91a527ad0379d8b3235be192175116f4c37b7d7a0e73f054262ff338c452e02f4eecbf1518ac3a8086f22543874bc93df54253a36370a56743811c348e2e28a50d5a4333972393cf3ad8b8bbfd9217b7c1d67a96ff100addc8374655db57c1ed81691b1f9de07851cd33bf685cb623cd366e0a93ff71c229c2290af79c6645fda906f313e96a2752c24249fae781265afb991d3e0a195645414afe677651b9b57bc391c3ea162fdf30284146e7e5c8656d98ca0e1322f83fa5971d43bafa1b5c772066a4bf90bcc2a12bb452a12ffd1e2d6821e98ce9b97a1853693cdeee850404ae262a2ca509b26ab8e039b2e0792d93dd2c3220e1f9e535c7319dbc0a0974d05f8c1cbdad145af311a0800e6d551a8a30f2c736e7fca80a5442f82b61e9a0b40bb7e5fd978926f95157ec1f02d6e721c5180037561159d5f1f005caad229c11208b9302ddeb7ebd898cc4d2d1dbac2d31da6bde74c9681dbcc230a8f24ea18dce622651beb7d204cd6a3ade72d39b29575be1255932189c0daa1767cb4e58b95c7056bb1cb88228498afc2b0cbb4739dfadebe007581514a40ffd7b96075e804176bc45d505e8139f61a58585138f4682c7fdff86b277864b67fe6fc0446494838492cc4c9a430e7053740955186ef74e30a3cb78c71ceca8ca56f5f0d81496fa6f20577c7fcca81179226e820005a37c7c6ffdac2d8f55581584797c2c7e9ca558313adc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd3a336c609eede1fc2e12d9f0bed346fbafc6c60eb372be41b1bff3d80d79289006e8ef3997d1e0c034766527c7816404dfda016b06f6309e336eb1a844a9ab80c5dcf65507f312a55b0327f48b364d666d0a9d5184d26f847788637cbfd3df3eff9c8e34f7e2091a3ec5596bd32d886c76bf8793e36686ae2964704eef4a26a3dce9d1153cf8ce9d680c289c3b4b87e94afb045ba371eb79ce1055cf1aee318035ef87d3b6d51b260e00351adfc19487d4baed658c01b0a96c20b1874e981619348effba5e47156a6e4b49dd50dde770f034dba4cdaa9826fb0461aadf314d169766d2fd3e7ed669a1af28453647694f4e768e0a893ca66e3f82cdf144ccc1c57a808e058ef4f3675fc3abaeed154d2200eea1ebd5ad3b3b4f482a00093d5a90ebdacf360896e35dfe996af0e481980994798e5eb5ae5a428123b9d1cf5aca72bac86e2dc03c4b72488ac53bf56e9727656b0df3131b96a73a96af81e13aa3b44ccff78ed99d44ed5f3d222943f6f48944543c41ead8f09888b4814b7d435baa45bd3d7108845e00bc400aed5dfd6d941e691d7ca0dc03fa73cb59a8d0ee536f0ad890bb557ac9218c3d59d437cb1662bfcc41257589fc14b98647e57bff3beacbd4856c308691e824704826fd2e638f8f9e9088edf9da2722d994de03e0f4f490674b1b677d0c1ddb920ef62525dd2a29095087f5af215be0ab8bb0632d68317c452aa0b969929d18dd9b368e2a5073a586e7c00827fc7547d0ed55f1336f8fb7ed041031fc78f1963ce59d6ae013cfe2e2b4328421660473ec869649d0929465a1f6a3350e49834674026f012b53e9bca47acfba8a7aff7bed53f9401964428bed9f68a64612826010c9437609d212c5c1fd9870f09f8e70d6b4b9438497d91f53b86c62aee4b497e8280a21ae1bb213a3fb6a698577bf79d8fe0fa80bbe0ca1e4bdab610a3e6d4cd5d1fe1921af17576352ec6337b41e2a5bf1387de4cff0a1276366056580c555750b41e3ba3fac309a0e7c8e33fcbd64c41b9dd03f2522bf2443d280e21a71862178423c9a592c4eb38cc52754bf401c5dd12d71938b00c1b1c9b4f14155fde3631fdb7dd85205d0d62c59caef26772a94423ca08690e1ddbe8bc037d5c2564da3d5e32b4a19bd0fe61916a85f57e3fd8ffb9bbc991f16503c0fc8f8d4c9024ed3d88ae7ea08b2564759b3cede0ba610434ea5481f8108f8d9ccac43487528b2b9f8bbe917cb8e8f23ad1c8603251f7ed8f21ea633ec340d792876ea045624337a157bd849d3d1860070a9ac3e27abc10f013c9807d3495cec3689583da37e9088237ff1aba6dcb29fcf7d4411658f7617611f1ce43a3d8dcd8973ab30ab303b9efc3532ecf7742e5aa510eea3cfe16685ddb74512ca03146545c895594685609c12b196e12b115fd4fdf31f9e4b6eccc467cf966394a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdb8b01ee2ba20391c733a8198ffca015f0492aaceea9fbd60b8405704de8dcafa8d10ef4db3051fc1c4fb31adef1cb250a2dbc5742bf743267bb8480c23fdc35032fda2edb3e6a956fa45e0185a2a56de28b20622c7d903bc16cb5fcffe01a6393834d9a1b46f2ab18023adb3f26e48c0ff0de9b9ea59cbe73c013c02bc24311cee2d7d89dbda4ef193b4e188d08bce4157e7df129cf73a50a792e8c91e4a7388ebd466c2669b66da88ebf35b8f35c72a23392eb47a43331b622cb9817db44c849e9cff09297bda4441f3b518c038c9b119e251e4455128f5e7381d0c480be4b16a6728c7a11292d6a2d34cde965414be44bca1a717f77bc2f7384e96cb45f3c3dbd21461f23923a789902d4a74eb99f230cc9b3901d04544225abdee72049bfd976c98a92ceb5056083e015c4d442eba084a4bac590cb9365b6ef54bd3bd942cf5cc8202ca0bd5920a6c4e822e35f0cedcf3e040fce19dfe563135deeb1fbe45318bdde30d6f16600dab473bbd32f34c42e5feba2283cae69a3b3661d4e6867e1e4057116f702e3ffcb0a14432caa7b88cea1d4514f627d8e57c5e174fc5002872eb4c4c96a1b79d393d1673adf9273dc838eb20f8de73953e4f38f4eef8220484885d1ad4b842db61ec3f7a967e196fa28d0ec9e8b52a896f9635c333ba449cddb4aa16be96d1a1c691db9f21e8f73677bf59aa87dfd235162162849bdf7c19f89fd1df2aad88b21039dc78b0caf04ce7ce705be9189a7893d9732bfe409aa5c086d3c1195089fa898c5e2db7d53895d0ef65fd0011914bc646812bb9130c5d2fa339a232e081dacf4c04300afe01f8bfb113a31d5c25fd393ae3cacd1c6307853febe5ddc3bc7fd5cdafb4eedbbe78aaee164f7f37558370e2dfbbb3901d8278917ad577b9ed5d773fed5aefa101c0862b610a221964dc54363362fb3d605e0c20a60b3f42b5801dea416302813738882ce1767251042f8fb19a7ff5f6cf2f529741473f5f41e9e25684ddc54a7295405e8f386887fba8447205b99e0bf96c8164a97f8aaf0811ca5280367db0de7e293792e89bad3e0e0a28016d10b7ab8d85fd88172d522ee63d3b34120fb1a555d2608256fbd339f70cf7e5cabb278192c402055cb6da4e116036f934b205d6572e3f2898fbf046a1ba94c35a3de15d8ca3b7de2ccb4d90e5d9a3042c69ffa24d79822ba47600b16795693846bf0c17fbcd6c66c3257243f2f6aff0bd7a3f3006b258c61d6e022a42d2abf2bd24933284c744dbef1809e0056fd01cc872f426c75c76ee9463d4d6f90ef87d78889efe275adafd23b533e5fdd95383364378aeb678d6d24031106951446738fd01b96ef3e17d3572108ffc543f3060596a5990f10e9cfa7a46ff38131ba1dbf2adb92e6bb7aa6a00970f44ea11585fd9dab89918972f332776f1c58834eae7134aa87c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h930c54c0631616d9c6d7b58b6dd07c08db04fa93bef7397c6f609f54b467f1bb1407e571505e009a39458230c7abc403a4a841d31edf527ae2b1aafc7f95b578861d4ebf2f0c46e1241faf574a467468580cf515387a7203cfffdd2c95ae974de5b0f280ac8567527a7bb0d79729a67bdfa01ca06204edfc21f9ee72871972beb0e1229ccfac1a1e4b9a9ebda8c65ccf3f29da95ea2db1a4c5117f5f5a51cde921fe48ceef6ee686668694c5cb6459b990d34bae1ef3d1a12c27ecec497e017194ecd465c7ca3d846b4497d23b81f4b33329c3b6adb14ce3ab0193c2d3ee2a842d66349b5a97997ce7a2b0eb3d3f85de7deb59deb321db5d06d74e6837e32a26defa63979031f86ec65a472e63b90bea2c63f0eaffecff3dac9f6b0bc4c1a17210b51d23206698eca3decc1b5f2db7021731894f67ddd0ef8ecf53457ea9f5d9ef1e2dd7c0321fcddd5c88a845f3fc1bebc123abadea44db9fbe5b719ce0865f50f58143bde5f423769166f20747a90068a6653b91f1518bf67e175326054c5a033e36f533e1a3f5e0814fdcdc7eddea215dd1e0bf23c5a50a0669d54e40493415a42675d41afd9f217260e3cdf2adfa89d7ddddaa3f8700907e3746125249851826f0cfd13e1c63b3a710d99f1bcae2ef638aad5fa8b8ae5abf00ce52c955f3ca2ad21e2025884b32e5d5329f767ff74c2c161e758ca5b16fa1d94de3ed51690c4227dad5ef8033ac733f80c51f6258d3b09e0bf1a9218ae4f50be7d72f653ea9ad46571c6bef4c910ccecb4be18eff37e3a9f6dcb993cf0488aede0911104e668e98bc06b434fbd1702ab9f03a054adb287f960a5cc2bcb74a0d564d523a6c7890c5d2664285b71bce79d4c8d6e04cadcecd64638dcd5b9e9c973dbd43614cdc7c809d4f16081b65b8b94cfa095be27d0ee120ac6aa54042e8b857bd42714e9e4c54f721e102bfebefb32d7b4295c50730b6d7fc35d4c731c30dea2161c026b6038b61ee55be4b4b642dbbd13c6db2f839a038e4f95f5e1917e515fa7fead16e1ea934d750cb1fbe07818ad827be9ed4f5824ee0354998e0d76cf1d12d0d904351ef60bc18e9697a34b6434f611c676fd0f5329e4284faa35109b2c869e038298d949b3ac84ce784a8a90c5863f0e544bf8b85380b1fff3256bd928c10b336598706e5cdbb9e35b2f31803ac5c76746ed2b035572d66bf60af705610fc839b2355c11ccd01aab88b0c61c76fa0a17c0765695ea408fe9beff15b14c1b0431197a83c3d4958eb3cc9eb6ee931682f216d213fc0ce4753583160ab5617faee795e2e7050a0079ef30d65c45063365524e958acd8ced1e38a43f72b0d292c60c3010f1b77d8b9ed8b736ee41632595f2cc5c83bcd686904600e5652e4f303be885ea01a6aa7339b9b5b4455ea2dd1056f7fc9769d43897ecba381e4f0a899ef8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h41f1baaafad3a0e476dd4426bb106533f02c30bef88c4d5406926329a4efe06502d931324cf074ad63bcfccf16aad53400cd94f0c163f3b96026328673e62f02d386e247000025ff4e7ac8604e90675175895388da641e22d00a0196168b5d150132b851deb7f071c3f564905747abd9f5166b8734300e66ec85051505808235a2d49e26f3bbdea8ccda51ca570dd38f46af7638adf7f07c60b7c50bbce3dace13721edb484ebf52b5cdc7203ae9be555a4e1eee8c6962eb276cb593b1ff7c96ce7e893d7ff4e6a8caa584fea7685b13ac432a82b0ad299c2f2f758f5ce8baa8723c0da89f1deecb5fe8d5360d5cc9d817f8dfca6bc92893a29ea576e19777e67f2e5800ec1cebfcbae1edd160258002d240d5aa4ef5546cf6cdc6a61624d38aaf4801250856788f91938abb5adb2dd50f2e17a97aaecd2e95fdab0574cdb73b024b3a2d730fea437033b0637b35931686c066a5e8bc77e34eb6a89f98d277838b06a65abb98f412b5f81ed4e4a63e104ae134fc2da9c8ef71c6a30fd9b22cda57f6967c6e781cc287c129e1e0dd6eaf7f6d8dad176a645a5417dfb4081d31c8cd6dcdc70b4baeb07ca92b3534b89e477038285c6a26c55af77d3fdcdb02b6f7574d3825a618bcfb905c7e31e6ff9a055b666c9b90e9e19c3fd4e186e50bab718a46758e490c58e0230badb790edfbf125984b8c5e2bf92c6e7004d36df8965572de821ec590cbc13ca716e733c18436e9876aadb742c3fe098d9fde352e6c33bf5b192cde10d5fb86ae4b632f1c1f6f219723eba58239586a7bfa96e3db349b3437637d85a2842372ae91b6ff8ed4a65f2d5009c0d6c4b07edcde91e734dac3949d72e9f3ac2f96255fcdbf97994873c53e3d76f40de7c8fd9ca47d686f2077c999e4a7f5dd6e368bd4283daef7a2bfa7c0ad69a9f4dd9e2e1c8235a659e6ddcea1001af9e42d8cc034a5a226ba0ce7708e44cf5f049ec97f82aa8f4d2b37e2b975a281a5bde3f79484fde0cc8aa3ca28e2205455c7e122a6c1f6c5a09f043daec5a6b6814e3e6caa7ca7166896c24755840f764ba16b3b7d75afe6979bfeaf437d0ca489d971053f24569e904b496dff722f54797e78ad06101f4ec0a9ebc0455df99fe2b855424bb90f7f231f05db9e124520e5e18360af77f3caa32a194421d7b8168dc97812361d8edfcfd6e17ddef2c2016e2951151455a0bb0896d3fd21d30d1670c2498d2efa4a1245cb489c9c217475acffa13ced4b23f32ecfb7d3f39d76ed492c45d92acb3bb7a62650337d6ac99968f61ccd1dd5fd7dcd67f02dbe74e682f9a370454a49a787132c827cbd4120bba39a4a853bdc7a64e9559f944ccf5957b2a0052fbabe927563ac23825dbf360529f9a48ce0648b83b20c8b8a8e0230963c06ac4d4cedf75b68688968988ce0606b308eaf1b4f0a337ee3cc31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21f43858073c1c199a996871cebf3d1a2c2a7c91029ce3ccc80bcfd06700ba04b7ceffb6c394e99251d7266ba6dc9c043f2f72eac2adb224591392bedad4c799fe03656383c80f5d79cac673d41462b7042570a1a983bd9913b8894628e23568e13b5fd849396ac1f2b4a6d1402b501f0a538a64b1cc7d657740d78df42d13aab2b4454d2a0fcda3ee6f63b28874cd33653efbc35af8f8fe7e525d4fd7d652210ee023770d6362889c91715c3353e6ea80be0a08c40a72e687768f50512be72e40923f49325f4ee03799e89cf067deb7615728210c280c32403b53645a0745be28f2e1a96d68a3652387e9c5e81f95e933168e608d681d7f12dc6c8370a0e3287cf373216c35ca372f77ba13f3d9939cf878b441759e2be2a13aaa2e0c52e9c2d66218e695f42c52658dcfc4d0facd96583937ae8a257e57dfbc7db327b85a1755defe7671582277d4b9d6c823e484cdc2a10893228be7fca1e4a9049a046ece0630343610ec0f961fe086b2b8eec721ea5b466312e94b33494167afd04557c83ac0942266cfd0701facf25d8c0f710955049d8ff1b5b06dd2258fcc9d893a65925c4affe8c17fe69cae89387b117143184083a5e7c9ee861f8e40837882562f1c81ae6520be1768e61d3b9671513392f30a4af6f238184fa4adf55f6f47ca702f43f02746331cda7dc217a7d3aaef8b8b64b7c6d8d725a019dd4ffee4b8ca576bcfc98d105724371035ea313a3b4fcd7cbaf1d54ba9db4e233ae3fd63d49b42a3f59b81661c8825287a261e64f57fb1bfd95ab82266ae7ee8ca0a6e044c70e04d9cea7f4f21fc8d611848fecc64965cf74fe2e2423330bb2a5301ebea218b9de776083ea8102dc15694b9434f570b7f4912aa8d34a1b5ddeea75b93142fcdae3416599cc001268ee9c4ff00c8c50196576b610238ff43b89cf07b23501ebc81d4836c27557805d97e63b0826dd3c9e33368853c059d29108e25973e8e7f1af1973645247d9a8d8441f4cbc190684d65aa9fb79600b52ca3ec0815c1a3490ceea13db867d0e380fd7a976aa77ba1a3e18e488afd816e68aa8c0f11a26fc8b6cdb76a929a7985a14687ebe3978434deab883721173b14d4d21d523af1e1956e10768c1ce8d51bd21e375dab0d3d74587ec4cca821aca952463696907d35bc9133e8189d4e61013d960765a0688ede216e4d468615e701facdb12d9ff27625a36636d06048b475cfc44073eded611c29c8a5e5ae448c64f76058f36f6a60ed5bfe025d93ac8f67e039af8e738d7481fb367489de86c1f62935ce85dcdd0ff3671545786478f3182647c75c81d3dc9b7e1daaafc9ff1efbd265f446728f95d887893e4c819b08616c62c5de5b58581a7d8bfa61736bbb7c44ddf159b9183f293d657acea4ab35e96a33a4c69f4e6f5d3eb4d6a0ea34a6572fd67e30b3e77f3a09a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb2914609c1ee90c648d19bf14ecc289086d3250b980dcc2e37dd8426063c1cfb37103e000bd417285750632e1a0353da407768388fdecf420414f29756b8db012ce80ff270c273d8fd3b445717291bd8e2a25ce73b9d46768e5ea66eb795f9550e5df5d726598b24426b5b4849b29a06bf162dd72e949acebd369b52a9433fca08e4b6c8d8f1e79a712bf90ce03b8c4915367dbc5a983f548610d842965876292078dd745aed0dba4811c5d13092f322eacdb34ba78a8484c78c068e5d35b3eb1a5fb7fbda76a3a213fecbd3f644fbce86dd548d50c1cfe8ed8229182ee82f774416aadaf152a40c377c4b7c68afef2a3a3497db8f11c639e979f36da14cf5570ed12bfb8c2893c6b7e1a0cd9c9583e6f035e16c07b2f2f813a4a7d8322c2aa0e6cec23d85ed686b4f1d9ea1d5c6c3454390959a732ea579f22787873db8f7823940ad67056f4ea50172f2bf92bdc7e84cab7a65627524c5b6fa2531eadfbd70396b6bb107fbd0e5d92fef1487e5b336645aac639f673be80950025269f48e755c21a91812fe8ecbdd7423f6d642320943e5456f13ef87fa5c057492c72c8b8eaba48a456d741f9077db5e497c147db00cb8695c90a7e4c0d7ccc77d689780704751a3627339f01d1de7e6ca2623cbb1f773dfcba054855398964d23bdf4592f1c3928626a560100ab34f0f1f3e47007dec6a2b86615cc721977616fd6ae1e02be603c7b60c532d1ba6d15fe95effd89038eef1d4759daeb8be195ea749bfd4e40f7dc6c9fdf2c42fc2dddddbdb0ea101f52fb046a510d6d0307e6257fb26cb0091e55de189767e0dd46e4ffb6ab9079fe2a8e8a89790cda0cea987b5369ecd7c9dce6289688855f3f03c36d8c0fcd8114935ae7436bd377f4dd85c354be5fe2e183b7eeaada98f786415f384bee1a25895ab0e153bce0f56b69d903a1d4012e17a4c73e70ef33e082bb8e513f04b9d0a5b562968273817ae6af2839f5dc99a63a24e1bc00b67e7a693d20c44d702f610ae64607feb425ec855556c12b9a4e01e5a2a3532af65dc4eb7f1f9d978331732a9a73ccba8471b2e9d298fb3f2a7e26f6952be84ee205fda947cbb235af88898fe048868c899f1a4057fcb5ec833c72a5f1eebd5f752ee3a25f9c9338eb34b145230a4d99394d7858ea22d06182721cd04568fe2ee756049de777e8fa8e71c94eb8488f9531f35a3a134bcc6465aa760167a331314ad0210e3e30371471420ca2c3e55a5771c862bcbf587897ab30ccd4d3d9c3b52f9fcfa88264b6d1c3b0bd29000b3c5b3a2799798a1b738275c6951278ca202e763f1169552a804f2dab5caacfa1de5bbe50853fe514ec9e14a778427986980fbfba51b7832ff34e36c9964736d50b852aa14fa9c47377f7eef8ef1e3db279607abd4d776085475b079e16ad07ff24aa680df4d3e31b6f3be4955d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h613848afc16208122e535a22bca148e142129e1cc2a1194492bc75982e3d09c5e97c5aefaceb8be56f09efe4fdc6c523f296bc8c2cc324ff694325f54fcdf80a7d707e4b2a2a62c5b1b901591aa3a112edafb08640b92f9a018e2dc53e731f55d956231984c99da35bc442541008723539ae0d212967ab3442cd49249a2fb366c8e7b1819b9118f6501d2f96b7753780919a7ed38db7e4efe79f53954303ae8ce9bf89d6ba11960492dc0ef7ea7c85a8dc48494bcf0a23d3767021d832470aebe7502833e94107625c335fadea874968b5eef9aa909245038479d4c1fc676ec942aa4b49462ba9bd209309d4a0cff20f0370696681e1ca525924f412920696875c9ddfef417016eed1516b6a16f6467df9f5b362f366f267b368f2ca870467db6be6f1e1b7e52e6523033dcee7326fb5b82632bc8f9673863a90b276ecc390e392ca8e0825ec3dda270dd46ed7a0735a0bdaa673da1a57fc7d35f56be9d35a7ae9c8d94e1a4f94cb5eeb017360f583d0e71ed9cd2d721c7fa7927a13f8556ec5851b76a608b8406e80348c394d7081b26bb8af1c4db12d022913a7ce005d9f2f523b83644a1fc41edc0ee7989ff01624498e93756cbfa386f7c0764fa19a4c8354d759a2bd73738b88ce13b9594502d135e27c791eaa2fe394293829dac6da4818720f472eeb6cfa873da87f23f68de0b4f6f484a69f85b098b64fbec04f92fdd369608d14bc2be253aae0ff2802498ae3a99e7f3df8c2a82e7ba0059d7ce5e208296cf6f266f1fce3e9da12ff429cd5ec4a505d0f8e41836545f88792aa025c553ac9cdb2b4c10b9614b7c09f7dae385a67fcd1d33aa36d169f3bea43e9fe83f9a0b89c478ecd2503eb1001d9563bd342a93faf47db477968e4c5052caa6d4cddc07faf559895d94e10b08e6d162fd197426d501f6af2a659a10017eaa33254a8b6f815decca9a337d5a8c1a7465b64b218d62c0f300c7e4e5fdd6e89e84e656b208aa87fbc5183cf8f96ddb13f9e3ea5b2b17b84d36bdf81ce62623375a16b5a816cec6c187bb2aa42730abd76e23d4287474b8bc974b459c8a490e70a523ca66a006897103738fceff602f6c9abcb8134d454096e5dd4914eb304cf4c08b366e472d10377d0718263699bfc66917027fa51733fed8e14ed1ace7d54b2f8227f6536caa84b7ec19b08533101a2c0f503210bd51c0242a57f216331996bdd995bce979355a3b24c14c04ba5869d781f91994725c78aa76960c2428eeca1dcf6518ea14ad6186385a78a65dedc5524d8d9d5f58a61320df5f1b3ff0a33656970732f30227966488f609e2d71d32dc28cba5408e35413756a5c104ca86b7c6859201237a0e4bec7a85bc7871ee1fcd4acaf7a33c50c324b86f06cda8d70866fd927a16d461640f89f2c9cd09e3162d5c7f9167b443eccb6c1b4580a07adc488e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd300451a5d1963acbfd0b159c84495aa6b10a5c6456b1b9b4afd087648e37ab0cbd93fc0fea61d940533a1a16e9b828be75b9b19d891880bcb11a4077efc49a52e1294bb8a6982d83ccf631c4ef79df70952b1c6bceae86737759edf5827ec98e394fcf20a434cc17b6ef1fca9b06a66aa523d5b33bd4e2a21f6b2cd9ca6a78cc2760f73975f2490de6d77dcaa11679664d92d87d881c6534c939e4fa97bb4d3e3e8d0b34a8485ade0215405e84f6700eadd7873f379cc3eaf12d2146d8ebb8f31a8f766d14c1e1bf5a92cbbe01115b8e5cd9ac9b27a4b8f4f02823226b327b7461e2640773fea49cab173bc52111e395db511d9e4afcf8384a7eb1398821db5c6e95370d14b44f74c6c25d1ddee5dd92eedcbf7c35b57fe08ab2f067a3712dab86dc1df4520187190f0b86a08d7eee98c987b1ebbc469fe2158abc1e79c97484ccf64f05d1fd1b5c9fd6b8de2cd598e01afa95446221ded09b2eceab7cdda4fe6f43af7ca3ad434acb2c69e38696e51716f8b61db395ba5e156655cf515edeca04128b18eea4d73415e81f11a67d5c51ffa7581cda8264a88bccae2cb2023210cd5caee4ee2fc7b99c1f3ccc07539e6887db662abf8a8d66b9f8e8dd36a9cacc118938abe7f08d6c9a17333c21771297a4a5d3b6d330387b5638d041c299b91c031154290c1c20fbdece736b33ba62aa3f30a8574951c4b9b1f8b7b36c8f8295d045e3705a511c471bcc20ecf190fea9c99a4a1438f819087d6ed4694644eda577b74dc3b4640cfa04d22c11617983d6bb5203fc1eee3ba7896620e5e622c6ee26e68fd938283a3d020e68333a761aa4f956f36109f3e0f5a5ad73591dcb9ffbb3330e293cb4d71ed9791195d56f58a820e7188fc65123cf1b248f9ec114a85b2078ca93f2567e548a105a67a5d5143e866c1f7de979473bb5e9cf8e357413710c1cb1382ef61f4428f40faaf8f6e36007e7037fe6cef7915aaa2f8e505ee929152c2f7e5c23a6faa3f7139a55acfd9c81b672dae8f30b4a4b4e44a23489faeba38a7dca04c61f06854f6fab953e20bb2ef92078ba17589bf61f8267c36f1de4526f2a84f0bd25dfdef9e8752077c848ae99b26dcce0f266ed74934572232f5b03cac1fa046c0ca2858936ea4f092d7450e52b00b3fab0f5867efdf2cf4252499adabe470a8ea7c2008314b23ebb8e5c8c4a479b707621a18d91e55be95ba1c6f7b361c7bd424de0bc09a1d3268e2a115c89ef712a6ff9608ad77c8d428af68c576f90a411933ce9575a30e11cb8d9c6eb63780c32c560ca5b17a0ca94da2b108d361a5f6d73f69b9b7922eeb9830f370a99f5d2402530dba1bac5476dff7f260a31350951b7d33e32f4415f24d149751919e76d0add0d903300afe819debcc2950fcb21fd391467e2fef6558888fa289482643949b22353dfa4855431acf93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6f01408b9d1b3dbad2e5a7460141d1071a06fa7e4957ed18c587fcf313ae7fad329d95dde443cf3f492ca2ac2062447dd61694cbe4ece50e212bf9ef32b7a690d8a6332c49b9308c930154a2d3b2340b49bb98f2a56ea89b2295a9fd813a115b0fded27c12297b8090b1c80cd31e5966993e7adf30894b9ab6487d39639674ddc20e320e937e447230fe775fe64303f6e284ff53685b38f323c22d2fef1d95f20fecedea5d9217d50c93fd3a8beec3500f576bdb301fe0dba5b07009543a5b104124d198aca4824b4903039c702d1432ae1092ae58ea776034cc6364be3fc24892ba5e9bdfe0dd7d751bb077f8202a87764324407be8fc64c00d586dc904797aa3b41741f3c5b6ea676f07515ce6c77f3648fca57728a7ec795293ee9bfc228b038432ce0978fb1d89a66698c47edc6febafe43440591ebcb56b011c6de90b937e9ad8bb35a29f6d727339ce0ff6bb6d7eab7cb871abf2583d32e00b194db151edb71948f95d37563ebf0bc228817a05d6e5828e59b6e77627a3b51eedde4b480237d6a30bb918d9a0a080b909b371ee8e7e5a4532050db7e0f584d1ca2b677b46680a887a1894abbf788d6416d44c3693464ba6837d0bee68c917f0c9d84913b6b45debd60e1e0bc610089f9076ceea059f95f929525fb8af6d58c30ca8332d6ed265ac953ea66b2dbf7120e41a0635924ead0f00b85c0fb0558c090e3e9a3c6680f5658ef977dc687b871b7b5bb74748a53081752db7f1bd10addef549367d3915ab1058eabf34eb6a9e510e0cfc7fd9bc9ec30620c1ba4979d0c825f5b6c674ccdf4a8306d9ed3a2d1c3d6e64ebf837476a7999143a259622d1e93573ec33c2c55b08ae8497aa7e0a0c33bdc1d3404c336feeaeea6f2b062fcce84e74d4a83bfc5ac65b82384a58b8edd59880c7cc8a1a94f75204984bdccc4d24ccd684c410c16832be9178dc3e4a570cb4bfe12bb93ea976c73caf0112671cb716e345fbbf8cf15bb7da33820760ac5ade0fd56f1ca9befc44ced73c9b77c13aab95109b466e8d04266964536ed6584852c77514f879cf0117fe051e609eae50f565765aa267cc52ce70d8f17cb86cd63f913f45f3224f945f0b6afff53db6e36d7addbb9cf4934a3a7eca7d464fc84706c91b488e449188ac5f9385b23ca497592f2d28ccebdaef7943a5fd2737f82641d7af9a1c7eb61b35cf78cd6d42dae9893ac6a812c2273d07b68f5e19e1cd2c6b2ab3601d70d108835981ea11afca78d80ac04684f8c49c1e7764e7dc6815e76bc55e8bc7fc6a0ea742ceff2c074139f6c8d10244c3a4112e516731a3af8fc7f1794562575dc5515c2b882fdc01fb0c45f819520d68833fb13f23ce3f71ddbf52ef28af7c84d657b94ad44cdc6b04c8a6ab38d7afcfc1d9542c9bd7a17e31c5ec5b054075227b801eee399edbb05b55df3a04a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he815689be7bc45dcdde101327d332012bffd25d31b350462aec40b3b3c32806569a3315c91de0214496454f68aff2e01251657a151eeb919ec8441c0d2593ad6442bd4290a4e409bd8d5c059520d6deed5ba440203335fda3a449791450db1fed91450b0de8843e10657ffd8dcaf5334aaf1ccda7b89708f78ccf0ab2156d58009d1817f5c34a2752e26af8ca28c9c1c7ae928904a61009cd06ba64e63537bbeae00379416b4430ac587ea0118bc41c4e41ad03e84318f35a75cc39d3243f643c4f3adb47c34e2f27b88192cc7e79e65c3a20cf04be6e8952be287aa6e4df27885842cdab5cc64e74094d0dc14dd77e2a1c940b9245c11ddb2ddb57785c6a943381d5f5062009facacf1f073b1d60d7ec5a8e768ea304e2bbda2a1872e54147a1c2888e4510066814e0bbceac4c1a0f72dea7dd62e5d4ca9e72e5223dcd7950a112ceeb5cb4cd74e6531eec70bead405902f80d05b17b58f36606811dae1d64a60242a55f92d7bfe4be1ca6a86338a2ca3efd02f7e621f8cc4dd436217e591f4c0d035738f35d41dd2755a2c4ff48236dd5bc5c6d8e641827c980be7c2919b188338fea2e688e2a30599a423f6fc2b62db8e7e586abdc108cc5ab2fc1904a71809704eab0e848e4498677d64ec21f3ae553a50557610da22b58f4a5d754bbc838d8258552192e1cdd9189eeb28de213370f9717268667c1efd6147e34a7d5490d216f93770eb7d74369cc56e01ae71ebde0a43785893e880004322c1cce59af622dbff5479071ec005e8407b0b7df569da2b9f6240060f00f1732643b3762ab6c6b67a8b2f718caa8abd67846f5633232c371be41a5651905337bbe329f56abc022ff185bbbe59e0b01d05be7cf9e47b19e24a212c128353309a3056e2519dd06a90e1c4c72967c1f6a73944ac3a411a9c1c82378c328f43f6c3993acfeb7c418ece64674548eb88a0b99eaf90851807dc29e7c404119669e0152b385ef6170de43eeda0bfc8a120ccda36e7a0b0399e6212bbf1dcffb3e21a6d17ea70db31a7b74207d6e594599b94a2d9973abfd8b1eff72cb50b8c4924dcea40f05b54e10b4667660508db12f7f257401dca91491403735aaddad0b6410f291933e318e2bc6c03905ae5fe339613fbfd99fbf450a8677dadee8b2d27e10424dcd4f74da2f7f57ab5f950a1e010f41f3e64ecfef99655b61596c13ca4e7b18079dfe7c52b3be603a6922b44b6e70d9bf6fe7746ad8ebce583c8b393605838c5b1a36281891e329df94408b1d7f27d8fa02c882f3277ad422e6d9d49f44945b51c3fef5da60ae04c6d332bca6b4a0529f438c332303d84a949e315086d692f42b710b19d99090eb3dc17c2a847ef8716d3b56e10c0e016bf83efee6b45ba08ba098b3c8497ec49b932a2b35413ea371819efaf24e3220c4dfa6376e9794b0618336c988b53d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h17aa80c5b1c73d55493b694027fcf9dacff62a136b6a26d054b24a206196f0f6aa42b1f8461e9f38c067a41c7673485d2fb92d15a1b468ad6824e67a88594edf07a11d7f496b4ca7007e89b5629863ade0acc674cceda155bd4ff47471fc7703d7c077e09e767b350b68d1d1c004b76627955d1d99e3878e7a894d3881a64c121983bdef790ca3d8f5ac231de3931153b7eaf6e100fba4b2fff6b73aa2516850c50757386ddd8816fc45ecefaf058adeb645bb8128b27145e2aac892926153bf67ddf337213e91ffa03b924c6dd81c9aa7446fda6634a64f4d13167353441e4d7b91c68ceaee7e5542f5a72c86788e7fa5df96c77c0c93ee5f3d6cd8d21e6b3ede81396c21c93dc4f08571c9d8460d0b4fe4cdf09040fd774d3fb913d17da90610e39d54de4c9e959c55a290133e63010db96650cea82bde03a0ad119af16ac0b51e250ee5c72b58521387ef67280924f9588454e10d9e60a755faf1dd288d9639f231f40883bb6c914ed4c86526f23d3e2532ba409c2a48331563e3845eeb378ab06d97453067b65bcad39a196baa7da6b81429d2a267bb6a9696f83ef1dd2494bb31b8fc9534f40861421691977c1151d1df1204cf50c277aa16e3cae6de2b185e5cc0d8a041ce3ebd40fb1c79a26731db3c6e67ea01e13e222e96d98632bdb1e20ecf0626cdd5407e3476bca7db79bc78d4a2d33c3c38d711f0657090d3da839a700a43ef087810abb1290d2be8c881e3b1ac938f60a273a9a73ef0dc5a8bbdb1a72d1e07401b31054405adbeba1126df905976a437543058cd12386705428ccdab3d033d3054659e45b54c9ae2de7cddc1163e14de8abc338898c9b0f0c329a377b72ab19c5e903b165734a49b518075473d0684417f88340d5ffd6bc44ca80c8bbde6bfbe2a95f9dc747ed1efac5a92cb0bfdbd7441fdb4c840b9ab3865f7730958b016da4dd1c91cd7912bc16f26b58029f674e6426e9b14d8eda524fd6cb6dc341c3fac18ff8bf982085a42013a5535a44d9f2069108f777ecd6cf703476ea69b8f2544a5c5590f70b8aec77bacf556f879626bca39edced915bd68432d5e2f320177f5762b2777c15edd154a13fed924e5b1b5d719a106a25d7152ea3e2e6511656cc970574665318cd5272b3d147dfc33980483ff233e5001ac3409e6c2b950aab5c96c85bab0b4f36bc437d74739be680bd74819597a62de28ae088370e819a812aa8f724069e82629ddc450f9cb2a771b2ab5251cf96c8b15ff9e388f6007cb6b605689dad9fea24f1a6e3ef9668a81822034cf1c5443fb5731d5c151f3ce65532e462ecbc208dbfb086919eb56daa9d4bdec2c2e9e3245024d2a3183ee58ced7cbb503a730b1ae4cbb3a7eb8dd5984d5c9d1467ce6148676cfd75ba1b5eec81e64d8283b5e25e71085eeaf9bbd05e447a33b9eb7baa9fc1a563f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h78e1f60139f16181d77d19756d7261e90534b32f77d6509e04f9ad317b999585987940887c8f19a4b3595adb528e76ec59382e3f39b13be132bb7befe6d37bfc6c47a907785a3577825178e0c6bce2403676b8c2327d00f5dbb8cc8ac5d2e9754594d88a1d1adb50b24985100b78f3726699d307b5557e636b3b3be436b6a7db75b956bdc3332bffcfd895e332a7db826faffba7bec376db06a6f031fb25a904cfebd76149be97944f86160a251076afdd418649fdb2ce6be93b920a9851120bd5f44a08a9f3e134a191ccb29f03840a1c89a600f35c8a3ab3a80148272cd0752d512dbc9e9733609017dcdba520f705db4b8d59a90b945fc9b323e48e07ea775e86f502a0887b6a704565b009fda46811571f1ba3624b7e81bcaf2935008b9121c44bfc3d4ec8635e424227c78f41cea0eba868c13992820c53a111878cb3d9f737faf393f0fe28e047c5f3d879e9374be5665f687fb23abe303789292b5dd38be37af8cb88dd26b95ce46e6774fb308a01e725869dc40c7e7bb2c06633f3889f805ff66148f9c6c68aa6232a56cea7a628cac2a6be3a72b4dc45f39144dfcebaf29a47a6f426f0f4e63065e26a02679b53867785f596efa9c958beddb977cb02852cb0c7530bbd2d83d75e7e3c05bbf6cc7f7125b38e5d744fe166685e2a8fbf871701e9ed9fdc74914653382bf84ba0f2d9ee6fc3650b17a7e4e7a6f0d87bd38ff4fd202a756d3014e5fd317bfe689bdafffe116cef6beb4e7a5e42176fa75596f934c0e1bbaea2c81cb250239fed689f1c510c605f1d0af490fd5fff5edf08164b3e7530eb92e86658cc7e0e054476bd99adf16bcc151e9ac7b8d60ff477e9134d18539b2699e897583793739c41e4fa861d741be3757844762428755afd07d27d6791d0b46896848494c326a28ba6756ddba225504f1e15074b0032fc5e702446220261f55eaa5b40ff66627168c750a30909e1a1b5d35200ca1557ee2cc31f8fb25b74f08247e52781a1f6cded25d3a56587528ad3b01340136e4a2597616f068e3f7c5194de2643bbf10e9b16c9bbe177359c537f7ddcec3e59d050aac0ed2c15e3d7310e6141919ae532cadc267920533ea6aa65d78823088d8f89fd9d3f4cd039575ca14d4fab8eeb150d02c4f06bba4477e38eba3e9177d2d31fc8a2267775e5c7fc6ad21a126fc9ce6e1953a0218cf9bfaa2ceb9f817ae1ba74be7f495e873f8e1979dca06f88a7f013979411b24795b9f90c7a669304a35e0c16bef515a7679ef1786d4cab0344c9ca1b7a9a1ba5e930a3292d6d39a8b1b959a9d9c7c25c56d6de7198ca1d5466c3115ff0dcb0a3ea418dbf62a58f13b39aaa33c615f9e54b1e86bd08ed317431d70ba55761c249114780723789974bb3d4bb6a21e9fbbf5776c6632183a81893e4c7c3dab8736a12750a6e4e2b43c63fd6f0e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb025b43ad684d18b082aa0777c42d1092a396a69d9cd5d69d7cc660f74548dcc60f9ab07c35b8a3d32e2467730b02312d6145359be564400af4768b492ec632e69d2fad8353bc9f355185a1a92cd80ad61b3ee38b2e5702d70d520b2e00d244253f9cd634311ee3224e8bb62f68ce8e92882441b15aec8787dddc9a34ebd4aadb13063dd58070432e05e53d77985a70f0b6cb1f18334fb0cf00136147e265af09df1efe42bd92bbcb314c6970eb690319bd8d6ea7531e3b1a139fe2fe4ebcc8e299bfd91fb89060cc4e26d5a030c42b27db59487100ef1a3982fa7833bd29481140f28218eae07c279fb88a2e9a878923dddb28746ca91fa74cd0e269b6a84d8dc78bbd9ba275f6075b0a1cb511916b7a1a9e07c4058cbc12a3b0b708525762cab641ccababaa13fd8e4a7aedde1f7681c682b4394dc57eda956c67e831932c382dfbf00e2375db519bad06b6554f7640ce92f188b59c9dd31c7131fc475fffe15eb25f2d6970175957ba3feb08cd7a413bd04f02d7bce51d55dc33593dbf52f77b311c734f2880b6cc7eff2587eaa69941433001b46df84def0360896a79920d4c2673f4501d47db9c6d6ea2e4fa52755eb11d800afb04c28d4f2ced3c0f1c7539809feb766c7ed5621cef758bb8a70b3d63ca7eb637bfc9fe1996dc546f8c8fb1ce89214775272b45111473a15014f320da61f8b4d9b046c8d8f2e3e104fcbe686095e8ea598eef9db175dbf18f10df53c591fd0f1fd8dfd965f42aff43d7c1ed81ce7abd5a7096ff60f48e27ad3e594ebec172ddbb0476ef9d2c6365919bff3fb86369e3d4648b2522c634c92c6ebf80e848147daf7a1c06e1aa57bb9d1d4c232cb433ef09e507bd94db61b2e99ddc9417dff90078713ca3d0361221bb4ea593c4efb16c098ba70c3f29fc7e8107e0c24cbf8102705466fc1ec08e3c4cf75a16c3ef23929ccdb205481a8120a21e9ed9ef49f74077fdd3ebc1bd5960d4e0d8a3e4512d71e7d9f2c102478493d8d38f8fcec020fdcd69acc66e7482b2a22b509baff9934b91ec241512ef8f6d159003fcf8a31836726aabb77fbe1cccbaaa668e570c8bcaa32b774ca723d3a8a70a53300770876de21e7d2b1abe7060257c3a3ccad9bfe22d770f03d1dd21c813cbaff06845b4c5527f29cf2b7f8176b47f1bd37f9e948de2ffbb22c194176b071facc8dc9cec505b1c3f7fac865efe8299cdcf9da8c2b87efe5de9f1b20527e428d8be21f61df398fe57d5231dbaf0562e186de8c35b08348ca0f6fa654735f45c3e087c60777ae123997c07880a095bd917a884754c0a35feb60a9255b46b7281e17681303ce4d32ba1e5223e36174c0fb63488e5c5396de731acdd7297cfd601b2663b92bf52866bd5d2744f5c4f0403282ae5165b0aaf78d4b0d20a973003244474d16767e7769beef4a48a2cbd39ad7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h637ce7eebeb1b0f0a4efc06cbbf793205b924b12a1cacf129607c6d4920ba9b2cfedb3ec4e3cfb0c2a4e533c5f81f2740750a860d0109c9ff6ffb88bf479baaf91857f73c46712d0516f7dfc6ea01af1cb5e6bd9e3f0e2a7303fb2e194716bd2b1c159a8d67998e5a4b918679ee16b12b03af58aab176620ce900c8556e9dc737e27fb4555e07c6b633f13a75d244f236911b5ddd517ae37c118ff7a7959274911444e9c7b7dff8f3c54fed313e24fe9e1867cf508ac5f96b4bfa5a25e889582404b24c7ef839834b44ec6e02c6aa503e33469be3a90d4bb33ae787dfe3727c9299328d84c4059ee55d3e2b54ee695574eeaed996ac0e4073bd5ea2e94e5f9ccd65952740cac5efb4f27f3081865998db96dce60773c3526a7c3e229057cc0bf958fdce750109b26208f4d2c591c88ff3b06f6ffab0e02fd63909131e3577bc404c8c404fdaff9f88514e21b1f9afc212389377c92dcf073e0f2ecbc80732a9ac6ab29723f50c97026213c0981086267507cd9972dc06520629716c7f83dbe7605092e7355850bf5d804ad32cb942d839ab094b7fb0ab229db503846d18c1fe878584c3fcdc9b45312a3a2af553a468af44981d68b8000503f47b3a27b78ba86c633b9458b5b328f263b7b23d2682f37ec4300799e4fa81446a7118f0226039aaea10d2e79d3a3dd8f6750ead99f5ffe903181a0ca5e1e901e9c136ecbe1558ebdbd6b14dfcb81b2c8caf98981db4bd7389330732fa7d2e492cabd890cd5f39ceb6ed10796d63c2a374102250f389e28decb5deabfc7771764ee4094af9855b47a1c6969676c5d58b17cfafb2c300a406b42c0a1f378f1f4f20670c9ab802c57c3afa6c436cae41503c93e9556d594c9e9eb07fed20dd7d677bd4c513e6ba1f0707744ba6cfbec13a4f03d7141931291a20a9ae69a3335ed2213e8e12d8bb3dbaa3549d4edd0b903f3e2cc3be7a1cfe74f8af033d5fa92d3d88dc412c654ed12372c1bd944f37b09d09c31a6f5d98c00473496dd112291cd8d6f577e1f99be35b63b1346173567d72abd231809548e889215e0aa46ff897cd29a28a84db1061a196f9e4c618a48d9ab4c5837666cf608e2f4e2e5609dd9edc662a1d2ff48127d239351e3162ec6ab11f113511a1d3636b484c4351e488e8c99d1a7f7510bb5203014d2b74c139b882af98a273e6399cdd349f6571b5477c4e07f34622e37a41654158ac9eaca75382cfa2a54e90db405d3b8f62464ebf7c16ad1b13260cc6bd9ea619d27ae5bf09ec1562bd7bd64ecb50f10c400f21abb88e7a6243f44d0f2c3de079467cb2b99e0f1aca0b72bbc117ce2019b41fa792c4c46cb1c372a2ac1e7649ff103a8f9432b0bb04c3a088fa48b8d43e062719fa148fbfe0272f9352322fa04e9bcd319dd27f9c4893c7aba11c2bbab0fc805e99148b1f67336cb109110;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he96dcd9a00abaec6327c74187e4321dda08f8b64d3df61c3a421dc31d9b891a2dfed3730a10cfe7d146f3ff6ca4a41cf1f62e01d954b43aec0c8266f6744b32fa6387982af05399633d6e76fe69883afb7368be3aea41257f68ce29c886f2c107aa97421b480528ebd9c5199a678bec2a8b41615b5b182a83816df825940b49de00de7189ed32a43167e54180269c32d27199a52a963504b665775849a64bbad07d46d5823b187674338a8fed9800aae7ee208856313a9320b1a3d58d8cb3b58dfde96b9890df97a19465b2de999620256699c11d144f91a57171f3cdd66f326f55913b4c8ac70de1bc10091751ca0c183bfa048216ca735137b58685a748972b3f7fdcc162f26df47053ed5ab7eed4b4db574e203b33cc07c6c9afb6f508e944a2496160da2cec579ab7f1e60363fbc22d62ae18246be5b36dfe3ef5ec4a87ec12089440a28bc667ad05d28e925702a508c70fc490fee6fe5e2c8876670cfccd7c697dc86b88034e25a29812dc3e4995fe815bd5a178cdb73c8873192937ceffdd74fcf5b385ef8b9f16a86c7210d61f57a4b7e8e1f1ebe32b62b384217ea6319a5e93fb21ec31ee27e0aaccde3d48a98c5f8fbf08c122b67619011505375d21d958a96ab16dd45e6f4b132a8daf420215c92e6d1595a39537c18435aa64351cbe5b749c45e3130e4be582f6066a6917d6f5b6917ad4925a83374618e9a758626b17f163c38ac2db27092c6661cda8789a2ce692ae76f629043a000452c0214a3b47a5d39bea8170eaa147ec40805be5952ba5c32031a6b1387c29e813c6c7ec6c4ecf4515b7c61aac9ff9559d2b06fe533dcb22cfb2174cc4b4541376b9e6c588d8987650e7c85014970f6a6829f44eb951fd02c0f5e32efcbfd9567e1d198d0af7d20f48c8bf1a20636294c2eda9eef7b7361c2b61edb75a9bdcb3dab1fac6df8cc0ced5a3358e27f56402bb94998614c7b1bf0f8ecdec15e915edf9c39eb2244a3f1422c72702a188c83c485668e7815cfc84c18fd30abd33b0bfbefba85ea5c7435bdc83d31024f5ebb7bdd97011aa8e9181c84b953872c3328bd3bdcee9db2c9f25476379f6d8ffad8a77d23f19e5b07c127ddb3093b7da24920cc0e52bfa74fa4bc323637ba395a9ba33eb7669b7d7f96423f93913ed21d831a186563f48f1e2c97ac5b4f49b9ff2f79ea9d5557131776607bd026f7378edae2651cf3821e61816f75cdebdfb495507583c04dae7c2e42fea9cb71433ccf5b70ccef8f9fde504c1e77ef74f91701faa93b5ee24a266f9563de54c18b9f4ecc0fae80fabe12e62225f944008b39913f288ac4a90ab2969473b4511098db6d2d903a4e9b6195d47af79e748381577d12b75dfbab8322ce2b0e4d0e22c0d9c1fcd8b3703af8995118789d3adae1bdead6acdf6f2e35af7908fa8cfac2922927167b5996fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe9075b80806e923361407bfd9d12e386fd01a5204467e9e19a294944ab6f19b43b7c3526c56383279e474d08de93b8e0f4225ed40971a62da3fb76347d2708150b698e3f15277a915510639a7a6a19e1fd100fdac7462a996af7040113a28165688002aa99ee94d79faf113b1f9c175982ebc6400ae47059a73489e827b320375d8c4dc54d4e53a5b00cf109f60f6300ce52ad400a949f2a0e9d6972c3c20e6712aa38e89325520977a78e31abdff00a61aaa63f2193cc6bbe87a9574629eb0173c774d61e11dd3c8cf450e8c66a486f8f322759e0e0c663efcbdb59e470edde25c14ee91df988e4dd7e65c4e2ee8a9f2c12bad4b1ecb9c273866a738f4580c9c716bf02196c8a86a4519352e852dc73ed63128d10ff0784c00c2d93b1b5eea54282953a24664ccbfec0f559fe84034ab5e6bab9b06cd13af1aeaa17ce8a2e25fc633df19b2df233862dd9ec2f70962ae663220d3a8a7fdbc5674d5770e74b4b208ddc32e117b111db7afa71b291c54205c383a8acef80b48738d34ce2de00c8ba30e040d72137a1d448eee1c60ed86a26bb602595817c58ce34693a44b026f43958ca9d75b8333057253f4d3f9256bf61bb472c31357d00c2c36340b9fe00f496a08e6aa29b216a37d8658c02f487159e18c58e2ab1e31c65ef1bbbbbdc76b2f982796bf198679e0312d1a3a8eb31c26f5a5bae113426627f57ecb0b65e1f3eb725211c9dcd610548bdd902e5ff5de08874c658f945d8a6d037ad7ce67ba86a86469141fe19700d3f702104313a41f7d7f78e02c016cd10cdc23b1e3aeb46dcaa747a48e7510c0844788257d645f58e318d610d67fccb108496dc6ec7e5799beb516badb42e2922b95489c249525e87d72289d7e16a9e788c0c671e21bce7145e267f27fda4e29f5e70ee2b572835c6afa22c5a16498315f5b47b09517de6e4ce79810220674ed0143bebfadb855b37be9201cbfaab26494280e1916b64c0fd4aa72824cc06d34903f117d11a78c56e9e422db5583e1215247b9dcc854ed268b344f28590546f78b30fc14e73ef7d0f048259919ac6e6fc07ad913a0a600cf24f5defe0b5c285ca47c8c75f9112073e9fe804f04c98de120bef61a1a17018ccd0ab3b67fb455f70f39c9831c00effc8925f8cc18886608522c6b4d4212e349858fb0b22864aada62eb4b8b1de3cfbb9e8786236882e4c47ce7495195f6d1c9a26f8c6c1751b43db93d643fc9204b85aea6e55250a1bb674ac65fc2d5de25ae995b5b5f5740d42e5ea0249eb34ba48397bc5a696adcd1eed5ca624e2f44c4fe367f37978e38dbf91a16a4abd5cfbd727e40cab04484f83d8d0f956f3cb400c3c95048935b093d2380263aacd0032f2979c8c3f98084005c410ddaa0d72adedbe12a3a53569161cf0849780a0b98240a4d8cc3084fae55a099901b7ec25de5c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb40e952a125cbddf922563e745a7d01173ffef308c2070a2bdaafe19c9e5c0bc2e07001a512add20b96069e8684b0cc6ad68f814a5a3c24910c74f5cc7fb99c73c48d5dee967b56872a054519a5df939dfc630c3e45656976fa598a27ba292e42cbfaf87fb10a4b62ecae22cec7966e4355c0655683a5f7a9dfd3f24e3ae6537015b8cecd0e2b0c2c5176628f4e5ff85298b681633331a88e74f715f6c86ec932a9f822ecdc8b1f19e38209f3ff1810d5eb36320bf7c9637ce9aba46d6dc9a9b3e5d398d026f3373f50d65bda06f88588bd9266fa889b3ecf9a2ab1525c502a67864480d121614cfc2caef311fc0d83b1531928bcbd28e764d6dd95e311b97851439ba47f7f8d7a4b3bfa7e71d608ba9bb18868ca4669b0581f22181596c482a63bdbf7a6b38a8d93aeb796355c58ce8b42ed0bb80edb3facde0088f4a99a3d5ef1c87e7ed356571d7caeaf6cd305ce5022ae8974d1bcd0a1c51d503e7fe30866bd9a07b5f83f2ce558fbe67d5152f471de69c0575bbd88882dc75efb30387efed5f4234c6a41e05021164e08d7007fc69ba645b98451ff7c28b84dea599a05b36a72a20e41f793ad2d004a07805324666c3d665184c37846b0aa3d83f1459a883f8557fd3f219bbb5d4bf0875bf902f9d14fbc8ae55fc6198464e5259a70f3b77508bcf5093c310b2725b5bbb7ec5225437faf209d3fe3db3f696f02130612cf45667effe70eebdfe711b85f036e88b76e1df9c3ff4a0a71dbcc783eb52b4c190a8f9cde1c69614be244f68eb5949ab29a6832ed04f7d56d7740bde3e85df7b28382c2f3e65e88cd83913e1930a3452aef945403aa74934b8d82eb7fa69d34c696ff439eec786dc8c14820f9b653934a7ef320cee1ce294217c59ca689992834db1827d0154e8660b54635c7a0e9840e0098c4b319535b92735b40bdf7a77aa3245a2eecdd1ef88c8ae35d35c14a5c43f150c37ad62e72f140ffbdfab3df2ca57effb5d98e804488ff02428169ed281699d3407fb3f13dd652738ae75152c98f1a362e35a070c36c6c9a80a88f64a961c91274fe088731effaf4990144c9d2dced3434bd15ab9e25b77e57d5278ab8087b955c2cb633b78cf6b8777753195abe94cad8f4ac9a0ca85f111ef208cca00a9b1e59812782a71dd3fc8f0abf3f824724290a2d539d9b63d5b17ea7c30e6fcf0a482e614d9723c275de6ff2899077d09599ded213a3872b8c5b799a1abc3d8e63d12ded63b47c1f593bb537a379709aa5c8fd8df3a48802eed6f131e1b7abafe7c4d895480bd6126b779fe6457e44f445cb34a9effe889a7303743af1786360c588e3d2804dfd8483c62f3f35644e6ea9d30b28d6356cd2e2e0c7f028c637fe2a53094e314de1d2c23849e8badd191efc44dc812a3797edd71435b36bc44a9911858f4159453a3332f3cbd654eda21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h61cc0f6425c3004f1a5c7099ac350b7fb853449b3c05e0f687c32515b66543c6114170554b5d4fd59b7e7514020acd2b47714087b6c10e7b821eb7463b52987707ca24808c6aaac9aca130de44438b39692599fed656388904003046b0526cc8dd6bb0f9250bd87867276d6d5ed46a0757b33069dd22ed4d571882d0919b769496ede66ba547cf40a393d6b7a21b7bf1661513ce8a8d3ae4569ba07ac5d1b73ceb898f17594d688cbfc0d0d0b31be6ba225fb6884036aaa2270150d11748af6998b01d54c2c0e4ac1843ebb39f028e1ff4af024cde192d57f6fbfb8c8fa13d691a704185ccbcc2a2133172cabf4479272a105156083d03969c0218592873afab822ee80731d4cc7b9877b88e6180f48391c9726c1cc10a65be343d19bcf95b7fbad629749dd8727db32244be14791cf1ab3ca4c312b768979ba1b91a3e4d2181283fbd9297195ffd464bbff8c5d5c275ad1972eeb507bcffe06f8f80dd9cb7f1b48c8a81b6f88b2e0af493b938e528134b010bca61cd7f31bfbb9df9f710f46e555b939179fce87e86d304df8b0b5010a2b1e54702b123833ccd9cbc4f44c569682b65b0fc9f800430f67767878bd7816e538cb6ed7100d37e37d9c0d29ef26759358bc627059640dda6c59ac0595aeed130f0808c5bdf0a3b73ea795033b38e963991f0adf63cc0ac5e5a16dd8dc1dd71ae9c3cb131b456594c0d53b9210e54c88ca11f31b2d2bae1178172e8cc3ba74f43b6dbea67b3dd6b2eb665455dd0340b91b980c3774cd6130830e1149331a89ee62186a3291bbf23011dd4d082b42fe5cb12d624bd332740a3d6ab5736cec91bb3da13453bd262821d3dcef2c66e1f24dffffa001b850cfd59f20d62b5271825a7b499283de14002d8af130be3e6cb96eae89f4770c8a6f2c45cf77b7d9de08d4312baa13f78d7291f29fdc6f0e0a2f7a19b619b8d0e3e34dd2a5ca19caab4faab9336b70f4c7c88c52d03b42cf4b5c342298b95a961bf893123f9340a0dad3b6da386e95d16226f370a90365104824111c5d781d248c8b06cab0543558305db4fe993a9af661ef6d94decefd4885b27f9018defcd8162711243bae3be9845375717393b565bfac4deb064fa11b183807d36030fe0137d166d49c95494548e38b95730dad155ab643ef160cc9fb5a71c91aa57d2afc9612e248324dd22e612da73a8d7c42ee10b58fd50e9a9353e78fff0027a37d92429e67a681d5faf9acd38ac8a1f17d7e53a30a54253fe24f4c85dc6024d09bf9e8d7fe751f941c538f3267fec7e3d1f6053aeb4aec50e0a7d3926e17ffa7f4f90bcc99095e4d107f4d89994913f0bf9453e89d6ae3cd9d1000503a95256fc417e10faf53c2c3602c1837c9f10ebb93b832e1c05cded41399802fa032e93ac6f8031d507683306d155d6179f9319002fa54d6d5e0ff2562eb925;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h104a6a174573dec97efad14b3ed9385b202963fcffb789626a5b62bf95d8a7f5e2d769f9e14902c6e98035155861111f0d9e169dacf265b477e77675d111aa5818958a8a84f26e0d8cf38cb186d7f93f7ff2da2c345beb1fe1739f0f983723058a6d14a37d1fb474a2b836bcffb38b2e3d3b13840ff49f9320158f80dc83d0ca208fd228578a6ed73cb2e195c174146b336b598482bb45ef46b59c7fb06026d0721a724ee794a590a6c8822ac1437369962273083056671c479a26224b46cc82f2803d5b3e4393d258ba90390159e3c5da07586281483fe1c685544cc6163dbf240d3f958be94dab878f9a3a9c879e60d313b34ab7d5fadcefe518f52280719464b8871aeebaf159c885a1514cf81b72b20e16ad8464ee37eb7c860db4c74376edb34226e715dd18123620f895ec0dd4458a2eb1a1b6a2c3a57f87089c4aba58b8a52ebf2c820659ade0a7f9c562b9f986442c9bbcce935b5d422786d392870a716692f8707bcdc4491325269943855054a14393fa4e421bca682a6e7b0fbb9c21851b2720da561c7d74447887227b131faa1e69ed90879d076bc597bb35072e5f570c64b1997aeecb624c0804b9740a38b2c8eec81d26efd12c3e65d5f5810c4a435886eb893e31446e3c5af96323ded7269e2eef18de5d7da2317f35d722256dd36f9f2bfc2f3ca3b9e11637c79f6ec55c0e7d2a4cb6eebb3f5ae7f4f9b9a6a268700817c0e111ac5a5486a21279c5036732290c979d81646219e3ef116b59d48e12bb335c3f86d691bf277ae838b57cf9acefead38617b7afb9d768fbf11ac7674e901dc963f0337a7ffcd8457f19ec34ce2cc00073f692c52be21a82c5962b6dc4920e3994bece9dea9bc1001f4fd6f3f84f1bcde292d251608b6b3f06406a11ff91da932811e52189bb1ead57b5cf6754eb7240747cb21e288d66b71e9bfb49969d20c9a6e973b475e7358ac22e7aff1c63ae9e220f77afe4b46cc6f3469e104e39aad0071822b4e725a2d7f41c16f31fee9d0dbfdbcbc4dc25b60d832bb35bcfb870f9354eafd50399245afa9d11f9bc34feb648947b241f2337f6cf6751e45f56c3e9b6bdb0505a3e99c7a67858d1eb165c82d2ee9111ca16271a7ebaa7d9e82e2a8fec5463990f99aea0180e2c2419df56a6ba0918260ae93dde7fe0a995de472fb9f9d011acbb96a936719948e8dc55c47fa400191cf5502cec860a4d06219380c07acfe48cbd9bac1fe0af12525a47c35443972d239152a140b9cf607cbd219f867fe2137d2f07c89180269856eeaf26aa41765b9e7a46bb361ff212b0d79aa2ce0caf4ede171b2e45a1d318f612f207d66888d610f53c475f97fa575d039fabfb42e45ea42917baf4bfd6985624a41f663d5a02bcdcbbaae4b5826e274cdb3028ce934266a7d403f5a367515bc0b2ed76bd3e61c7fd486dd54c33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7d57f25ce42a6fb4330da602ef88e824f52822f40996e2322eded062ccafa5ca8da6d4e32dc981395275b522822f2bd01093b2ca99eab098c7e2c19b305eb3b57c1d433678639eb7e4bf0c90aaba2e2a2660c3f5f6fdbfcf5f40c9945f6219e3aa9315b6ff0771810c0513b1785e8e323d9d36815a86d7eeb07415f811efd1b41b9cd31a75b73969aaf8d3e40c60df7b31bcf327ff0e5357ae3d8301e421cb8ac6b959f1860c10aebb74a41cc3a3275c693b7d3988989bd9679ecd28a608b70b3a292843dff15a3508a86a42dc65a52cc08df3215b72d944bd6c5e1e01ba3ab04b2d931fa5eb6a826ef599eaa0b3c2d4acedf779e2c59355e4e9aaf9a137599c3fb951d1063ac17b04eceea7b0df80c64a72015e885fead62dffa4ecf49ccba9190ac904344feb66d490b57dbc716178f1930064df07a0c4bde0ab5fc6accf47ab1f3b15d63b0671b49c1ea4e7283e8f138109442c31a54528c28e53916e263bcdeca5bb2d434f20af3e260dff79e12630ba9a5308a5262157caa5f6d51822421c314a478cfd0a1e4d928db64ee160ef747002b5e7213c3d6c90ac37d9c16cc061e1b2da5892770fa31b5536f03144b1c63db5ad057babd90c95a76b949ef9eec67f7c75b63efe9ef44ec223300daf1f9e956661e4853b61c60e2a8f7d0370e226ad7c0331a2ff53c81a35f3598502c0363cd3cf96694a0b424fea6433dec996f94e9820aa8723d435499232830ce5ed3fedcc2284d955b829d89d932f765e876292944f13049e9e34a1b72c423bc78da35f57d3a518f6b60a7928077292b44f6b707fd5aecb5c22c7d71a09f12745a87a195edaad76381b16339ea93ca2a652a76b54a5f30dd12e72836df148aef9f0fd9ed00db10546d82db8ff9048c80d0e22aeab56e68d7c8efbe817aa6f6113a42fdc907c40e2508c79a1c98b3f500c98534e124b22446d109cb0dddea95f839a434ddab78b826dd947ca28a0f25adf042402a9a0a5772c1725ddf25dbabe2de920b79296038d149dab4a2f72196e905970cd70eacc15a1e974bcaa7b1e92e5a81398d74350eea21b5cc3c5b5e33e0b0d156e9a2ed9e2e7b82de1a482f7aa0c9b66df89483875b36c88b234722718737bef38b4b73b3f8de279e1267440f343dd5d9ba9f5e281e9514dd1c04a6e1f20d0deda815796ed3d9e786c6fa5db6ee4114d58b8c4d0012e66bbae060c79f48cf51efb5414ebb2efc4e549781b64cae46b35708a5f985aaec9233dbf1227b65a9dd87ad37bb3d5c3282a5744ce1bea50bd7f836f3cb4d0cb95541e1b6ad9c2bc4e5337c76638694daacc406b8213a21bca41aff2936ab61d72655131bd1314b8276cf1bd8d80174db9635fff3a1dbd9e2503eff406dd32e13df9b7e6ca3d360d122119e7827c89f99416ea0627b6fa19a071d05533f1f51ab39dd1eb67f43c73b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7672ae49902e5eb18c7bbaae1704fc0667511083dcd2a881e1516257358554ca1f8690d992e9f2095aaa9b088779541e357ce06913d733216b1f4f795fe64474c3210ce3f618e667e834c653fa1d7cdd62e0f54656808e1c983c961d378f4044f4362db2006fd1af56090401af076a5156bddc803385ae04db7ae91002c50eee8bae5ebbb4f239e4e8e699153330f636be5a6682015532ec849e3229186c4bc9608730ac4f8c3e98e927a0bc3de19bb7e0d24fcf98b8ed5b30ce2645aac41027e879c5d146df9afcbc8bbf818347e0229b39afd93fb6c56fb398be7b8bff46efd991feebe391aa446b03ed3dcbcec3122456f35d6bf06e7f457d274d807db0758805b78fc458641afda75c9322aec8e8aff129ed9c71c25a42409edb94b38da8e2ec5a36ced1b3232b2f92e8ce53f7152ce4174ee6e92a056f4bd157c36f91b737e8e707e110074d89b2a4a36a544c1342e1931e6a5dc695d376554d60f1edd517e2418185d2fd6ccef589410c253c01b67350e4c731632bee0fc0a677ca34a5d52de507e27eaa1ef1f7c77d45e52b29235653d977d23c8d213e9fe3e2cf557840523f02f10dbb25eb4cf942d6ef5a1e63f7ac65986163e158928a2202ec08edccf1bcd78bc039711cf3d2de9cf5432275c395d2c779071ba7c466b04a39cb6a34cc119fa09b1d877d6b293173801cf3a4bf5b6cf6c601e3db79be34b0f8cbf15561173d5e7afddc436ee5246e10501c31b30bf22de4631680ebbaed6f8aa298e64259e199c7e08f5ea6659f8bbc77415595d427c714c7ea29d1f2d340121067990da282684a27d279b170c21f3dc5f407eedbfb0ab2e4d4ff6bd3ae1a60223caf9bacc8a66727e77e3aab87c77ff867f3d90d044f614d26352cdd97217734207c80716e96dd1e7b4a08ef102447c2c968b9b000689e2ca10e7128b91b993c98539933059c2a79c4ac4f1bb19f5b2c834087e7a85d49ad173ec14cf9a0d3580fdc20f8fbb214044fc620152935049529c42ecd75cb5a171820422c3afa287f5979140fc3780eff6c734274384954d496e15e32022e0d758648e79b712022e2d19b2675efa9379dabecfc2856996ee75276b3db19b30f867afdbc5848ff6be55538d1ca643f5430d06be3ba1d25b9149cda4111e760c806882a4fb148524cfa891959ddac5a3d0d63a1499ed80bbc59c12644f94848192cc88caa997e7527d30b2c2a1681fb475945df4d834c9c037fba3ced6cc7815be3f3c3b90f4adfd86b8ef53a8415ed10796bfc6a755372dbc85e876482bd75b562a5b5fa74324af18d4272e830a680844028524294410156a16027e7ed8176c753bb5aff1483bd7d5501ac0d842b0eae4fd382022418b9a7a475351f64b257540fc7c6d8ae6cc18f62e4819c355a4d222ef37180f4bf62e6ee544525090964bca5a24763f2cdb8078ac6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8cbe4330ca2fe68978f615238b61abb44c4bb8860b12d7bcd857f95d6ce1150f3d0575e56c65761d84d68c13def928e809099d73d6c57a1cec4c29204d6badd99df6981d82d1a27893dfd7d06757fa3cb36b5e50ba6b94fd37a5e9316984ca1e8b3163d64ac62b76fd539645aeaec72dd1a0fd3a7988dbc85d10fa99ad12af7c37f987b69e1e4f4cf645ad3ac46afc6b0c9886ed0d46674d3d38a98fb2f84f238d4f239b2ddbda6431543c179e32066e49153d04e8bc7003b83fe64003ba2173451f895c171bd52a368ba2c2b15abb54a5e487f4ff7d32d09b89af63b6c3f10126d5156c3f87fd40ce837f609e9ea20e0df77b7a4fdb5c50f882c7d6d967deb359a1fe986713ab17ffbb63b377538274547a017c61f0e0bb92115c2a3686340e64a41463ccf4cd224312f9f775e8742334420259f7bf09d33e89806b6d0ab09b75c30b8a0120fdf065c92c4d332921fb65e99307c7c62bd5784f672da2acbafd7b989eaa025aefd885723e43325a43e902c44b3c268604cdae539ae34fcc483f22f3dffe1da4b67c3e29e5f08b0351ffa1b2d63c10e0f9e3d79b0e8e3fb46b7a30fbd5e7b9f83205560660b2de74e577af22c3d9dacb473addbc02370fd01fbc8950f534cdcfeb5b2eaefdb5a2c9ff427983dd5e4483a26d12d65a2f8529a575f01a28a3ebb93b908a7d17788a7ad16cc01706f8fe1bcb5183a162fcbebaa51afa4193bf756fab3f3a8e335e733137e488926e565d66056dd97950245af0a3ad61ee59db54784a61892e7775afeee8e0960cb21716ab9c3b36de489aa0f4b39624707e19abe45966363c7bf95fcafff79afdaaf5db174dab5426739fe6491bcc8e18dd961692df3065872a3f04f5a9a7ba1c8a82b1fca6b308be7ab006130985c3ca6639d65cac024d7c154ebfd458dd617d9856f6e21a5348b0e4db33f1d38e9fd3432a9a39a06457d073dfeb8f0e488a74986f90639d22758047613fd40d9d3bd6debec1aca5e762ed4039f9a4862d3ac62f008c2a577407c3288b610fdcefb6c5b3de8a3dfc9eaedda82ca1f496aeca83e518988269277d65959213f8f2ee39262dd26b715189c15225d17b4ca6f58e5d548f9b52c20b41a684081e45391ffd2975107a9956ea81f43c42411b75d78d250b827eb6793712fe97a95ae5929360ef4b940ec6180d3542f4e11f9a86fbe9ae8912f83dd22e727298a2c079c4575f11bef2681df2d36c21aefd0e3a2e217273acb8d1b5399a2d3fa25a6eaab1db43409dd99a6e8b454a64e38ec1c084ec8c0c34a6c1b4901eeb2bb89ada67458c5d8bf182687c41d9b41d279b424ffb171076f0d691b5561a1d101f8f54ab4a0f4c6d020c51a6844af0d028deebf4761577297fbd2790e0334c0c9f130eb788dd1fed2a2cc252ff5b30f1bca69034fed08ab4dc91f8a33c5dbfb24896915595e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h34948479807707969d8ccc79563599e3fb499cb54dbe72f3d70620fbc0185ba40c1cf68f3c6765c6b05056bd6a48cd43bd0ee05a3358f5a5d2cbd62b9d7d44c5591dba4ddf594c31d1381ef0d4af5f8607ef40e55dce176450a9a7f3076b68f83bca8faaa3b871c8ea08c89bc4c672b802f817c8989c293ad59ec366999542467d8a93e202d27c4b5c05512d9c94207d375779345a5a86765a6874aa6b281ace503bd614e6f3cdd08e0887e1e0e1fd82e2b8b022015111da7350fe215b497067949f91b60953699a8ad8260b6ae75330a367f5ae23c6c2c7dc0332bf0c663300ee727d072c12ce1922bc940b202406929feed4c170c528d87b5cb13cd0cde77cf74d945376020115d73524db349f874bf548bf76cfc04a7d247888ab60ac7fcf73084fe72f4ce5edd87d6d7799d0d0524e4607e0d226cc29427a2e6d81b415a2fd8e0e416c8b18848df4399543377dd1845cdfacfaa593ec8cca3f2f04431dab72155c10639e1254a699bd2627106503a7ac7b96d488c1b3b60b370bfa666231f53e978641ba06e334226ae7af8d9710c434bd55ab72e8b6acb69739f5557a2f336d4b0f8e85d79becbc168e2bd7a58578874722327ead80fd24a96eed730a1aab6a623ee9c6e192021bb8c75bad24a26319bc66ec84695a9d7575658c5e11a2588ac6d9443c23d6777c3164c7fd2f9d088e7659d2feee125fe5fd61747c977fc0907ddbca6618f13c5359eb555ba250b5c5f96c539683779118e8d83b5f2e5fedea47c029d936b88a1c6215048fc23c3b54bcd90fd0ab5a562575961fc096b1bb6c528a6fdd58cdf0413c8deea52dfbbf4832c5884675b8c109348e0aabcefec096679d23cb6ba269e7142e87cc06141525895108b3a83441a1f5111dae406219890c21351c559eab832663d10cc46f7371f8fedb9f9f28eb54ac6aa90b83362ea2d7a9f523f622729ff511575372d170c6575cf972c79e8fd925e2c47223d1da81a5a534ff211426ecc043d5a62069f5fd6c575113a5183d12d979635741f932f4c50e77d5a625b6597c5477339b887fa5e699919388fa527a17753ba7a4ef75b3004fb5488e0c5e6bec340b73bf7a42846572683b23d8710a81e127366b7d44e6d613ca27d0a731c3ff60c649a04797941f479285fb3553d13054157b59aebce989191442c4ef9a6d4b427d0d8795cc5898b2ec8782b737235420d0d4201ce51cc3bd7b415423f0ba789f501ad48f348464808a7a1af4e2c5ba0f3a5afbf14c864ded8de1e4d5c6dc2d7c3b07ac6895429811c4bdcb9ede0f24d85983f9877b0fed2ed331b63983bc72d5511ebea4fd18d730be47c0cac98a17acd7e328711e3d5d0993c037e9a07d172db6b88b0d802072530082ddf0200edadc6f203f77f633cfed8587d37416d85f9210ec5dddec02ba8d07b42680f36b732b96d6ec3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2167ceb7dbb5d18fa9861dc7309da3637ea80cea796aadb2fba82582bbd602ed8ab929c55df40dfbb517e80b8c39180e7ff238e7298b416dcdd238dedee57ca1be467515874077395b74a1a4d32ff0efeffa8d98f51725571568d588ff3388f475ba8ee9c0af58b5ab6e46184057e9fc9da9d152c5abd24d30333962fffa9abab6496ec1572d01e8b1b41e5a071f540c7667dd24a3684be3a955d0cb517cbe7540f6ed19b4c95806620f6227f1f3f59c876cd7402e7b66572ae46de9c2bd8ad83bca5fd7bb332c55c033a2b2f9c079516a271cddc064a1e3e4f46578d361ab44c3f68fe955767910ee74950156463e07a503f5ef77fbe1db63644c67d607115ec07793613918baf2c805ab9cbf8a6d8eae32ee809514533e08c24bd123d8914a354e7477ded6ada8a93a7d71039dde0911e51b894877c06788a87d8bb14e8b693ec54a5441f0d58aeabd1488706afbb425aba2038ecac759de1dbf27f0a680973e84f29c887603383c9d9ce87e155631490d7443e5b627720eb117f0e46e87e02c5ab22fd86fa2504bcc2d9fdd67e9c688cb84c1d01d6b1a62fe9c463c237cbe8e4790f8eba3f035878c618a3bd7028886eeee9c151d39f4bc0eb881eb05a956055b6ed8fc9f700496550d44751cc0c8aeb5f11936ce15c7982fb7c3238145866e1616cf7f5901a3652b343faf42cbc528f6a7a7fb684b88e4693bd51901028881c504bd4383ff2ccd19b80a931196898030ebe202d4eaedbad76ce7cfd14e25bc2baea471eb6fc4074d482286b6600ee6ea137d4958b0a642947039eabbb28ae979872ed5c41dcc6160b6d41872f5237b6a5bd57f199f73669b0f18eabe5439cc43f7d121524314e0c0911e4d075f478123e509580f2a14526b229644b9f67a2411385c1b105b213cfd8bf4235b575c420b004fc5f5d07578a5356d928d63203efe6b0ab7893953adf14de1877a1fd36cec2198520d325474e8e478ff8bca77b74d9a562657aea72ddfda8e07dfbbb408efc07e4e5bee9d170f03bef19b24e83a995dfe5eb9359e20dfa3988be9af340da2d8c2c7824a5c82f68b68db820a3ff1aec6a0f124be0ce2aec089ebef3823c9d9cfdc88dc2d89bb6b0cfc714df469aff87dc4e7a259a3b178ab99bc65936b2dd0a47fead12059a928046073a57b6d18a49663b7b602ae900e853635dbdf773fe909809304ae75cf5619e5f64ade9d8bd72362f28cae84ccf8bbcc7be9a166c04e521735084a261d6781c3d11f375fd6425e24ac75cfd15149e51f3cc7b2be752257d7dccc926633158fc9dbddb00c82406b0fd7ae0e900fc18c430f565809e6b8d84aab75e6561641f9a20189e6646dc162c941d7a0a8b1663f119705277ec7f59a21a59349ba45ef45b15054c24d2d7f92d7a5ccd9be72da80706a875e268c1bac8c37f4f35dcf0c351438c4a967;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8d4af6b6b251d46853c78acfd3135906488754f23761ed3ae60ed4ff2c6e828112926d546acc36170ca7400e1dd21dce739fcd03d45eba700b7849820f1597c7f36db6115b2d0d25cbf95c467dbfdfeaf90ecaa18100987e4fd31575b7c0ca60b58132904752d62302d9a530aff66251cbc45e0737241a1b03fd2014da73cfda20c0d30e586d794088ab92dc519cc9803031889dfc883dfe4b8631bc630757dfa6c52255a16b374a59921dd46b798bde627bbc897544885703af8df57531c55ff1abd06a8b6729995486fb00d9458a765d41944ce27c853b3e4750f0cd1f4c2b567735e4709e935fea2589f93b8e15e430a0b9453e33e1e1b5cc7c5f4ff28974a1b23917ea85031611a6d403ac223f97d39d3c87396b49dacfe57441bd20774a7cf7caa355bdb49e7c6e405c205bc4a95d6f9dc09d1bf39804492787acccdf0be18396bb4a6a13079868aa728f3d727c09058fe0f792e6a4d3819dead8d6f5b45987bfc5cbfeff1011cf9690dfbcd481f72892273bfd49280e0fa79b418f7f4559a3baa4f62dfd852e6f4dd7605378db25e82896dcd8edf7cd61d7e0070f41f142fcd4cc811b270fea48b546e1b75b2129e4aea9ff8ff9156544b604d270f32815165487bc56421dd553c518d01d6906bcd30e831966333ad9aec1e2992d0901d769229c153a4d257c62c20f0fea4b0ffc477bbd6981a52ff3748db6fc2ddc1070d77b021ed96574ac07e984d9aa798e1b8ba9ddfce8086c6be94696459f891c3795ab5a1ae9ca2f23c294a21610d6bce3185a2fffa388b0de3125e9522727c186943503f302daf90fd938beebc521d62f65e7a142494e4f89eb856fcc5c87a76ae37d52069e5ae14f37b7407178286226f3139fd0198aaab04beb44f8c61f8e9b937008ce616fec957b43c70d2cf4e02438daf1f51be5e200bec1edd91ca3b46aa67917c523830e2e41e68352554f2ee6d3c606b5fb751bc415610f19ece60aecef1ea2615ac725a215033fb94f28591162e3c804455fb74b2f6846ddf6980be568c4082ef58222c9e16bcea6382c348d8b45f546c4f0f87ec8af5dc4c8dcdbe6236efd907e792927e68b8fcd7f4e9e2f636f630e5fbe75f48551c2553d396718e0950317e3ab769c46a2375704b59a172d80f046166b1c76bfe7d72f58bd08b2c3363f41ae7c41c99fe66e7846e5d9870c595aaf77775455ca4f2a60805390fc68eb3357daf11f7911b085a757232ecf88e5dfeb0c4d4eadb30745a49e01b42921613dd598f4389b96bb56dc6da5e88ae5dade2833d2b573f606021426c8d60a4bb3ad6ef146f0c4e5f184c2763e74d862a2e9a1f0dfe451672545bde57d26fd654dad46f7327b659ab1bc21d9cd6636b37e7e0d90b948664e1443b5f18e7c750d383b700a08562781fb3f8d6189f6590f7335236849a0da7ed5d6e4f6a777;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f19037565a885272b171c1e1e4fef49ff586cbafba526b3a51858905727f34f73c6e0312ef83a24793a836b398ae751b02ff52d2ee92ab4dc758440696487449abf5ebeeb90a84a16b9dbb4a6c90046c189917de0009df724b008453d16c0863b0361fb465dfdc915f80336973778268c4c1352aa29dd3ea9e1978d02cffcec357ffe1902ebad7f02e65e31b6f34fe601c3f412aa520001714661fe34b862cd6126967485fd48530a27c1a61478ad10b64b136e811ea952fbaac6ea99837a272929df39b79ca22deb6f6893f60c491155f7b1079961c624ee513e68fff6612cf68cfde8cd386b09a5faa6898d79dedf0c1da5f4292190498571116d207172d674c82b6f0e9af26025693241b0b0613b1bd66ff873e332130b47319deebdf4dd2cca4b8e90fcde080e4d0a43931c4c6de2ff28b908954621a493a70a69741448dde089877ab1a2219ef87a44a5e62c317173e616582dc8bf6b348fd814afc94f33a3008e046557c403704d2c920c383a6d4a9fd283987d0469eec9b9ba80f51b2ce54f65ce63eddbfdf130973f5910f330ec2ce26005a890e2b22472ef92d0e161fb2f631b7ed37889abb8b6c582f5fc84e9b2357f794656c8fff363db4bd204baf5d867875297aac506796cdb836033d5b25f00515b5e31a8271caa0d0f3b6a0e94b6aca6174a6d2e1dae9e0ca224f0440ed4662721edf7193827255be70a4c2a87aa6820059a577f55ccba94060f5c5390e83b1fa3cb375d1b5faa7f696d3405fbde0cdba0cf41376d036eb63592f61d24147358517b0a65aceb2ac889f86f2c3479586efe50156d4be987dee037c00a6b8bfe0ac94e48171ac19f5aa40c72dd79646b23cbb33da34b6a3c5efc45a39a1dd26f5b25ce54084f6f57d3c179c739ef487e29b23b51a1d7cdc238e8c3a031ce1ac731d9b3d6477361296af982901d79161edcc5978db589b10867e81c47e5725075986a51c71e8b8abcbcf88b4cb118b573263883cf480896ea04177e87f7dbc2fe0db2bebd7d3def17ff08a6268e8714cb8fb2a22edf823f1d74e2f826a9f85221050f46d56f9a6026b6b0d14abc4a20c2953e9ccf32ada36c0d2c4a765941e136289aba9730752987e530f6df2ae0624df8b87698a9584cd0cbacff99b64822de3a87958b1203487475d79caa815252267273e805c73741ce6650ae62ba7e23f597c994ef5dc333345b5c370ea4731bc59d63b705eb0614a71d169fda24f388470377742c12989caf8fcd71e70de2085976c88130829603aff3665fbaf4e85f7f2fd091241c96ecf1b5d5b14832a194da40529b8c067a2742b02ec1f164e8450d293ebd105ddc7d28ac039515fbe3f40c0571e74bac5e510e7bc0dd81ec52ec543d9eb650a21aa214c0c317c99238c096d0960863d34de767bd5f2140aa7da6214726fd29466c306ecd5cd749;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb8e8df545d6311e1cf8b08fe7bfe1d8579001ea4928d6ec9f45eec044db3791ee9dff4b7f023c0f94e04023cfb836be896dbce3894fe9da0bb387bf46c2e826cf09b0eedaa46e832c8b8fcf17b0d47e61de48caf8230bfdae1b93819076eef9396b954ad2c1c3a1bca7d672e8c590159a885e0945dbec74c358c077d33715d89ea7bd354e2d07ad51f2177be8fc458de9934099a1799670ef218ba783de565c2e3dd80238b1f75151c925f661d7053676449e2159f9b1ae6291a5561d1eb1124e06cb6789af956d81916f9154c1b2cbd3fa3fcd1c2f412d47601987eac29a8cb3173fd5cb23ee63a3b382c7c5c74eae2016dd04a9a846b10f988f9c69248baf7b6bcc2b976f694187c2f899e58787a6060d80e081baec564aa4665a9e5d904b3aaac34e350cd350e6ec7ddb52e98d9ba50f11754c232452119e6c27a57d1c1d961880249b5afc5a0df2df2698e31b30829e1be43bf3bca24c8898f2b7ab1a2a442602fb3bba57c8c0d6ce4bc4315d039fdce67c3c743fbeb10b6301175db2d3f49ac4c033ef82606024f4583890e7889d91e3c605c63ebe45bf853a3b939ea0fae2d1506704528eea3e6cb7ee824c12521f1ebaaad77a16c9d089bced374546cf6562eb4b3df7be1f6b13426df8cebbd2fcf977e9fbfcb37d40445c3f557753e03942537ff2e7e1d23f95d12f05f148e7fb452f647b358cc5618cad8e99fcfbf308fc6c240848f8f2bc44b607cd11a3f3e93360a96b2c9fd12f93f1ff5ba4f3a37f636d9621729fa50f35dc153b49eefe34c740870e61c76362f2a271cacea7996a45f51b6989dbc878bf2f5018511a502779ba4ce9b8858312c3cb09e8dbb521b725257300252e1ee349d2e54d6ccac561670bbdab3ad0db59493e3cc510a6f8c644397a6daf55bc56fd788070f5bd536286a702253d0b9dd76abfcaab46170d15cbfeee74aabe809340a970c5937e8623b21493b9dc23ece50c90e5808467e5d76e672cf43211b185f112e5b611c1005c13b60907110be0bccaa890b002924976f36ed0c887505fdc1be5e458013c7cc2bce10222714a6b76e202d40c755876ddd0cd1489de153736527573dc87918cb53b4fa4f36482c9fd308b037f7a9d22d4563e493b55a86585a3a2237ae3fbe872f6618dc8e930a15bc20cf8e157f3c53086737d7b45174166faa6fc373ddb3cb126b56e51a4c08a5d1c1dbde96a4a606d6a87418016d8ebc51384f5cc9dae94a0da7437e4f052581cb85bc6383b194453f01317a7929e7eb46f7cda39ef15d746e64173394bdb1b8b64901a157fafd16437c61b8f524732f40869a1b825ceb2d8b40cc6ab639940b566393f867b285d51e22455bd6cb7f52ff69664a280e5638edcac9070431aff1f4ff7377ab5d598e711927d94fdccba79c5442c4bf051eb3609c9b6c293d859b2164cc330b64b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc20d6b79b503aee48a23089e0248229b1cb60b3ef8b14be5b6307f8448539bdc36537bf28dbc18561d258c4140358c264153cee95354a014b214ebd27b8fc0368d41773dce4179c67ee55a70de46bb9784cffda5fc883ded5708721d941d2e4df8f89550fcafa9e0dbdc227a96270f955f2d3324fabe6f07027c59ad926051c42621b4f261c96206a16e6d489d924ec45ee9ba3a4476e2da353264ee857921fc131ec1cd8e6ac44a0fe9ecb4b5c2354d5174162501263901e63ac6175f3f23a02b0b35cab30c5ded68a0e2f7f9037d1fdfd3cecb9b4cb481287695e606a66dcec764fd5038c0e2567a0764680f9e1e14ce55aea7f846e20e312b5c5d8d65ec29e4be8642b59ec843f5de1400194201bf487b695470748d49de0341e63871ee662b787077dace35a9553f3b55e97ed8635b39a75126684a0ea3e3d473403cfe51e36a70fa78b762d6f3104a1f529bd71466cbf194c71438d86ec9c832023568eb8be8db2c13561eaaa3208c687054c881b8f25eb25f9e65ea1a1cc8de194909aca25e32ae0fc5c72f8bb47ef8652bc18d2140d21594bd4ec0c1b991a344e42d3f2c941956ac94cbf319f54fb3ae56b06ad6d52e5050f56a04705b604e51c935eb7964a5d2798798b876c2fa24e48ce9bc9eda3113e5d61478e92a996def72d6a0d0ad2f7b0512452838cc64792df3cb218c1cebe85e70061089acc8828439b87a9b7bd76de0350e29d7f9b2c051a142839f4d1b9837ba251f1e684da86257a09f1377fbe99b3e77bb09dbafc9556b51d57fa98f74cdbb282d25645787e4f723e943f8cb80add9d473cbf5b10d1013ad0de347b2274b0e31cb7693765619241b5a7b7014ae908bb73d8fb850b1dedc75cd5a0ee5ca6f1c8f2eb09d699f3c8eceec5833429dafbc87f24c13e67f02c9f06fb04f632683d9179943ad6b725cd16c531ee60d3a6542e12c8b67a8e5efc534cafaf4995e517626eb186ea47c83a8d24f51cf8af4a569bd3837dc775b71e22ea9e34326bcb458bbb44544c852da46a7a689b482677a0f874ccaebaa3cfec8c8d4f84c073fe041b6e63bd899187328780aaaef04335ae700546903cf7ad68d9282efb589338a112a1257fad1de53c19821d955b0dc34b97411d08c052f98536f8c911fc996ccf5eb391efec1cd3d264b6383cba0fadffae73465f89ff766516741ed7bea7372454ab6702246ae32149697e4ef1d813e1066e75d3986f1e7df3def1ee262889e7754c0060ad086630c64a0542a0dfada6732daa36c9e396fcf070acf206420650e77b193948bc93d281d72b9df0bb4861b36963d98699e7ea0001d641448dc7e711e92889680924da187830b59c0e2b8102f29ed564ae65b6f11e94ba2caad16a6c73f24c6d405bacf679ac0a633a88042ad7d19090c2cdb68eb9f4e3e928543e0e3aeb9b872e570bdaf4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21a9fe5a4811bd0285ef2ca57166b1967939c00ecc5b7212a6a62f0eccd01df3f420ecdc050cffc59d40acf6ff432fbf4d505483bde8d008d0a22d0f49d3ac1c79a0bef967ee6e556281b703d0ea59305fba933e0ab007787b39531c89988211a7e05f899889a764583e5d3789276e8535b85785210b61dc9522ee7a9dd3967daa8131519b712b4a5c09ec7130c578842218060303ecd0317337460045a65ec58eb708da48c78aa7ec84e2ed338a47ef5930336217d580b112b4784cd997032cd8a9233aded7c5702a2ee32926db1abe1af6165459e12fd2973ff3637e40136fb0c128a2fc1e530bdfd7b6fdf11e64739ea2ee4e898467d0217812db5ba074f60b2160be986bc33eaff8b3400624e319e7e41cb7bdc2c80e480bb725d18c4abb8fa17e77674a495267c7777b01c3286a00a0382b2c216339dfaa007151700a363868511276dcf0da0e5d35f38edb53b7fd0d0402aaf86fd7a04f1266f017cfbd8bb1f8fc71fcc72ecf5f553236d368b16dbbcc8c3ec7dbdbc66b77d45bf504f06dbe9d05543bbd78b2d820a979c5eb9fffe57f93ef46a418d2bd1438daa97df9d66b70a761c507dae91577d2458956560788292ee74028e37558e75bd63636dfb25f2fdeb5af4dbe4c32a7d9a94eb6f126e93dc650295fe2bbe9d77100fa67c79bc78ffb969e8ba578d1afee23019a759b2d7c35768b0479fd5d28ab79eb16f328ecfebb3bc6625c2073e45e9ff20712a1075280da2de021d3b71df06bae24c41e3e4ff68c424da1ebf48d81d9a3d9cc3be576a452ab97e8ec38e394b647c3a95bbf63fcf90d4ede2a5e6143b33c0bfa851e9a7324d387c860e0eddda539ecc032882331336752e4e3c8dd14e4c6b73f1b490693c59dc31ecb06f3218289a46197b0762e10e56fd1ab6143c36e0d1b76f446ba6715efb317cb7f84145da4f288e828496d65516b21a4b519bb3bdedde4c73bd45c83003f052353f21ff6a0673646e68c3f7ade8833d88a6e804a74fa22b05fc756ecaa17c9f59abefb541b93a036a398f34164952b396719fa8e6b6f573f7837b05a9ec000d1ccec8b57356cc8bbd357d1a3a5c3972d359a0955435caefa4dbfd838622fd500a976b4b816c2a2aaaf84125a28d29c2f7c7fe38a512b9fba55bcc4498752f503b1147559662f439bdc9ca444422e737d5c1ea16285602466b88e8cf8a8f7f66d65c53d33ab15217e527cbb95382e5b710a93290ac02763b5b78c776b5db0575281aca4384f898b6fefa515c182d716e33f8b815d33dd6d5a86c6e18bf6c6727bd5d2eafd94da674379b59fe88892639ab4c76c7e790c26d6f91690d2b6f6b7376aae9561bddf9a1335284961239163054ffd76d774ac9508029ac88e5dd791fea07adb0ea3a12f12f1b0a9f40192976e224ea83f173bdc3ad75a6374767a0f6a5f02c95cf97de3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he2147a2156b53d3400c056cc651cb70d22c00fedf7f300e1436b4ce9d44779a47a5f5c54521b01b7c60edb7b5a06b977cf82a90c48a19358ca7eb452f8fd9973ea9393c2378c545908f7ff1bba7abbe1a2ec538dbb1a12bed4e33cb4c87cd9452cb686e9165b5a86f6401c959f4da238fa902feb895fe6984c122958aee68ef9676e54747944ba384564c574cd98ac4d8c33a5ba9a6748f4bd916da19600bbcc944d5dbb1495ba1681007a2cec034c0242a2f6c0140126b1f85c70ee40d92432a5a7c9f11f1cfbc07a4248d3207f7cd9688682cdd444bd4d89b1cf8ed3182566b09f32b341bee7bdcbf46b5ed7620cd8d2df3033efb7c4ef30e3f1cef1e21d11f95606dd86abbd341cc142d3bf0146f52c65044bad48fcb7ee229835e5f6b0c27cbce949565ef7d241c64fcacbef7e9141449344471aac9d12814e119de8545245bac60aad6a05b3f041df4e681fe9df953c162f210d0f34465ab4ef3a0edeef8303fffe9f3c0056cd7b33883d817822afcb699c1ae0370170a2e28ced15da6bf02c129ffb34ae88d00131389afb14ad25194868b43e5ed4f516ef139ce9b62e53bd057461e63b8af34f01301346514554a8978a4d858b47345d58676059ad64defed076a14f7bbf70c12a2fb38eb5bfd81c7237f478e0933093e1b7923fbbc25bf9abfe9fab629040d9e9ed886bbb62784f0d80e2af8ace95b1b50c9492601ad0005e56fd54ed0161fd5b074b4e4d04ffdd641744cdc27e0f34f330a2a27805579b9fefad297696ec7890775fe473c69a4c6d9ca8270e258c63b29739e1c81031b9939ef3b3d052eee7130373a099f8f998a737135424a28f770b03b499b2b87eaeef9c603731abafea8b380eaeaa3efe3159cf25c5ac77d3117c58c52b7eeab24b5c53c67d086ccfc36cda24aecc4bfd26f352b7c8df9062c9e34a8e9d008aabc50522d39674f1fbac487673b5562d0440c4c5d2cf8fc6a478bae6b57c0f7678efd549bf13e2945b1b7b2a87caa6b963f3eb45dec9b1fe118c1fcbece99da3f81f0b39d46ead5adcdc7eb3fa37a9a4c2b4a3b6022e814a8acd29d868ab975c43e6c450db4f4ce71d06493c401be44fcb32d79ee018e272bf56c16d76983c46006254e1baf3423a9e4ee13c1bd4bab0838a00247763a21186ba0754f5220895b54cc1b85235d91d694fe618b4dd4a71faa99274402ff4ba9505ebf78d6a7e178760670abd91ac6339b0511c71aeab7c733293f23e25f2f8537f720af2489ef941d94c5c1559e596168fe75523e82e075aa5b73f041702d042ab4f047da2bd1f056f736cab81c54beca925e87a6181afb3bd85db0f5853db6a072172f0b02408119d297ac9f370abbc0418b211afa0692517a601f2a84588730cd3fca4bc6d0fead9e06f18eb2641a4d2ba07f977a505d0179adb884435c3cfd4ae62e5071316;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h788d631878ada871dda31720387e05113b5716125c1b1bd86789219ba3e41c46953f227776202a253fbcf42c8552140341d1edcb838a9b271d1d33b56c6730030ba4f34b7cae1bfdcbd678eefd49b76e4e336f4f46652af38df7fc0354a914d2097a2ece7d0760bc24abdd7072123da6414385dd91198f3ebfb9c9d3096b8e1ab9cba1912366efab48c41104b38bafadba964de89dfa5ae98bd9dd13448ddfa85c1e5f60f98ed2b3fed2abe3426467591c11ccad50ec40a5f04d9a69d8fab02e8ca7e8ba67e9c4c34004552ab81815d844d38901b9bbab134259edb7885dd412a9ff8288895c40fa311e653007fe2cd68d42b8efe661d8265dc8316ef5cec21a6f1ffbb1017e59dc69ec3d39dd5073ba3fde1d24016a95ef43b8d104a959d741c8f46ee70a8fb8b5e8fb8e4e17e6eb431bf558944f4a7aa4c9880e086b7ac8f819328fbecfdcc7ed3b054df7a19fc13ac1d01508122ec9b04e448ac9e13afd65819c80c095fc3b3cd5de76eaff585815e0d68130f196669724e74fc318b2c4fa318feb263a90989ae478a0516107681858344787021ff29c6237dd074231d5661090d3057b7d8b5d9bdfb68dbc5b4d370fce1aee2366ae880e92ec4b2748ab3102bd6015d4982d004369e94b27e20c13be250fc41365d5f0a58603d2067c2a2a9fd33947d7f1a7678ebb388e9c079ac19fb98ad8113ca3220aab5d925c8c082d5a1205ec1d36aac3a2aef2664e2a13e2c3b474f360e0117be073f55b786b07a5a10a8f473f9c4b84f1be09b7adb28e96d01c8185cd77c0551cc3fe6d1b2d090bb07fa937441319c3d7267aedc0bf4a39bc7b359561cbc4750e6e98bd46d353e95fe8c4483240a12338f5173dc1a484afbd3b778d9a573d68c36ca3975f24746ac3b7d0f7b0c450dff6570326708608582de0af8dafbc2915e706f990af860038e1ae30231a16c0198abebbc99401b99ed99fa090dbcc61b810af270e3a8b757a04dec9710bca56adb8684b1ba20db0309f8e0bcca4c180ac25c4783fd9ff7d8a975a565fd718c4b6f686328de4bdd2ff7095bcc25b0065e22f0a66e56d3b667b881a263b2cfa88b50ed13cd6070ccc0ce8910f54ccf82d78d21807040fec5f2200e8b3dacda858b6f3c1ee3a6580b9aa3a643ba8ea77fafbd933a8f329943366ff814f7f6234f15eb26cd320ec4c89d04041a703b6fae5fc552394e0e2e720f9e1f0e796ffbc53b0b4dfd036adcea1de93fd11d24bae97dd137092f90568ebe35204663d0f0d6fd25f0bad9d10eac9fb437091e0564aeecd6ed21836f11ec88184da0a7963a8fe5b3dad5a9e5f73e880acc3318b196dff277dc58ce125dd1725cfc58982ddd177ce68d2d1047bcc5204ef3aaecd1a07473eb4c49d65b53a2d3e328d3e2fa98782d243010a75ee3f17975bc7bffa23c06d8ee9b3500441881e38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ac70b44147da72d6fdd79217772cb31021f8af7a69e8cc245bf90b3bf2021242aa87256428be9fc3b7b83cd809167150853144d45ba02dc8c052dfb00f148562e67fb8b63b54be286eabf9c969a09ca7ec35a1c8977f9c84776105151e81774e9a8cfd82c0bba75c525a98b548995322ef13b7cf097eefb9f3a452aac570c410739ba90e7116e845600233af9d18152529ff70167fe40d48ac3230061da17336743cfe8bb896f1329ca5d829baf1dbc13fdcd5e7d4254ab0ee336d9ad6979245ac21ae1d2ee3dc94904a152f5677b5a0eaf1cecd79ad30b669d0f871072392c43a8704849ef67ecd4838d32e69551f405e7c24efa888cec0833188fa5c42ce06f836d66c8ab8499fc3065154b73d6729171bc580dab0217e40b4200497c9e5af400ae3839981c7219f6cf91802ea38abc5f2044ba203813ab9b97e85c58322b3a935b2ffebb2c4c65fecf38f24f0eb3a36165e31b59eaad62c5af6b5e39530a66bad5aa7b4cbdefb8a9082c037b0215e7cd5d6510af449c0e5959cb6cd5b61cf4df95d1b36e9281b4e27045ca9ec9a748a4510b268bef190b5c6967e38c611ac3787ab65d2b332b0f5cd711169e7b38cdae7a0b3623795f748f7fd3683d31431239c540230292fe6d8c57eaf490568a16e05c80972ff952edda40a63d647118ac70bc2bb8ee8faf606518aebae4e090e5e215deb79450d201579002b3f6f610a6ddb9bed87552345ff0962d67c61824e2ac9cc3a757bb2613af014b37cacb9ba34619f372ba74d0c880012dc8146d789133675ec3d5b74f87a0d8fe2b44f018aa37ac75a44727f1ce79b33809e614cc497f4b2bd6511b52c3ea34c779f9d3b726ca3c0392622ec43acfd2597d5c61141c852c7b24bb2b6600717d7bee3297af584dd26f068d29ea4f5627fd7a483330d2dae04e146312dc34e90e60cdbed71acec97c9b3cca3a76dc8876c8b05498f8133124b40fd40095b6b6f4b0e6c308681362c3fc2596fca70097675125c7abffeedc00478c5ebd77f5a1cfab59ecef954c9965b01dd142a4cdee9d30a20642afe8b14cf18fa169408806b1549a9b39ed31067feb7bba1df926ed303ccfb6d11f12c5aaa24b788788257d062c7c0b79704cfe655ea79cbc18125c65a29383fcc8c511b7064b277955d675593a244c4e83dd4ed31d12b6901ce67e5e02a36291333372270ffa2a3f95bdc3e672207113416aa48316db09968b054dc8f6755f146c17d2c5d4beecbacc7070255b444afd706ed86a1a00ae4e8ce0fce4fad6f10c935dd096b7150a34e4100a240228115082c3ab2b404d405e6b003220f820875f5b8b83bcfe5fdf2402d447eca0bc5ac7725788ae7d3496936361a54843661edcae654d9a6c7976ef64d75aec5873c3f03f2d02f82058266dae2abb091927e764ad6984ce2855cdaca73df66a295242ffbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52044262621cde384367e567189148b79c103a84e168a05750416876f01ce0962503933e6b26cde83ae7463f3f01ddfcee0d5cd7189d1c9dc330a612d88c05f0e4e17e8fd6b6f8301dd72b4de3213e5f7be8343d80cba9efe72945e8c32babce4f977f798c8794413318b9cbf1366c5bc4b1fff9d4dbee4f1755d7143bbc43d51d490949a72ba38035bb70fe7496e79d80c2e1061cb7b21aaab73f939c5453ce70e28ba1354d4e71e0bfba18de0a2169fc632bfb2e898f48e77377640e453976606e5683719afde5fe290337f250138cb4e8fe08e025a89e25e01fff84690a1ef2184cf0863120bdb0038825f5552ee62e23fa6bb97cc971596646c85213957f57ae783426809b1d297c20152b6a2652c4e32f67d3ee697e5c94d4cdfd9d41412b2a39bdd583b25941b52176b1c0cb469153358d0b36cb6c0c9a8e9f3dedcfba9cd4e537db212f9881b5ecf0ae9d375d2db7c9016250e29515ea87b6dfa384c7efb49d5ccd7ef7065927ef52d8eca5858ec879df036cdcafb684ee8bea85facaf86d48f80bb2d194abe9cebf7b16a23789d8ac146d14a45d3df900aee1c4952c4d71ae11e3b8c6f297aeb698880df6a4450aafa3900a4ab62dff12e24d54f36127ccd0af6bce4a81bfcb1bd5c2e11dd479453bc3f34390bb5155eef1d54e4eb8cbfcc9df14e266b2a01cd23bde8ec63a759938235f364d5ebfd12dbc27e1363f1d6bfb99d56863928404f98a6d88c96974d8fa5b72536cf524e178eb74d1c65de2a20171274eef2f19b753358dc33aa842157fa5a405571e523f92048d84d85363aeee14ec4c28c040f58fe1e29be3f76566bf92378f36e7b335ad84f79d0e9f8e1855df4715f16bfb0e45f50d08d56f9d17d3fac4f0d840c254e9e081a96e38a4a2dc8f2bba978333852fe61797c0f97b92433ec96ab46e0bc684c012725b9db5a96e7cab88a2ea25667ac4c69597326d60d5acc7f720bced06cc7b3d3e4ed362ff3437690f2a189566a14aca15cbaa85ae4a41d76b9267445167f352dc39be5694f2dd897307208a7cb9e75f07bee6abea16800a061dfb3a492b914a54c1ddf9bf61730c64f32371c2f3b492917d2b122106d75a5bad203d205b80f91480e2f55809ca4559f495f4ab93232af7bc443c4e7c441f4fec2bc6e2928d31a5a52b2e41cfa65671dd5abff5423f4337e659b82f35c54c6601384616486b7f5e83dd219a7504742490dc622d72c8989d6590e529c8ac721d43ae221b1831d7978847b17231114ec5db2e642ccb49900b1589b91113856e1472c32d3c0c48cf88feb83bc22e7556cfe6a95588bddcc891288e1b9c1d1653fe04e3f3066d64fa264119c2dd3ad4bba116d682a05d2976d1a5bcddeacc32ec458c67a7a07ecbc8a02fa8a29008168dbc477974aca1a0b822e3bcefc2ceba2bca7ee0f59d8afa78a81f47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc6ca2dccf130744079b056a454d8dfa49c0e38b54bad29d0025e0fa4b2419ae92332f2d60b17e2b3bb9972deac1691ad4d07e50447acc8555d56805b12d42e255e0d5a04ab1e1026513b7e7d214498dc88e7c87eda30dc61f30cc1cfb13d21a602a08ef261cf0305d3c5bd8c81aabe7cd759e645f05d48b0909065f9c5904a042d14a57d8a194f91aa8760ed67087a4b64f3bcc9779109c58c25f1d230e2e582e2330a40961ff3a6cebcaca5dcb8e19508692d1e4be0940a492b43b0125d9b0c80a9f1e78c50a9cc30b64d45847b5bb237dd099869f7dfea15eefd3386eef07d3987b096c914b56cf5c67316d22daac03264ce3c207f087fffda79b6bbf1c9937cefc9a9e6ad4ecd617185fcd2079a46523d35e2d8a91032ed06cea1c82f0b3fc3aea09a682d6eadd41f38db837e16513bf9cbfc5dfb93c1021a34e04ff4e923fdbbe1f2171cee7157f2908aed13f3f467fb61aff74c9da2e98e3602bba2d5f95454b16a72a144942f24ee6dc83d37eb6ed6a157038c02ff44a619088606304a740d3549e2bb49163e9416dc52fda20c643b4604c80cec15e5120d6afd4ede527ea88e70adb4181c7eb0d84b7b4301a5cb1afb88b584f85ab32d5da28efae3267bee2099b69820a4a68be472a15a1526bd163e2b3c6e0fc0600872f75411c61d3cc69f21a61852619a3d0c6144b3c33cefd6f8144be297792f2a562f40bf1bcdf3cc279e7a32582d24ed7c3c20842dc57ce91c9c14e3d9b30416ec0276b5b9905b986c1edf437d46838434872335388d7888d25aeec079412a83e5c7bbbc1b1c9a57aedc110afcbfa97272037928c7e94550dec2b74be9b60ad632f3f162848335c6b482c7c4969c64bb4ab7e3e87cad7c2f824a1d845275c7813b5231431669ab34d382759023615b591b0ffae9e8776e4a9722de432b23a18e3dbcfcd1c1103c32e405bbbca03ef11e6db0bfa5554e5a358e2ae27e74c6e0713d3ff8574237d42de4336a68a0d1b00ab1c2898e70282123efcb94de75b1f6f1d584bb6976da85bc48ffc0292266be848f7db73ed6cb490e9a2fde03342c33eba833da8d9e7e100639a6d84d1b22b4f4dfd0f2c17be11d4f604bb3726599974fa5745fbf119ee2f7c058b6aeefad9f9bb13cef8f8bdbb3e104e1f36ab0e48b777de6df580bbf500b94cc468556a48d8ba5b34b1782ca423b254e29179ac6bb56bfdf8ba00a520e05ba045a06a9cdde9c63ccf5a62ae7dcaf5d53f63d15227f9459324ce779d8fad8e1216e3350c4e38c22d17800b8c8c6f4faa2a111fe7d987eee664397d235fd92308900e98a7e642526ba4a51dcd1b65fc7f1d9e448d8a8c5752e53247e24fba96a7b112cb29b6b8a99df46dae9857e71bbce573e3c9114a911e6eb4cf5dd6c8c2fd39e1454b8e6d857182d230a164ecdf158b79353d1eee1b02d86867d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h29a467791295fb24afc147fc6de03fbbd5f65cf457ac3441a8de31363dde68d21d50c620d8f0e09f4db424492cd1282b8733501591f5be8c7ac0faa7b1ddcca704acd77ed3e9393d82789b9b35ee36f515568d0c75243cd2cef801d72798652620a5f32652c45c881c81460aaa224177e9e6ab751aad805d1cac8b496e9405fc08de9c74fe9260888be3375361b0b960a7f8416df8d65af59cd0b57dec5dcbfc76628d90e1f40e7a0b128c1ceae53d078681504e8ee2e843fad269738eef278ae354bfc8238eb158ab9302a0132b01772056f433751fd4931954b13ef73b9e1451bbc3aa5c45e1a8dd5100e4b18c0b2260788d4e48c09841fedeb3df09892f8042c398f49a07a3a472ea9a62d7236387100e348a7a495ec0724ab2e948fb4700924cbeb4d105dad0f86d1b66bbc83121af39ac26b93de60a4d7a0311fdf6296dd351e6b67f3b4e2556f82115b7404e4e578773b10b9b30510634762cd44b04c6b5311cb8020d0e4a9978e9aef79ec2afd19edb6b5f58e6e45aaef5b7a78896ff50a9654552ec628de30ca3bd0048a0a1e6345e79cd85d7da2abbd4aac76e32f66ee2fe3536df97a8bdf2f9a958572d26eaab5b0fe7a3f3a4d4e068ca0b3b904f1f7bec5d6f318adc916e358fa3c9745a1ea50ee040dc4e2724a8bf68f61f1bedfb34d0fd13d357a013c0a43a5be70e934f4e271578f326ffd3726b8d955c32bd220c89531d158dbc13fedac74b23a791b7515e403b296313c2a06db184944fb63c3b60022eb380438bd3f4a0b8fbaafdb0b9e4b3316c239e9e28d7b6f5ef66c76fce5cee2ad63fec4403c4a939e39252e7cc76e6de843e40b54ff4b986d60574e89de0f8d822f1926a2026118115266bc389b042992696918de0a1cead782da5cff36fc0eab6f8e3ccba0ce98b6c93a690196f169a6769d45527d4755ca5c1ff24f09bac4217f70b1482dc21cfc68a9030aff5cdb7d48298f165883ceb70615b6fd7aa10f98bb65ea1f6ddbf344daab6ffc919903286d08cb9b7ab6669f7ce18fc5af735d09c3d7eb21f0d8bd431fbf612f2324290e4e122b6fa11d2c851d19fac51135979f1c62dc105667a48924a19767017e0d87c41c4b4a2eb9824c0561cc49d125b21a635f5d5e5d7e3d990a8393924cb839a1047046472d5cf93ea23363c162e8254b5b0aeaf766d6db214764c98d8733f332f5ed28645c6448e7a456fb073b3134ca4e02e81d8ccb835fab34f9a12a954e361e25f6cef885eda1bfdd5b3214dc647500a2cd2658ca6ae0e5cc967cd2ffcfac1faef55310821575a9daf569087dd7badca5cea00ab6c0c9cf9efd2c6e30994e17729a31d3e4870a23cb4e65b06303b13d65f579fc39cd15e1ec2eb96734f36eb789c2a81df8fe6c2aa8d8eebbbed17cbab1738dd6801190c7d3cca5743ccb45c2c80554ae348a8c4f543;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfd70faced7dea8cd5406b588a8db3b7e223e618638b457af40df530160ff54980470978d9ae5ffe5b34591a91a1024c7b4f300bf6f018bd170b5144797c3fa737dd49db57538b90c08d59aa71fe29987e675eb9faa52690a269055ffd4d30791afa1a46588ff4e9dd41ac8f358001d29b1d7da0a6a2598a5dbb16837d28553cadb7bb04c35c3094896c4d657b35d883f4482d16f0ca17c46cbda028697f47b6271f8b5b01e030d54e4191a59cab90b1959341ba86144565db30087f73d18c422cd0d1fe7242ded5906210889d3d2c5a58ef1396c714fafbdbbdbdc4fd161e38d69191749030968d354edbe0f2865e2fe81758e40ed73ae4abecbf2a4db3c6cef2af43d7de2e2dc547058a1e4209b68af4a8d7f7117cad6f7e18242b3d0ecc449708e367fa5b0a353ec5dbd7086591961d5afa8f6fa1a32f143f4c371c7101ef5452d3392078085327f9389c469f18ac59f5f345c7cd283b025af3c9c178bb623167593673e44465542644c3aa3a1b5977ad1fccca7d16ea9384a565ee1a57705132c11fb96849dd77638442d01e8032e68f54f37463bfc8f320c6c24512cb73d3835cbf43306ef9a35194062d869b393cc8d639689e4480323f77b6a5c053a7921142662d6281c2b649cbce9c5d45c37c7f0f307110f15868e65d9121a84b2705eb7ff656311df460414a016f5c96bbf8c32b742e057ee35ed5d3c03b98a59ceffb428af6032de075c4e6630fb773dcb3b0c0f7864d1a1898b039b05bf20d6fc9ad4186a13ccf12f686af88e2daecb4013c1451208557b618a8fe46aa7a10726402d07a72d1055f07577b87a600ae03004d284c7414458a4a44a507d66723c08eefaf5b401ffa01a663d8afa7c7c989d318356c7abf8eb8d1503d41a55a07b8fd5e50deb121b1002f10be470240329f03e3a69c532cf94e72f5efec78d462e35b144fea69411306926e8a2ff0fcd75fdf24c5fe19604fd8d21eca1e903981834d3dbc63c45b7c9f289e141044a9ba413d52a9a2461363c609de6276e29ef9cbdf023f8c39a2c42b7f41f7ab8fdef74472e8a53d16c1921a506ce641d1a53d76f00fc78007fef813ac9912761dd26fcb78a2135b18ab8c4793d54db924131a44e901d0d566e916f4edaa110844eeb6855dc34a6d3f2eb5eac47f88e005ad28ed8d23f617cfa1d767cbc59f035224348804900212d6db28b17fbaef36df50cd717b2266223897d8327ac2fd1480aeea47abd2da2157dbb86701a4017d9b3fb1ffdde9f6879d10495a5bc24faa0630d4a71012772311ac9547f79c70b4a2f968484dd8f2dcf990d30173840bbbce2a73c370ea49062fdf16edca96b93909c96a6f95c8e90ac3f95261635ea716662924701d39ca5cab01f7f4a67ae4586a3f9b9001c5eb46810c174c4d34f9da25e2b3baac2f3d9768f6f47cf2f9d8ad94407e96a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6881330e942f23012b5f4d01c08ddad113b2a3420b8a1eef476163e92e732b45fbe2287e25b28e99b1fdb4eee4a3f927584a90a59bf6536cbd4cbda6be06ec87cb939ef93732c7e083a4c1cca2286e8af31b1cbeabdb0d5105913ff93d5f40ab10c7188ba956541e62f80126f3b4c343992b48a2bca028a8155ac72cb102853d6a93fc8fbaf24aea93f958606bde05bbe12015926366f6ea486b421eb39b6239d8ba02af01e26307c8a7c8c32a87b75685fffb11006210de7b1f16903e7b96c56e453a26d94fc4f7c13a28b8cf34d34d8b3a0e32f9fa97b1de2a9df94f724bbf4a35ecd7422eb63c6857e7c87c41f07428ec13ee2b66617276b56a864f57929ec4823979ded6702f4249bcde645c32820f2f2fecf4c769cffc48d9078b3876e2e8f95e3748055cbaa06ef68c6014cf91b650f64f8a9638476b53ed8d6aa9d807ec3734419e24d1ee6d1665d94fe3d8393092f3bcd930b30d5bd71aa42436792270300d5ccc2f41fdb706e54a6d3842e613afa233ab82a50d4a035f2ee8a719e96bef22804974007d6cc1040474209f0e3698e57452f3eb965829d43b0cd4c3ce59d9c814ccf9782afab95942ea4f4dea645007926b20a757fcf9bbf6f11f8b7d19787cfd20372846cbb4b00f1c1b6a8512ae95e9df51a083b5a2d0b791f3d77ff461b654e12252c1f5557218bd3ac826c4c18ee7532bbf1954684d4e4963adf27c4ccbf8c40fb8d0f186896ca47ae70595cc78101c98a6e45835c3fe612fb745ba2a45f4c6dfe2204859667deff97d262d99b6c3b1a16ac2d8dd586f9787c0ac65482cde1e12c00239ecffb966a420c1d1851a801922dd90f05ca2d0c2bd3139ed376b2abd485686897c5aa8ef9e91b4297915d32b043ae7a1b57647e0323f5299352bdcef9412fef7f8defd0be2d018faf7d3140daebf414d082745fb4360c1c88edee53811a9b1f3576cdf731ba65de033eff7626fd2079053c57a0c009c4d1064ceabf7f874e9bbdcd903a1159ceb1c58cbc8582ef6b717180fd70f7423ed67cf3469fd17a7af81fee247269bdf58100ed486b46ae5cc5b1cbaad38937b9c7e436d93ae12ffca888c6f27e7d4c454596b258d4f9a48dd82145df916eaa9823f25592f9704c9a3556a74ea5c192fcd1ecc055f2b84a68a2b14ebfca7383deae137a0edba6979acf0ff46631f24bd5fa0a928c938b8699a2cde2d91769765ef2bee7886609026686428f21f0e8c060936a5b60d41773bca8bde78afa6d9dd8a707704799ea4cdfbe650ac8e397c061efba6bfd37e429146b4ea72c9c40e1a256c807ac7be300ea08833f631199a3be8b386e0b50a3211a87b9070ba07a1aebc534e01a78d7d251f9c50cff134002dbc0d9247e923729a8cb0a58b881e002b8d67925d5f7f2b5af25ad28582d7f21ea3bc081b85145bfa4ee9a5e6088e26041f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h500b3ad9658dd286f54161c68728f0d2822c6f03c92c76310abc21542d1d7a98aa31a05f950f11b28d3ec51b7c0891209fcf6c5e5568bc6a3a58fd01f843562e88c303045a9f33e3729e3d0d6d49d7ca0f4c704e011abfb4bfaed52fb09a8b7d29e0a092472884b22883162d98c282247ee719f52610245bf50e02e8189a343b523b09ea160709441e9560fe4c20587892de39cc5963c7b13efd0661a5315f3abfda2e7bf2a6f07fcf68f80b9b381ae7ec3d93052c72456d7976149788f7ddc0391b03d2e215a67390d5530acd4c04654c678921b6aaf0193347cffef5d5679dbd4c81e654c342120b9d9d4af1804341702c3623e6439a2754bebf87149fabcc8e3e37c1727d4b733afd40320dda046c08aa257e59635c27bf2ca8fec626e71ed9cb4f18e4e30a64882390de7e3c9a3ef5a446c0e84339b3dc2bc9e05cc3841fdd426870a5bbf8b56fc858f11b52e539201d162b57de0fdbeec8cd9041ff1d7236087d858d4233d5190fb89a43be0f83b8d41c280a0e827db5aeb056aabee8956922618e087aec5d006d6fcb4ce08040a68cf86a0aeb12959fff4bc13f9d0f6a90378f13ea35e23d3a1a402377f36ec6bff93db85cffe5a8df62d0ead7f33af90d049ec2c425657c49994562d384c73b2ed25971226647ff51656e06de1a7a15487d76e924f5f1474a59bb5b393f7c21251dbcbf9b259b62bd489d9ba88340e01b753f5e612c4d6aeecfe7b166549d5222fa5b9fee38adb8de7ea0abb878ddcf11fce2a6f33db268604d81f95e6136491c5e70ae32596dc5ac02bcfcffbe97493924a33c31608506fcaa6cc23867d213b6b96a278021f5dfaf4fde333475bf058043edfca8c64dcbb0a5c6ff791aa1c38e7df323902396a30c9d5e7f09170dc7cb4aeca68756e5f9c09da69a20855cd580463cc88565dc739a037143698adddb562482b8f336e1626db2003388c6ade1183c643a291130bb0a0c14d167a294a07f498c9a32d3d7563ec03b4aeda9bc9cc2fbeb3d18dfe003583f2db5cdbd936f1b9c8517c27607ebc39c5131d15917ab53af62bcf984f397fa6d561c04221a79cae7b2ea64cb5a9ecf265542be90be7246072c26882ebe3bc1d905f8a24a36afa92cdabbff39df73c90ae0086f4e48684a87287fcde9d9c25570a0cbc859cd7f0c3c81111fb5bd1b2acc95d732eb4eaa85f30da7064922b6601ba7485da00f5f7d01bbc05aa91bb2781b21811c048b6cc1759bc7ec34949600110dca320e66e520371409ab9f036e9d6c3d542343e84dd4e90cbba52ae2c194eec1b2e87000388939ca8cd5d435c64daa7a9479e42ac1959eeff06b2765dcbe1b35029d7b8cbefc5e9588117ddc7cbb6cccce6a076fd5ffb42383c46272ae77a0768c2f123d3929ff5b0257ea79baeaa91ec9af6b7418c466125809605d1b89973b0710ca7b3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h934a065222dd4e4d97bfd4289ab6bcb7c10ed58cabb27446b7712a902dc0967ad0ca3f8985621887e9ff5a88e5092162b69484742ddda2a2c3afe019bc47111656330f8a7e71ed5846ba6c4b8465d1f111ca7cfcdbf925a3a90d53a47ef1b3d7b8c2ddac49fc47d58f70e37c01c7062b7c63b5e318d66e0c2bf3c59e3f347d3827c465abc2e885dfabf3714e18b0ba460df2a08056dc563a64f0e71561a88414b076f62c7394492b0d63ee054bdf232ad359aa32ded789a4e6a9cfd3e8f89ba0ef3a425d02ade606b572050fd7e6bbd20e339e19b95ff1113eb1ff13bb79f5874750188fbc16d72be27b07de009b41975f24b448f86ed62efe70b21d039450ef0d256c3ef01e5dfb91526d1e77e03bd73c02ee7a078d941037e4512eef54d4f447a8b35f6d3b3d7311a8d980a6525e5a78b1397615d751bca999d19fddb6e4a1d7a94c12307dcc5e0b9b2a7ccbacf986dc76549cb0ca9232303de24a2928c44c39d3f872ca2a9abd897e94a22b2c7ef0a1a96b3a07aa74c6197ce34d48a9d6adef103a8cb5e46c56bbb19be7b9c60a0dcd25bdf3ffa3cdc30bb3b8e9887bc75295f1303f994cb319bce6bb7b42d4f3084e6b2636ab7777e3dc756034aef95dd430b43a924d61e30b43223097a131effcd91a44c5cce16264be4a96e16edf13b929cb3bedd3812f91039c12e5440b83f9ac83a17c2ccf79feff9424a348be216042b33151f6fa74c7ab9cac4ae8b4f7428bba47faf0a19fd3fe4066b3a0abcdd69e99c0cf44d08c023d57a3dd0e4d359ed280c3c9c747b22a8e286fe9da256c3e2aa780b9e42427d9ff471ab5329a558475f96f7fd2c5faa76437ab9046f5203ec6c677627c694232cca9138a752ff1858640b99a42d764cf4585e0eab8036faffab8797e288c25254fcec1a104c2b705b500493a8fcd697dd5981f24f03991a91e4c1245d9f218f7fc2607f729ce64971d00e7281648779854f905cee1f9a777b09df0bb2c9861a5c97fdd22f817c22cfb79c5a2d14e74a9ad47a83ba4aa10767643952b7ad02fa11046a8e63f8edaae386849422c2b48f76edb00371e4595cf8d91416e2a456786751eb0751e3997803edb50271aa411426b4ebc19a333706a7e902f85d2f8be4934df06fbfdfdc438c4f7198b1978d58dfafd06592bc87fa2c0915d74c3e8ca193f76d242438c46b2b4e026ee543af243e8937ef2587771e188d0fc3171d7a87725a629746f01f5200519fb851bc163554807f8d98b53bafb285055b2a3218cefd60a87c9b86b5a3ca0d61e54c2aeb92c1608ef3ca15a7d4bf9cdf7f55179a04c47654c263dac214d0164e9661534ab96a8fa19ec0b03fce24918bf07a73ea020c219d30a793d09c2faadf451d685f9cf386e6801e0d875ada61156eadd8f0c1b45d2a2ff4c95154ae787c39ef565b7b506d5020e7a34f0f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfc564552ff2ad6c7f2cb8afdd9de4e93cfc36c9113692bfd2fc9f6acbd2130c72ea664d8e1d74d0e80ccf62daff1fdfd153eff39dbb17b5e34da833e0987c0fcdae1a877044f0ba61472891102e70f3cc38d53db8a71a4f9c71b029fb312983af01d76f24935a95e2839176b3a2f2d5d6d8d43c5b54a553aa4c91a53aad1ce9b6ad72f1bcdb54ac0620a809e931f519751ae020846aa081dcb03d7febd0ef51885b2feb005269b990a15a31169e0f912e728a645665ae77a69aacba729423dcad76b99aa83a2ffe521bb97a1f7e35c9f5280d3180aba68db1932b7e304714e9a64b06f99a23ed5f42f328eabee6fa133c92c0f77653213d6f3aeb610af6c57add38b3aa612faa77d2c1e6b162ecf04d3fac480a03dbcb5ec0268b199233bf001742edb05da3ef60fbaa7604d929a72064ac077bb56cc240f9e2c47efc6208c87e5f70a55b4a31680e7bcd582c3d01b5b797526341412edd8dad2d7cd1961fc2c1c5daf06490ea8b5a4017d9617637cdc8ef15323fae91715f4e9e21904a2c83b173f4090cf8adf8f049bb2e181f6f1016e61a7b40019f995e4d6ebc16924bed9941af53788230ea8d13632cc49d061b41e54eba9a2cff035d290322a850e85067858f0c8f7df01fdef3da1b498cdc278a0cfc7bb485a259e0d78d51f897456eac7ae775a815cf321489a45644474a0d08c6d1fd908938fdc1dde3063016bf4b7b6ad426a377885e0dc9dc124c84390b4bbf88563d8e8873c916fdeb2d14a63e6ee3ae397b48077664e4f2001d30dbc03741a6c0f656a10886074248adac2a7031247aee6f3a7fa2139a402ed553d5b06136ef80bf9d73f9824fab01469b08ea96a116d7cac3bd96730655f3dd9301d0cd5774aca1f51d6150bd842322f22b6cbcf209c4c57b0600aed0acc42ca1e5619093e5374afcbaa7327bd140c8e301566b4d35534d3805a1f65cdf3293e16d687c959d793118e31ea42d12119fc769519814759aae9664f9a5b2a475b7afc03546bbc370d303491ac5b4d75ad30022061e50a191792e16533d5e2a159c5b3b75df0ea00edebee7f0c9ef66593972e538ec8ab4932f512d76b0759f702b35dc6222022dcad8d238ff08c9dbbb05bc6e1e09705cdbd5a97191e4d99d442f712d734f8bab74e4aa76b1e03d41044408fe05064974033ae821b2bd5b086eb102d762b50efb4305469c06075c526da1180d31e314f730c3e7dfc0f2b92ed78bd1490f8b46321a39929a043b4430b553aef7f143d9f1cf8dd644df5f26fefde77634e5d82f023e1123e814bd389974e484b0f4003bcc54a18d0234e8e6ed17f154e1411f6bd1572f0a05d7698aa7fd044320bc7d89efe337a94301a558aa44a14aed8b8e17cae87c199390ba13ffbcbfa8cca023de4679d87ef9448c0e7c517476c1db5ad38438ef88edba7185297a73ec74ccd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he4dfd6c70d943fb608743fdd0496be8778ec2096b8d84aeb4175a42adf4c21ea16ae66746a42339b5abcbf1044965e10dc9775a99149a21acaa93d810dfe85cdeb83ff68cda9cdc852d1ec4cab348e8d72d2a264510b816c2489083fcd0bf3ec99daac444dd5e16ec0bcdb6f1b4db0aa66d14057a6eb94182761c9d959dd29c7033bfef5c78057f51e392d3dbe0314e6c1e5f64f4b9c1393beaef182972bc9f16bd92e63816f2a5463bbefd0ddb1983ee8f452a18d7c8cdb67b540c5910562710d52fcad4a7da51fb87da430619e1ca34389a0f12196147b68c9269d82e1b516c22b7c61ad3ed871964d376f15110247c4d215d08735e41d5004fa94940d349a5ee16368f15ffd7f2bff66115de3c5812caa0edcc481b4cca413208c1ca53d47fc56827c3f34a0db2d6d08335db5211c68d7b632e1a644484e9a7179cc1d4eef1c136475e12c94acff58f188552aceba18c8b19fee87bb776ec5a4830ee5154a5e00c1d21910ff09195ebeb86cfdf4bcd19de627642f44d2f7816a8e82e9efeba069a06beb5d450d37a308185475987ff4c6e983095fd197f4733133d5ae50c9d98caf2892a130aad65e9e62ef10917343b87f4260f94536d57dc90749e21138aaf2e80a645df3d452b01c5bcbce4935bfa4e00ac9037498742ed3c00cfd9ab9cd0ab79e122825513dd93027cadb4b13bca6fbca98671c35ff3db14a9cc0074b27d02cd7337fb0ca0c859dd583a7ff9ab41d378dddb6d6729cad3d9c3a33fbd1df981b99e7a4a8ed9a46a8a0ff03d438a74e3ba8b2b844a7eadcbbd757fbe90be0038b448154dc4a4df2b68e0913044e8f0ca366a936370152fe0c8c31fcf3856aae0a2dbabea1df7f5f6e28bc604fcf291f39b31a487447618f118876810f4662c10225d9d18c48621e5a58a816229c531ce6fddf8ca3f511127141e8bd776ccd43a905a65e822eab4617baa644d267c841b63b9472a213849524149ff46376e4c972d90ec5db9eac9c55ab4090f8cedcf38cedc08fe68dad884ebe4da24df03e43fb80f28e721e19e15dc95f9c609d0d0bd7495cb6f9c5558a8b4e543656bf6ee9ed766b3eb06002e0b12f58273536ca87cc88616ddc4ad2f49ae272f4f11090500f523a0a20d03213611688d1578016706e2b48588e4ac91518612cac2938d0a1ade45f8f435a987176aad126b31414937dfdb71dd3506b479c821b5fd518313adec55f5adc51b6deeaf3c928193610c1a22b6a45753366f85b04b900caf7ea2e6c829f0bd16f48fd016fd6b3394387aedeeca2cf638f02a1a9955a38e4cae00bac794b7efc393f312074235443edfa06e2baba1802bec50976311a41b5e455cf9aba7568c7ccab87a93453caac1562bf6f67e8c07fe67bc8770c99be150ad0c4eb092fb01586b4439a3494c6223e2d2868498dfb9289dfbedf2b33de560f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h38ff68a923d789f164cd792b0406610479e7e21a85dbed0dfa6a2d74242e4f9a7ca6596347a3124e84d60d739773b27594cdf8657536f67b9cd4f19baf57a4db4990401400ff91677e75087ced28beb408582da17dc0d5bcd559ef1e0ec13839ac1160a688ef0641c67e35a049544c10f0d83006a1d567a6ff9ca72f54d3b9e4dd15a8e7694edb87beb860b5f3478cd5f44a5bc58b1ae3e7fdfce8a87d8908fe22993b538d51f367aca18b43f2151e309ea0c17d46d0c1f39f1570cf619f74e02fd95e724d449543b9d613a078e4b422c9f135d052aa6ad260e6187bfc8f175187fa037438061127c97b12af892312a42bea08f66a6018faf65a7044cb9b7c1a3616c03fc652536aefac7e7dddbbfb201ba4e2cc5089bc4e9063cdad67f6cb75aa5f24a7b4842b7b93fc34a5674081f898e18c0e6023fd390664f3b51903aceee768f63f9d7117ef60cf1704654b281a5c6cd671d0bb9f63f517aada708f7e767bb477fa7782abe4f6203de9d72eaff5b601fc13d94df4e4501bb3eb7e9a5804997eef45acdf8325e2e7b9780a493fc796bee1131e9ee602498dd5235cbdfc6ed8295f24ebac92a56ec31aba7201516549d6f39e3ba6552930e4b19381b72eba52df7197a1da1570187e19fc484097d9c98e64a49853bed9476fb38504b304aeb66dfe290e7843e70b1b9a25419e88d8eb0d9cd1bd91dc69ea781bbecf5f72a28a03f9931addb52929284ab48959979ff834aff623fdc386ba940b0a6155e59c1167c90a5145eb607b715470839abd15260c6fd9a7e4485830d1962049d1efeedd7ef4de6ff9124599159c5d7e965723ebe008cbe643a1f5fddb8bd5426442bebe8225708e907ef505a9665f843bb5630a4c4c72699cf7a74422ca11a11e3e18525dbd3b838e8d39e606bd7c5695849da8a992866883f9547e9cfbab454120eeaa34caad89b65d2c7f5f987a8b3cf56758a1a65a7d0f48a900e639b7cdc9a8c60260635f2af864b1534f0aa89dfefad33a96d00dd17ca99ff2b2bc9da1f3b8a43d103af050c8b44929c272f73bff3e46101b433966638dbc9bd60d639c5185b15bd9d68278e0079293ac5e306a5f58e59dfa73c286e47e0f6256154430dad2535dffefebf3f76732fa68b22348a9bf804ddede7981159cc334fa8f4bb853d516860198c355f60dc6dac480db7558e2e56eff5c425d31dfa86d2f874bf04d36bbb619326e646765f2bcc18a8b7064b83fd4a61b9c300c3bd16dcee4e5902ed48a87db93bc05f6d5faa9e9db0da891a2368a5749bd0223e47985ba0db05d9b0ea40f730355d1f1beb8ab398627e91c3e2888f183769c6c7357d6f4003368bd8354625bcd01460232bcf8dcc3885828d06c53f596ee2549324ec490ce8bf1c73dc5659521d36a6c53aa41b5862146b09a08e8414bb8145d5b8fa0c75d8ba02b2db8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he58ccd612138178215c8b6bec11d1f6614138a8df1bee0876281a25baced05c2ff770c466f8654a74b7b7538683bab81a400cb2b3c4f1f20015c2dc1125a7edb1323e12330e232fc8ae6c3d037144d9afd90e87a1895d1e7764a7a9ad9a3154b04c406035b13b454b82e438600765e70a67ceb6f007d33586a57f71944540d428e6f9029992379d914fa5844f219c35979c93c023a141fc8aa24e73da9e086b82705510f83e365f61c5b6c710bf795e20f18829dda503f09f981ec02cce58ebde13f27f467fe01c5f1e1eb02e2cd7da830b66087bbb64d0d18ed183fe0a7c8004187ffa50a9395da350617d58feb42dc5a9e44c11eac46f45271805f12932ed8923c2141e70fa788d6872317c738e1769d34fe1d629117fa1e1646a131cc42f8320c01331dd713a00b5b0b2cb000291b90eaa8e3e92d4415a0f2ca6ba9634e184adb0cfc35f8f73388fece00fa16392b3c6335acf4a1b94847480e427f7c7dcf7a0df1190c5d65ba8a6ea22a982562d3e8babd31a5bb85f17285cff6cbaec82b5f2bcd63271f337bedeb04aa7bc35fc7ea9c1dbd1989ad2bf0a29417d33dcf0fc985a68095e520b7667a1805295744dbcf429230fb6741e230de415ccff57c2c9a5edeb6003c2dce5ff358f2bc09ca5bf7bed00aa5583b20a68e327861efeaf04a169f639549dd0be454ff0cc4127f6f0c84b7ac719010adf09b852d5afbfd798e6f3e4a2f897b06edb0cc98525cc3fc143f80745058bf40f92c4b3c4e78d66caf81fbed9b1baf2602caca6c3a770a38099c2b221dc9d4359ce84c842c7bc3d74c84cc2a2ea661649fc639d7b241638356dbd064c28f49a9381b28fb5f0dafaeab87e0392fb339acbe85f07e9d0995af7d9f1a9f8f182b2dc60ff5ab26fee766e2fb05720ad636c0451f74f944e5fae51b465ac8661424ea21507ae8cccf2aab5bc01614cb44ce5568551a5f9cb7803d27f3cf30517196c06389c5a59a95c303750e47f10003c3600f95c38b342ada47e1342426353c8033c93696062356b77a7ef293f8953ac02bb99b1df4bb3e486af7027d6c3390c5799d1e82a889a513ba7ea37c44724b99c65b1ae35d79826b250bd5f45b5f74ed94ca490217e6b8daf51c7326db3ccc9352082e58dce3051d98dda05b0449e8c67d55ef793d49c984f443372085969e8454b5d2b573578564734c8940f96781865704b14c9895b46c5e858468342626720d06ba09a471ce0154518e0063097beebf94deffbb11ad90cbed6748532f2098dd33e004f5d6f59c5f6a87e6713163f876fb7d3e27bd35ffc7d363bf01553e685905d3152efdd5d1c866434730834d703d824114466830e45bd89727eececb8af22ab8a76a4855ba710741b2cd46c42d2207fbc8e89eab4cfb39fb110a2d7933bb9bfd11e100834ba7f830c78b3f96ccccdcb42e609a6fa2fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hab39fe261af932aa0cf0dd479f94c38699c7dbfa0297360972e9674ddc738a64a9ab453e4efbbe972dad09c8216ca309ba85fdd944cc10d4108684c52f4c85ecdb50d57f8184e430ec1f7de29f9ff6ed2b477f76b52901ab31b86e471177e3e2f0e7e05788817244e79295742e74529c49d9b4c62ba68b3506176fcc7d06fd2092254511537c1cf92e33f6101c29850578e64f933cbe4ae20122839d8dca5eca9ad2e1aaa91f5e4ce9f3fe8aa8e3603156cdec003b10d9745601fb4a95c258f3dbccceaf71d0738096348a781180d0532efa5c6429d13f80da334bee25754f1544c1edb1ae55d50242aebdda15eccd3a380400b6d09fc317acbf4bc2e7c49baf9080dcb1a8db145d1323c01ba019b61fed888699d3b0ddd519143cf1e0e213093d6d65ae9cc7c667d5a3efafe0e4535ea1a2cb21040da05467d5f88087bbf0b0d838d3958991a466c52fccbc3c307011d5429ecdaafd37279e85a21a75d1d09b685ad83d2e40bea08f5fe5846b3cf08fb57ab1e312616456763e6f5f91108fb6e303642a088ea04e74a449ba2b592a05f6cd47985f27e83ed0a19577b82ddcfbdfda7c87f7841ab6389ec3795f5158d9232a9157057f68221b6d8efc1c696ccbe1963f69abf04b563b5a10264bfa0ef6d59308652c1975dfc683c21bdce8d66e3c57a82b08452f16a81c708af7363828c76c3141f69718e74c0d7e58015b31045a9e6b05d5ed627f343cc4010c590a3388fb22e3c7d2e0518adf157de993de3b0d55fcc1cd3ed3ade9028b04eeb3b8ef69176d040f54ced1add2bfb07442d8a1d069935d0635d0e5c7ee85f4554acdfd631c95d73b3aa88ecaf3de1f345c314566d2cc15768e5c7c9e40e36a6233334d9210ae2a314cda8e5ccf0d417f2739f089a96eb5eea701900a1cc52b361020d5c3f070b34a349e9a4704c735684579c76d818ba5660b9c086b02cea1b48b23e1ad828d8fc057a328396efe8fbe988e4034a4191758ddaa0df00785b755ef5b50a6cba81e5627b80ec095b9b0372633c2aec2078d56bb7ada86a3cf3278762d71e36e3849623a328e4d4413212af9a2d18852218069e4a846669caebb26bf560ac29589db879eaabfa38c63ad52df4cb72f94e1799be3779d30d70f115367cbb52f84e763d8ca40ce2d8008a3abb49db2337e19fe65c502c49d68bc111a5e119573f3b2ead19a873656d60bf39b8be169d5f788f4a9c654abc6a4c89f16e385615eb7395a19a320165786bfe9d1c1f5308a050f81cba80c3ebe417c61092604d700e60e0e5cf3b5b7605c06c2057e80d3b0f79b96adebaac517eee798deb5b289527a29933ca9c3ae48a0cf59c27104b90a8e36ad56e95dfa910dfd2e46b31003e9f857c71b359f7727e805466a825f87f1ffae62971001718a70853c11076d40fa06cc53dd8f332d555173120784b80f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha5869e0b141bc7fd5924e06a2bc9ee787cf9b418fc65e249e9bc602496bef68aba4f7276d914986f797a069aef8a645fbc3730a457023af003840393a9e7ed4b7ae1459847bc509e9c7373b57bc2cdb25616a21b323f795d6ad62b1980661dc21adb9239fe69b01bba9cf3da5fe0762916f6141393cb9f7dc779fb4d013bf30d26063023c33c74215efbcf426c54d31b42bf4801320a7422c91b4a1994ccde98a8d64580cebaf64b375154ff7933b4aef7b5d16ff271b4223e295ccd0a75ff9a1efd98e50d65619ef710e56847a63e0e944bb936850adbe572ef712b59771c2ba977aa72888f41d7e2d0e624957a78a9357ef0e0eb9aec29554511a1141826c407feac8edc8543a2cb1c4465db448aa5dc5a9cdf9f86adfa1e0d76f01c388bb47f776b99725b98de959e136692a72be7e088244cb6f711947b4b0434586b09cd29aedca9db41e9ef9cde5ada051e88247582e07627589839feb0c7905d4b0e7ba269774a987d3fdf2adc42f5b736da0e56a2324ac879f58585968e018f0e686e9dba3ea0ec7f2e2af4a3fc6b3a5ee8485334dce6d88e9cf160a58c6010012b2ea4c4cb3d6c628529b8b7bd598c15e802347811f4d0dd638eed1e61102ee58b4fd65020d8d7489dd4db636cb074b366a0c2f578fd6c7d17ae7858d8cca84d518b1d85dd3e3ad1f7c4b252ce86999f2f87b22ebfe9249084c1fbc53a73a704baf49062b4626bd56910dcbeb2f05ee99f86e53aee9b625a911b3f034b420d59d97721fa0333979c2b4d637a3b7316f1e9603f3e47548bf6952f2009cf055b13687650151b265c675127212e5104ae271091b45bec84b3222d764f7ddbb4502abde6932bf7362203af960578c938e5f252566d3eb5ffa11d7b597e3f1098a7d03fcb644da54f027f839454209ef52d53076983920c92ec4c5ba13049d33142033e20164473ebbd98da89a0d883ee6ddb57f9330aa0d44ba6bb08e19558c7fd9c9db6c92ea842f5dc0ae1fcf1f33f4a777c16507b318cab1ce345f68054e6c3fa5f3fbb0e6f17a695bb8549bd2d1562ad6755a0573c23939fd14632728472243d15d732e5cc59a613b92806045ddd958047ee0903c6a459da037299bcde31a3864f646a9510dbf1d746272bf0f976cc0b8cd1a1da20a5a1c0d452a36d13bbb756183b9d8da0cadd06be67836a2277435a42985a3818788979634f871d4e7d4da3efd5bd1670e56992d2e356703628a1c92da864b93d2c0e3bd436259929fc07c5792984d09f0c6ecc1cec3be78de77a29b557b741d7b162260f02bf8b89ee9261d7eb96e11ed95cc3437fd7ed181e90ea06ba95893e5509a4ea4ef3db281d7ad1231738a0d85707be592f4e2df074e062a119d0f4b721d08579e8b867ab0aa366a08c61cd9def677e10e83329717673347c995ff67319a727e6129bda08a44f3e9fd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1072d3a6f666ede290d89130e11f53240bc0d8e30256a00658fc081737541ec26d88cf00a0f2008eb340012664baecd01a518f5b9be81e74cf0f5d8908daaad38cfc13b3473bd2b3e5eb41d88c6cad7d905876482c1aa2430c58c36c29f3adf1ad2025c07247f4d0a9eceeea30b9e1b1cf36aee39a367157f628f2068cf3f32ba78ce40f3cd97c13ef69aa5f6c18f8117e07dca2bd5693a91411ac24d156aea9d6794552f8d816cc667d2b38b367554c7723ad125276a0794a24727ff391d0894de5dbcefc6bc28328cf6b5e9e3c72a00af863733d5bddbac64d734d29e18b40c692ba42bb3a1aa3341d5004eae7d3a7c2cdfd84508394fdd072057af8a4d6c26e3355a3eb31273bdc55344872a66879de8972ff60fe1692bc5ebd4b4d4fe2027c5adad6234166f75539700ff1c9be71b9f7ff836048a80e73f9f9835ef953cf5b802bd96acdaf7cb7a27aa33f735edc012a80cb84219a11d819defea309827010c79091d7d72240a8da678a695fa677a77e5261596c9534c3d08fc6c02483f60d0be87a2cc1a27c599739def467d22b6b753cfb136ceb837f2940d3983d03335a9c5c97a59ea9d9cf0c1807d561b3a6247ccc76b8c61cbf4bf398d296180b0d5b76c241d1e39545d03c145486045ea8e9a8297fcbbd6bae9b9c6ecac7b13fc02dba06cf43ca24f6549c8bd8814700937ef8d3d7071a7f0c44b172a72c5d8f85bc51c6b2c9a2809bb45c94b6b05a18afa2d33b5a20ca35222f2ac37b42e9e7d3a2f5797ca93f0176ecbf33a43bf88ea61b48fbe21c7a644726024a9d41d829442ab1a280b649709637b63d966ee1aae9ba0ea210e1dcfc607e3a4618949c2361a97f9c094f9e53f6aaf865482939a05e7a451b267754829b69ccfc56987776f2aa2505705a1ccef3b3676a2a1bffc5d2c3d34a0e868650f2c68f0d4f9ad728e6e60523b60bb3a50517202b6509ccfa1f692da7d283111812f156800880c4a133ca6898a236217f23b5147072cc4f82fa86b90f00476b3ee86bb80beede144887c4f023295f6c9db7d1266e825b7ba3d6db77364814f1e90fbf9d0503e369d419fcb8646b0b5b3021a0b881377c049dba37da4a0c886b09f3b78c2391493a6a053816dceaa0cf1f6abf9e5eba75e56d099f70e684f7e8e46b122a02472c8df0027736b99a4271cad43f126c6b85f42d6b5480257b0eaa13cd42fb2e1ccf7159138d783d367a8029ec4ce667700786c4add19e27c9871090195a45b3a72271b2f97b860443b20a8d790a0f116072bff9c0de26ff19caff7a42cba9d7667b0f9153677d0c78080ec0ed9a3481badd90691e459a6e3926d728c6f71710d4a007017672a284e67b7a8c647e2da65f1f20fdbf3fa16e542fcb82c3e52e36d96a147d20be8891c831030524b5f3b45b7a8615af13b1bb2512fdd037a0486422d582879b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had11ce85828b2c1d694cca9abd0200e0bda2fc7fa027b531d1867867b69772e627bca639ec9538297fc1a2806842734e82c078dbc9e86780ff97b73b4938d8de0d64e10ef072d9710448931455de3ef7fa81ce888ffb85054da30367ce92fb0b8dca5e4661bdfa4b60363745b0f960a97ef7c045e2cae3a7c652b98d4d485ef9ec82471efbab7f95edf7dfc3b9737a328ef7ee3bfdeeefe0afe22a74a82c5a157887808c182758a6b9db91833186c79cbd0495a6be7e7238b08dc95ec8501dec22a32c03c5e85597b63d731515ab557cbf179b83c4d3230ab11a9370d51b7119a3e1c10c11ca8c9e0cb474bf31067783cbe64eb78f0ce725e1dc29e581b5e95439ece421e382b3793356c7e7bfc2261d484ee4ee94cc1f8e9d93a367272fadb4cb6e702cd7cd217d66c116f9ba0f3f7fd76e1747ab2b117fec4efab275f165de4f42bf7650a533b656d252c7cc205c074547a05b45e5fb10bc9cfa01ab15bf71d30e880cc3be40d927f55886e2fc388fb964f9b4614b649525f535b3928f212e38b3839ac3f40e5762329d264f7e9ed06951744ec79331261f6366cb9d70b6e23ae5cbb33c943f96c50c0ee8d2efc6191c331e9b72174536231bb71bfe7bd8bd1320aa045d68a4da4c4a5063d523206650bab7527409b2622d50180b8202c0f99b76527379f0a0837dc0fe15ddaed747f367e5be16d435866c50f459c57efe467cb9848b298b120632b5aa88f7f02507332fc56b1faeca62a49201107babad9be4cdbbacc797bbf9a34462b64691865ab9f5919febe89eb640a32bca43cd9f2ee0c86733312402265faaac5dcecd5517ad45d7ed1df4acd7d5796f2204808cd9b70df8bfb248dab83e6ca6d0fd066b8b9b5d96866553704e5f365c1d6082390b1d1f05eaebae51aefef3af3351383c4dfa112c8a454daad4344d95036c6172ca7e41e915b4ac1da8634bf62ea500b7b3d9f9475cf99920301a1806475eef0c5e1d48a72a2a4992803da061bf0fbc0c5f775ea07d55dbf1fad9fd9ae590b9e054805f5eacd6b7e2fe76ea1a313580a6ee047472daf6442aaa20290b84f8cb789b8bd48a0669ea715258d370edfe18e82824b3e522d2cf8727cf6aeb2dd171f7f4fe62b8a129c185ab3dce3230b3856b8b186bac034a7c1f014d3927c94dc8052aba38eb34d831cf4ce138f3e92e81013b65f3b39df1e6a3ec4fa6eb0e3a851a50126ce3ed25e61e4a515da2606482f5394045aaddcc789c74363efa21471bde5f6beed6621177f9bf608966c5cedb5336563cae164905f5e8854bf3a542a5746145ec3e9e186e01bc369076e510f379bdc93ce6d8c3a4664a337e8c0280a15a0d5a04bc74f676c564a13feaa22ca0129fb7dcee08cd7a70efe524ea38aec0b55345afd35fb566df1708b663123adf207616609b44dfc05e7b13efe2a6b0860ece;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9af4847a9f2f45e706e54b94a2fe03f9a87bb9cf6032b81b87272dcf81682165e32146a8ab3dc845022d0cc3423f4d0b3ded31f00ab23abcec627977d8865c8bd42b636cf6ecbf377bbb072ec05c321a05805106173b0b0ed87e08daa77e0b5721480cedd3a72e4f526caa7d0a2c154d895f8be74c011540095a96ab32581e139525838f2b74327c6480aacfa694f729b163eedaed772a5ae7d458764271870150b9f09c812b3b3995c5bdf7eac5e4548a394de969b9d13cc2401680953bc9d4eb785afcbd148564316383c40d3ad27c049975e3a6e8455ad5421f224b469001e4db2b395698c8d0eb375187cdc56ae29f92b5853ee64ab06daead643e9c470012dad5e8e0b3c50136a310855689d0b50844ecb161d01af8e925938daf888d4b970672307b8088f77e67d5bac0d3b38b78b49ac181840ad34130ff3b8d7d5a076d4891f8789161bf62e42f92a1e5a9b78162a4a366eed8fb66b1b22ba41c0eacfc0b1570a5558b691ecb3be9eb020dfb060c5cf6a4c014c5e44982dc8b4c0ef6dba8587a1256d40e215f17d09d298522cdb692fd63a4bce661fedf7e7233693b0f168cf34c1d11478b183e5f6e1bb05cf27c145d7ffe4cff7145ff975c8951589d76c35cc909cdbad6676300b480ccaaed0de13453883c3fe7816ef63bfb7a896e626ea75274ca57882c11c97674f5765fec6826d1206689d0de03269924cc0764d433c183cc16cf3d348efff8b66102305d3b2d434411047bd5e1861914e8785ee14ead035a6831d7f7b9d501962d2f136643c6e1553f17c90e5f217cbf9f6bfd672f4c31aad1cb19d71770804d0314bc7de47178d68e2120c531d418f57715870d92d9cde234816ef8820896597442138dcca840f816002ebeb638d25dfefa2cac9c1192319d9287d0bac648291f6c9139d37b5ae5714b202227b4be6fce5aea72f0bcfa7d7af78ce3f87e4ca4b15a2ced25f44d0b5bc575d8dbb000ceaadda73f403c207649308b60f1bb97eebc79ef9c410fcd7f63722832ea3e72de58d5d9ab91ce2158d901df8e55dc6435ded3ab8472c2f2b59c66383ac50cfbf826fb4e71865da3b0f472ff96bdfd163b8aa6b08593b2ca60c922dd00cef9ffb2916a1f7a7ef3214cdcc0e39fbd17edc4e06520ba2886ce1cc52866e708452e8a4c60c78269dcc1634e3d5c3037fe4687f45e752cd3d0a39641ee54bc22f6a86292852a562c2217d9ba0ecea36d088b2255fa927694e30ec2c859b9efeb4107d083d5baf0fa7dd1184fd6daa4ec017f96887206b23c679138f5323f7d42ffaed781a4ac9bd6c90877cd0c8a902f258690053d00c89ed7e817af7817654b8a03527ce0927b157c9a041df8f7491742401d72b81e7856bdc23dffcaf39c6f31e459290b3bc72f2a29e82402de6399c03792fa9636fedb4af592f333069807a697a4991e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h829305fe707b309cc375ac6937a6a29fffd9bf153cefcc84056e6e3512c82e12410882a749c3fcea3b5820f1339ec8e9723de7ce75f1c90b731c9aa642740a2f1e161c9bdc06b3b51d0d7ca71d5683956748e2a8d5fc513497738dd8b2a8b344b80c39139c24cecc5de31723e3c613c6f91e58a446043453432ad865214b294f137968953e86772c6abca62848941492254c658423a8d783e005fd94205de3e11ded75a0fbb019e4b70c857b4e30d558457c27bfe295bc252295b77471c8181fd745f526b26037f64665586e12613bd0ca4216e20eefc5340a8e25e0f49e141a305587f5a5911027ec633abce5f7ba811fc256a23844f814c079090976d6adf4251227891a2509a56d382a9bbf86fe7b5c34cb58f0c51b9cfcc930df32e289201b66da7db8ef21d88b02271b3b43e6d6f54d8ba562256fa724eec57493d371eca4dd57d13d8e35dafb2398ce04ed9187ddc0d278e98bb23cc5f83529f22c5c07355220655bd4eae1f28d79338d5898143465ed713cdd43d7b4caad6ecc1282fb0aa3a8926f3ab183985fbb421d431302087fec70677121b431727cf74032642e8ede3594bb887715e0e5678ba6b16dac999e1283c1b53facd6ec6d42257224dc539bfed9d23e2a42f594576c9162f7071e15cdd6a02ae7032f71c28d3ebbf350a014a1d4304678a0805de541130894dea3c451a7bf47b2dbd4195880145e4a36a3dc0fa8600003b708aea0a1b129836517d131b44a4375af192e295b68db0ed4839a4bbbc3c821ff41051c09158a1616eececcf674f723240a64aa71563185b6bcc6985c3f63e1c7757b3dae6e3a43836cee21d06a7ba95c713e0e1a6296784c39084868739631c8acee6ba62a7ec53ae6124b44632faa6740ba36a537047e70e524ffcc87c6605681404edb769d6c25bb3161bc0786c278d5f228423cdf94cf331b3c1c6a0455450dc36eb94da6337b393be4cfd23ed9e42526a934b38dff48d557903ce0e1b3b1275d811165b49353a946a2f5cb70adb0e86067cfff321734b1030058ee2f55d30453fa7317f1d94a3ede96bcbbadc32ba3eef227a8b5bf764e136a9ea49779299f47ca2fc29cb693c8c3823e0eb0255b7fdc9db95e328038346a9af9dd8cc4cdbd91b4eb5320890568ea22ce863b711f3fd5bf19045a5791229e38825cbfa9d4acbc52792d5df12eadb12e5dc1bf5d78393c5971feb9e37b200266b5c1d36a7b95465be531cc3b63abf772967515142ffdaa1a7c6c67d1f8a5f4c9ef0bab5bf931cc5a576663800bb9908285766d3e9234bdf0193f530ccb7df7a68788f1885efc21c553c27c761d8e5e23066268b1466f6a888bbada5f5bbe0847dd9b74cc099ebd57b37cb63d13cbfdc9837e73d59655946c96403c282204ad9c701eebe9e9a85db7ad081495f67937a1b8484e4816172e327f69405100;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he399f3b556816d0ec39b4f8565e66e67e61912ab5ec61489b780c68b13a9739c53a73831ef2de11d7de86820b4f50938e38563aa93e2b8f8a57d7e6b2e3e2fa3e84fe4b8cb208ca7cf5643f09b17029452d759e59c06c267ffbec4f06b3ec7af428b3b0dad06d3d29a038015f97efd58ecfad78ac0d6e6bdedf9046b9bb360e39184fefa24f28c2211db1f1c4725076ff02ae167f02c62c5ef82677e919588ed5e912493a44d15b4ade5917cfb3c2fd8775489ab05a96dda9354911be3f6bf3d87972a2cf76729768386419ba3e9ed36d3b519893c0eb38e814dc704f9bfee663efd2dc19506f9d9a532e7519ac765345d5c7cee2c19f39318d985fabe1db13fe547ac7dacb4d0e65fd919fdebc1f7089f02bc17863698c757cf38683e2ffe93adeafacd2189bcddf5a00f82fa6ae78d48d95def8825b3e2352dc96dd2191dc577a9914d1d3e52c7059cc2680c9ef0cc20e47249a6bd639a36934e6ea7ff77214486f2da554fef199eaadac9e82d5d3c2c2f828ef7da6970e9f1eca802ce7fe56d83bf9d871ddd64a023b6322df1b6fa2d9e4316794598d97622e45d97ff2f133b404a988cbb81363e51321bf54cf2d96c54ccba8c2bdc4e8addf9668441b6d116c40ad69d0eb5493ea43cf5c4acf7dea6e2a11bc8a6e300a08ed083d9620b1d13e22825cc2ddb2a6eecdaf0d46c65ec44bccdeeb8bc52cda78cccc7a1d55678fc807a506e6379aaeb11ca3168c5f5d60a8dc226df01e1f14ae9509f92cb1384c14a37e9f77088802af865210c2f4655dd4d972e9aa541bb6acb2a56a175a762507f194a3a1e73d62d78246d9188309ed9dd6acca9bd6e871efad77093f2146e8073adab937314425e033c1c0caef37e4e040c7e711757e8575f71e561bccc1a9f321ac3476173b66a29363da9ea5090adeab6d911bc70cb87f5b64075ff2c34df940a1ec5a5957d425ae9f16df01421e3324af2ab111e2ded3c3f987d935e5161dd5516c432fa211f59bf4ac9e95cf3946200e7ff0e4b3afa09789fa3df4b9c249f887b6b1c3c21d61fe20f1d85ee0a183d2b14de4fb55bd302cacf6eb7ac38351fadbfc1a825887e8a929345d50021d689c5446c6ffdb333a24bb5d86d5dc60bbec404b167d772c25cd3afbc09b701069a091c9b2113112f819ee5b27d4f1f9ebb0b51de4fff69adf70c572ad26d02b46f98aa77c8a2dccac9f97c8f911fbe20ec7945a220d478be5f137eb5699b8e43d1bd90ab97043c895543d75fac1eb1039b43279e2098659d349d386f18d59db3bd163d309bb5d63d48ebe461275a800e7313e7f5704578d8664fa7285d01937c81f33c304253c001b24fed7c7d03f017b52f411812bfc7c5514d4be695bea95dc6530759d17365d44695a7ce67a0a2f29ea39232f89d20f8a8658126f9f7cf2051f25001695b9b08c13de70c78fb60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5925b20020049090229496834267f0e1f9ad78a38da2a0f82fd3e94a2ded5f255b8b81d8cf5881166253baeb07810f09af9fb0556cce0e591a8bc5abd8daa8876029ebc92a691e1bf56973d09c81eac54f39646eb1884d8647a36b44ca6d0748ac0242d0f6a787a442160db7cbca578b56c77304555cfd4cc5d9ae9f0447735d5ae107de5d51d9770e6dec2bb0140dcb5c49fbffeba0e1e6f4391c901ab8d9cd2c05d53a3d60c27ed07e47605e3ea01af32d1429966bf1f189e3d24144167343dac7638ba0a21ffce6690152af85ac85f1337b09b3e4c61c6a323c2b7717cba7bf5cacce2148884aa194a0647038b32234d064c3e9e09ad33c9bc1340d62a60fc9262756ab9484740fbc7f97e837ce37fff0e6e676ff919d13b3aa0d48ea9686347ea1acb27346a0587baa1ca93101b98b4ae1793eabd950e5bf2434676df478bc5ac88cd3067c2ad10c72039d4eb69a859f6f363d44816e9c9e4b431419d550720fdc2501dfc61cbe4fb7b9e67b077322c94e60a809edf488437dd327e106005e70b59ff0321082f74159cda27f75ced6c10edf20b1455640fdd5bd6dd2945a6db0facd92a19ba00205613bef044579ed98a6cebc8ac1722ad40cd3bb903ad0aec3e1c3de8e9343cc4db453eb03243c00808ba34297b92016716e6e201a69355f841b4634930c4180534dde906805a8fae325dd68b8ac955fddb0cb3b0923200f9f697a60f098527dd5e3fb760e9ae4d308583482bc974d49d64aa28c7a21b8019ad86c476f6b218351c22d250b4c6bbed9e2c7cfa6d33ced8a233ce98dff9ae09fd2700c116662b954d75e5954965678354ec5e928e0267fae2ee7c58930b07afea066c9a1bf68ad0e2ccc21a2b256c8ccb87ca6652c3414dc110bd6d78a5a7845845f0596972ef86985d5c8e6ad8803f88a4f57756aaf433227ee99ede5f8fa2bc171d7060cbc309c400931dced2e9169bb2b9246b779af7555cd3e34965277d4b9a095a6aaaad5a00a4da58d41182cc407a584eab35b425ac6abb8d3b4c41ff4d0943a436579ee8f2e5d973f15450bec51b260b960644567ab66cab835fd935a55b0d22348ec6bbc428bff7638252d58a31ff9f122da571e12940b44dffd08e3a0508569e1a443daa46b0f190506cfa9edb1da77d1ce742bcdb99af23131085582a9a2ba8e8994c4451aa1856e391fd5a0033b92ae37047ee555021845797c21ed3714f2685c607b3eaf3e914cc9a4e008b4d7485ab47536d04f2b8120efe7121aab5064e36d1e7c62113b42a870924c8c3ea308156db14d14f4738e9144ee62ad4c0a8ffc72bc89aa957d348fb38959d53779c17ff0931aefce16977d46ff0a48ca54229b0fed6fccc1c8604fde6f06d8032553dd473d32a4c636c9ef409598e00e3744c92a6d1a71fca0e69fb6282136c47c83b0e33a882b35423a1ffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc3acf55f81d2f394a759479891c66a117e325717b89460adadf1fb6e6471dbd1de7e4d4ce50245ca74cb4abab783670ecd0526d1196f652aa17da5c4286ff09822f5b424575d0bfd206e775f40352d0aa951f3f50ad49dbcca8760596832c5300e6f44feff0cc64e8f4c57eb8ba4fabdcd8040379c94c2e93bb84dfb982184f8c44303aab0a03b1f57bfc7766162c74d94b6b20268e4761404619718bfe349a70aaa75f932a0c53d0f6f55ad11b60272efef85a1123fca7014c323fb582364aa19cc723a528e24d037dac591cfe4376b6db6dcab451eb8326e4f57ed460e3e1a277667cbef1ec7fde217c35eb5cababc6bfb28662f1d84f6285067d7bea60812034c08f9f8312037589872169647b8b53c6bb87f35036bcf45ba74d17ff7bef07657cb9eedb8e341f3af661c6ab66726e4d7bf61bdb69eacb93634946b93e53542c49cce13193ff32e42aee28f62eca3169fceb016c259d72879aecb6eab9c295bfceab5cbabefa548bf7d5a1158ba5d7160776627e27903a9ee21d6e655d41d26457a86371a39e874c4afb665ab075031f8cadb2c094487a59bcb09e217726c8d07867f12d1f29d3df27fc02ee436e48a84955e81ecafb35d00d35323aea08e7512aab871963cfd579a20bec12b71ce6fb463e40785c60458123e01ecde4aaaf8a1352fb22a6207c4c66565074b323aab16ed7a92262dde6d58093441d519345d26cf53507a36076ce3c9955c5be672b618b9ad332cba6b74382d31ec5d95e460164a83965c765e7e898d780c1c52241d92a560f9aee0efedd3e41fa2afc645088c9b7eb310045053d1d0164a762a8a954f2771e95cc0028193dfc7822beafa85fd2a5f1594eebbd6425234332b611fe89f0bc31303d6e24b6e42033ee0536229147bf8ea0b85ae88950d1ce234e2339926a2fb6ae329b52acbac92fc724f5e3baac4b71c80e09994cd16552a9b4d37253fdc536d57fe57e247947b9152f0c091ae40446a759fd3478093bc4bcd47c6b5b5ab1dee3b37df7f4faad44a213df6df315568670c5986967ed95e6e69c6b8ce7d938a738b689882b778c8e2cfd02d067141a51295dd8ff676d36b11108f112dc9176781917e20259ca69e2340dcfa1d8d05eb51ba4883374bdc6fabfb02e1a21e2fcb30b78e15401d80f3f5f83b96367c9c15e79c3a066db2c92ae1f632bc11e966b6771166336cfe4d97bd2dcd349702c56764fd98cc30c0b2e5a3a4780e64620b585b95d412ccd05f3732667823407137e04edac787c4b5c56e36c87e67b1663043389c677335d64fa57e72e83e9f0d2fa282cf42dfebe4287cfd210550a1cb48c82095d6bdb4bdbd1b074a38f9d73b4593c735c00f561acebe8fedc8ff78094bff0c98921330d25474b8df7b68d1e2a1ff62e6a57bc2d1e47382f691e0c718f1e08d807f8be50c58db454e36b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc8f6a263032595cc7768b7e0a97d3aa581f324f1e0e572360541b99f2881395360b936ab16ce30b898b5f938c5094cb41d9effab3d0a4c96571e0d7186fc9d7a0fc66ac491572af86200d81c311b76b8319011fa93bcc968bcb7b46129fe2c8bba513fe943b89c2e5df4aa3e59076ad9eedf85ab1eeb5417194c506b0a25f9f48be98680d2acd1235696c9dfaf44356045aabed3ada311bb3f54c7cafc3340a95f1598990c6b79aec4fa6e65ef14b16446efdc1b517800f4a038c60ff413cc60806646276f33878816bd20f36b6eb1acf0f036c3c9ff1de494974a3076d642b0e2729dbee089520a104b82c146cfb1d48ddc67cdad05ec01cac01692cd16af5047f61d6d0f59df1ece4708cd51a668d02e74b985a46a3eceb5d825744a6f425ec70f563bde500f42236cb38ca0c2a894a828ffed126db19b18e50eb6815f4701813726df426934c868b88f5c2e2e63615fcca3d152afc51a8a2f6f9fbd927dffb75e259faccd8f9dfff9624a383bbf504cec453a769b0fb822ebad42f2eff4ddab3dcce9359ef740609adb9d0724c86d88fea7957b8d5f6c3d6d04109190ff2b17f8f65e8d52837ec220a3a35644a61a2dc72e0b231ab96125165eb01d76217a33b5886705b6f83a58e4401df52ebba3d73a322cca6539a97236deff1751eaaf1f701855ec6525a712cac015e3b8b5bd0a7901a0b5d7d82563b07a1ca49a3f509933f6018f55cc78a12dfaedb87a9ab009314b9a4df20e1d9eb5a9652a2e78241ac92282a7607fcbf22f6d7d4223e007b4a2ab9eb38df2ae73368d431893105c0c77cc3bf72d4e79db37397e4f4e50ac4a2f0da3124de84f931fbc1a29327db4cca721500991c10d2132132c341a6eb7e171ad23e26958bbfdfa0b9bb30f44a74ffa600aea6b4c82766add3c1ecff20b607c810143d6e14f325f0c9d49982b5489aab6290e66ce01f6e00bea4163d5bc1c74989e1247163931d6027835716b349f9088559329995959a183fe577192e66a3de156917ef4b70252452543704f2cac7da38d8e17b71e956934b82535cc1e8a0ab1870723720161ee2db9be998e0025798a9622e900f116735572193115e21be3938ca209e363723baffee06b4511aa421e5d617a33fd0ac7cd3ecf24257a0ddd8a516a4d5f428156203ac4dd7fa6ec9fd040caeaea534499a1965e7f3ca541961f64fb7297e37366890809e3b4a009f0d6b081f433ceeeb981c294633e3cd646376d33615c5837ae935309bdc6b67c9c0d8d391e87a674c0fb488a75c2c8427da82bbba6133fee1b0a2e490a83422d0249951eb99027c255cda2a4c656a246449dfffdffe2623eb95ab19602a05724b24c83652058bb2a329761b64078d29bbe018619c7d3c923a77f0065db9724d564bab2f13d43dcb354bcd49f97eb0594107197ef8b059513882a0a727edbf2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5217bc1f3ff728f2b6102d843192d4aab6d5f2cea0551079639ee88f140067cb0ee7c8d6e806208ddfa558178495d835a9083cd9bdbdd95321c3cb5bbc323df62a6dcf753ec5e4e68a7483f8b92aada0f6fb301d0c0136d233e6c0846d4c3825efc8d210168fdb1b473e0be59a603a3185c5585da44ef244b64c0e9d6aa459540d43695eecb1bd7f46e751cb7007b63ea9c9afce16a3b7e7f64dfc5ebd4d01004cb175d8cb425436d1f925628d65df380b1397bfd6b0486dddb9408419d25901861ee7be7557478255ba178039496171df7c9a7c222cb54ce09795d6f37feefd7a5f714edfd887b4efb7dcbeb0678a3c4905c08294e63ade11047bcba19975a1dcf45c133c738ff260c9efcad378138dab8fa7a4d124279830e814583e1a6ccd6b959e2c40fc25aa1a9a98ce7f83cc771eb496f64cfad9592818682b552b8e53a83811903804fc79840c958ab906428db9bd1e6172b0ba0bd06a4481a39e18d5ee281087c220b6f3587074b4e58a090ae34726324636fd8cc7a48d4211afac756b0bd9d09d58eaecfac813cbd27a9366e41105b65f5a934b2e883f8ce9136c6646f62f7da4f6bb6d3345c997704fd8314d2143379ad85ec785166636112006332d5f8d6ec58af1f91af2eed9311c386c1b5f5ae61a26a8d7f3101416ca2668084ebf8ba2fd4ea9831214ca58858df98b4a1ff115010dc83f7c2d9242ea6339a5ba77f9760d8a26f50af2442597e7668865ba178f96885fed4ae333f5d7cd08bee4237385265626b29043b6465dc02539b5eb341b9ed5a7cec96e85e2b1efa990ea093a860e5c13ac3c781ea4584c62e258d47d0d1dd9b8a538c041c0ff05a4c74c65a38d2c6fa231f591dc236f152b875ef5947782fc5880ba13edb74d7d8316223717ba9239f0deb6d8f9d8b859fc0d664984bca487f9206a6a1780cffe4317fad76030df72a2bcd950dabc20e9f720eccd48a5da414e9b9de471f4b261879606f8010678efb47170cb418762011c639b1096112760c895efab585adcbcc2c9e5a07646d4c365e6757a8ac795cbfcd2cccd1b48ae865c0658ba1c18a51d717f342c68301a0c1b214827fee3aba1b45918fbede8387304e48f9dc983c0d8272a16e3fd5897d2c123907c505d1b7c702b26a9db50d58d8b1948b7b7ba2362b8d470d79b2b8d4f876044c3b29b4588d9825650375e17f20e5884a845f9fc3662c05d8afb291364eb11dba68e7b288e3986f8137c01a57669eafacac04c8393a1a67e321d48d4095823e613bb01f95b87df82c971072772330fc287dfe380e9f62a77a1d2dfbb0e709639f2c28fdbdb340188e1450d4afc2375a90f9cd726da68bb5e9e5f417d61ee1a34d40699afad95e475a62e0f50f4a3e350859be44e4aa0a765413918e00287aa86bbd3b34e3c59d400c729ed9cd00d89779f4a1f9239526b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd11293293b2c30b670615570f1e9e34e0597b13f07a13ecd5cb1ab27c4c281afe76d60756196b9c382f314b606e3115e0dfba0b09d2b7909f8f361ad113830b22625c901dfa7c458ff226c62fe1be76b67b685615dec6f2e9f0e91b5c2279418b2f10321057005635eddd5e31106af45027afbafa7adbd19066992ff957b943614571033a3087dbe27652fc01729934a1a15d952f938a18103d2b9e0f3241897aa1a6f915360fa055b380cba844d68383c46604874410abb8162eddb05ba8f98ffd395bf0a336c8ba6eee9e3b61e08fe867fd5bd5b05c77cb0ff9cbe7fefc88940e41a0e23b15d55f140e8d82f3a013f1959bdbb2a72f34db88e9eb20d7b6afa77ea09d0ccc155773514b8e7bf832d969b0f4fb2645beba55924af88845910fcfc67b8bb0b68dc547effe2b815be450b418d3f66d874973dfb5ba7883e8177f19f285cd5c828bc809b03849a8bb513ac4291fc997dbcd11782d9e8a6582e39391fc65b164333fce13644cf5f3cdf530002042f50271d7bf719356f9dff44213ee03bf28d7deb0da8ace5f868ef188fa02dac63c066952b9b8a910bb6f76c67539ed9a79f4adb8abe434736a7fea08041247c94cb99481602125f4179f44d253349c0be6a9c1e806a6b74db2ef93c103bdcf9b304fee1e0ee965c9b881d35ed01b6e7671c23b851bada76039be8d7d374064dc922e288a918c76e7400fa92d3b1d15270279b502384aa4517d0d335a68bc4fa9589ffc769807205aec4da255b695756ca3ae3676906b644db0b5f0f9438688be19fb98a3894ee8a3e809310b54247dc59851ef1ae959d09a584e997ecef7119bc72d21a108caf6dea4be5841b4c29d392e6ce23baee8efc0d8ac98eca2fa9cde4715dd46e0dc60a6ca30e69e57601be0b901b58c404deca188851f521101b10ab1a5ccda46868b1c0a67e3cb057fcf4c62440d2c0373a8c5e2d499fbc66eb537893cb21c143c81ec92b2b7180ab54b0de985e1f56a96af983d32fe434d4d4cf613742cc4c38464f06f37debb548575d3a4552b5780ff8a72965abc171148029a4deac78fe44941bb415c92e7e42dbb2b91b139df429ed7ff131ea374b3e1813e0c84d5369d711849d4ae6a551fb2d4fff042df827695c09b65e3936edcda8aab3ff60a8db79f88e3c7b8a796127e0416b78c9bb852d5aa769a4815c8a50b071b8ad398df0a837048a414931a5cf00f31fe02d4bac18816b0ca0ec9720e9670e094031d5a8efa972b24508f476cd366ad2432120d930d5ea5b2b639e217d6265807d4b3f5633cad3dc6dc52fd9695a6de50157bfc783adbecf560eb89059089ab3957d55548e009391a9b2bf05b3e7bd9104bd006b2fa0b9a418a67edf8848478c51f812371aca13f3d236f5efa7bf01bd073739df6c67687bf317dd59270b36ede3e04d348d40cde6ebebf49b90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h51fa1b82520a1e290c36bda95f3662f3b75630256f4e1dd067fcf07837e279d8cf6dc5bb6179a033f2e19c81a79137f9ed0bdb8f0887d96c030eb85137d768cff92f3240fb406494446e448301e3b1277e5461152ddd44d86f085045dde9e0ec34025525392f19e6891f04a941c839c5651854e4a7fbe63beceab53320dc17f3a37f9d4a07451c30cb3fcde974aca30ccfcbab24ff8aeb20e4e893e520e2d0022f51b4f71932981baa85d0257204bf88132ec74f250e6995d2e77c90188d44f70d84945d69619aa5193862a62a209086cc267b57eca53946e9b1d83c843fa22721a9d737d4f5dc34732de78e887518ed6fef4f67d14e1e06ee5d95bc6e0392b73e986033f57d54907b4e55033978bdcdac4f57a27ef6d879857afef84aedb14c25a102fa27ab4850cbc68b928e558f60b7ee7d93e61c6db4fc23c4da859c32d4d85c845c2313f06f3b788fa901c85adb8b8bf4321c361e8afca5234fe49c39bc9f589f6bc258031cf0af1c018a1eca6f1b2504ba3a8a98eeeb71288cec465de26023bb5e20159d78eb88dfdc5042b5e544775605f767406f93a1ff3aa530d627682a5e96d79653282eba8e44e45bded3797c55ac4b8c127bf4c616bc5e3fcc0e62da423e5c88b1d56fb067f0208b237111df12b7bfaec0db8fe9e39988f5fec3201bc36157f93ba13adb1b26ada2d3031a3d7535fe6b5bccfda4bc181596c96d29e3b14cde95a8c095481c3fc5391e8328ce5e49f0aadf3d447c6ff155c1cd4b0f680bc31076f81fbbec87f5407f75225e84651a922a35adb79890114155839fed3be2a3d0c018f157d433fd66535230059f0735a58106dbb09424b4729698d6611617648eae94b5ae1d1da91cc0b00c6c2bfc88c955b5ce87adc931168cb5f3bb734f40c81bae23251865dbb6f49c19b7505361104f483ff24df40809b23ce572f0876504ba963039ebefb40bccbe4646fcb583dea4a2f972dcdd4e5873793bd707738f89de317b5d47644695d5823cbccf809f5d1dad89e89a5b0928d9e2e0298821d50d506f591acd8872dc2efb13da8ac718d650352f9afe4a5e420c847341ba7231d322576e5ed5b549fc8e41ba4e1038c8cfc35ea8cf882f66b2ed14f46a0af7ccc5e76ca510aad375d1825d0a46ad890533f4fae35256d69289b7b26258ded288154decbdf930e27811c7a93062081efbff7c3362f84a7d39da16c40811d968420c480df3e1a26c36e3308b195adec8b41b772aa5747b9b4b44088154a0be2a9d29dcb02f79f5642f2307d20c93d2a46ff7656bc95b258cab104f7d6e5f0389f84fbd1df4405c33263b0e6f458f87bb656bd742854575e206d838a9ab3005702b0eca6f54c583145a9809067e6e64f73980c299765a97c186c4741896018fbd89497f84204c010eef6f0d4f01e9cfcc38e97d261e8dfd7b87f67fdb27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heacdc5fc9d585df84897902faf22c9b7305219d954d1db61b490c3b03b4077edfed8adf8312bf766d0c4048f1c184124524ec4dd294d8293d29455ec58eacbfe0a8f77d74cc96700455f149775f929aebf044b307aafa2c3932d372c058959131de400456954c19defe02dc5e4a0dc07de8b6cfd9da93a9d696dd870b113a665c1ac5d125e9e2412421c0ce750d5d3621fd7ed5f85018db3c7e570ce6a94944b2e430e1056fdb1077a7cf016fe05959ee9928ec3ee70c4b6f18606d93ead0ce5e2f454aa42c11d2583b8ce3a77671539b2ca32d174d0bc35f922170b2f1e788af3c4452054faa75c7da978c1eca747aca509b58cdf73d9c7bb7820d28b7f97a73066f34bfb1be989154c8e536afaf9938d085661d0b68d11aaf63be54c48e2585092f511d43c5fdc0edfe7fd051d063cc2f046d72eb8614b88a4a0486b7a2c45fcb2520e75b7f1847c6da24487cd7cde55062388ad8ff3df1a63635e8a4e570eaa6fa679f8cf1331bcd191527a052fa5a8c96640f70a7be66173e703a182924f56830b02dc17abde878b5ea4d11736163e5d4b15996b70151857a1bdd4bb7aeb4ea402aa45a41eea164dab6d89ac010354de9c8026f394cd1b7285fa6b5c6351670edde5e4ac025cb2c88fe7c64fb69c3c8e6d4bdb46615eaef14417517f9b3eb04d772e5b63f39e885e7e09b69a376a13940c343b0ad636c5103ebe58eb5dc7dbadc2b79f8749b59e4855c723f21611adfa5bdc480d9ef523c406408dfff21a1ebcc1e5967908122ca9f2914e55d9e76deea329a580db3469bf227d4b573e9c4ae6a93858da712876b2ea2a9f566ef5a4ce167c9967179673208a61602ab154ddf0d07a033bfd1dfa3d222ccf9956c6e1789f2d6911773a8a727943a802b3802b1ce97ffc3bc4a56138e6aaafaa386459751907ad5027212e0d8e3370a66eb836a509d8582b121299ef5fd51e1413583ed2c8938f92419278ba35d7485637e18018dba1d1ffbd0ec039b052e85d4153ba6ef3a6e9623e5ef9eeda93899861326680654c4f5b9d4b13e5d73c8df1c49d7c09fc4be5d1a9fe88acd1b81a21c64758fd5db5ee072e7edc68f4820b51f536a8e73b7e577e9322c027f6730f98e64e8617fad1e2c91579a4c140b6e3000a263d43fbf3ab36e68457858c3b16a84f5d70c01b9ad8414dbd3925ee57f1a49221a38499ecd973fb7e80a15ec0bdf33955e88271b5ed54eabebf4845d244984bf0c7fee3f59f74334f98f1639f574f26ac8ea6bde2a43b2f485e3bdc2fa5a02722ca981c8efd85c5a2707a266c085b59604189307041031fbd7a1fdcdae52e45d4babf0d7271662a5171f6c62c577ab236929c42af54a73095470fcc13cff83468a5b0b5efe4b98fa31aafa2e13875dc1e788712f67d0d1f4be7a5826ce3cbfecca29620d339f90dd7cd95234f9c4a02cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hada42a070f0357005e09762ac9d9830472b20ea5cf79902daf6eedeb0e37153902e88fa3449e059ba5388a2da859a567b79c3b9563794d653c394be90e51124b2aad320a06ea0cc6be3042a044454b524d7832bf6f19372c562ebea37305515d15d82a0dae6e519d87a2604e1c7097bdf1b5087ec3518f5eb61ac75d1c85874572436ab03dc02f9b29dbf12f598f2cb274812c6b249af7492da7dc070f5f1c650e89a800de72edcdeb133f56e54cf1411256ae3247baa46d5cf69c70a1fb88aba8b94e49249a75936fb22f4ffb547484eb12110ad31e3ea846f78ad9724171d48ae84302e562c10b9b10780460d5d38d7c20d76dae2caba51323cd92de3ba79c9e2ce36924a4f3ef349de7a7c1cdc5865825e0b44f99cccf77bd50ad576deae893220de8c52abc7d6d89d865560f0f187eb4119540427ee1b91e8344f77964b69d149c00ef2bfb473570c4f82a8be43751358968f395fbac6c539783eb23006d2725f0ba97cfdb85d30f270e3b389fb3378e2540b4b3b4f29540eac6f12c4f6e143633e3f0e84ca0e95d6e5b99a7778eefb75bc1474300aeb60af8ac5ef86ab8eccceae0798caab4b93cd1dfada9609764ef6acb015bf1c16e76393446bd662dcc4c78dc89c7d2840e15ce93c98c6e7ac9d311aa7efcf8825f96dc4d05555bbb15e1bc2ea4631319efdf23115c32c2446d9621865f30989f06363ae5412892f805436f8b3f2a3bac6c135feb0a60b055dd5d5876b239e8d908847e9647c1e5e254da6944fcae35c328bb7657a35b126da1d68a53a32d07ce598818b9febe72afe3a86f2d04928047c04ba5f310a6f7d4d62cf597d607623c6acd37dc0a2590d083d4db5a16e53cb41a313b5e52f42b101f013e4344f36afe7be916fa0c58c70cef5ca8a45c12950ff2ab34c145a5b6cb5c81bf54ff44d2960a278a0fa37da83cf3360f7f69c03e15c78e38fbfd394351223535cda569c7856407dd3e93591ad3e5548082b330d34e7a9693e71ba59c8df38de0890faa7c0478039a5c731e97c7a8981a27c60bdb0a1343e30cbf9622061a3f3f482d6ce830305d33ed979e3ac171b137030257c3b989137403d6a478ff4eea909437847707458eca2ff5c7a0a75eb48ae518807f4358363402692df1a91249b585f591591d8dad542e6964e719e163374a6ef295db6eadec0a3f9ca2bab10a6f690455a766991ede0ac3347610197c6782cb0bc7c177e02dab197dcfa7a90a3898d087edfaf773876e6d22c58d77983b03d7841193333094e264dcdad3b8798181a854ee61a5decf58b01724da911f47e06567b3f5f1c58a28c91cfa83502edccfdaf4050f8057bf2a9ccc10ea47749973e148cc3cf4a7c445003337ded25dce5479536aca66336d065b671fc141704899fb5b6212636053bb3d8e1c8497deb2533c3d1e569abc57d89e105629;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0fac186d63e4016e8d4caa7491a92591eb81d78dc7cf3055bb1a54617bed96e6e56b6319835bc3fd53b24a5d075b66f4df5216672d36c8e66ca5fcc914767dccf6adf45b49dc2a668e67ac5267969164f4c0c6f0e700ee2b433201adf48e4d50422129d8e0bc766034f7fdaaf876355f28637df9499b64a46f8e969ab1a36af98fc2bbd895fdee57c1c7e2384889f5194494064a130f1f22fd9e87f5dbdb8fd31fdb37284c9ed5759f1d468df67852824e532bedfb275eb3179ce6fc02a120f04785244f98b1c0eeaeb379b2a0ceefc3c76c46904920aca0d6b912f3992a74f328aa33786fdca8f0452080f6f88cf599f834b37d10eb439a56c405544483baabec7f8532debad5eb11f72f6715203614171aa83e26ef2079eb460ad1c7d0bd9f5fcee27c93bb028ea87e4acb0d19ec13fd446b62d8fc65da6ce332dd3291cd21a02dae6d45e424faf53f1bd729506c60f114f9f297962d6ff00dd098ac0238040bdc598583a220be8733de4af0fc60e04250e76cfafa3f3014a310ad84aeb0cbcac93cf1359494ee69922e9d481815ce3ae813fd1823edc944d9e5e044e60ab62ca75a4d275a97231d5a119a923f17a097b4a2167cf759b343faea132b370ed3bbee9826a1ccb4ace4f4ac93f34b761f48f23171f3b45b247282a55401e242c51003f6596cbb5765e74cf0598332b5bb3f9ec9fea11488617c1ddd85d1aa37275f1873d976df81d659a52be101d267dde73c82593f1c3126b45ad4906812ebfd269110c621691dd7fbda5de1d60b02d56f8b713f5fb033700c37029aadc16b0c95ee39ceb06e64d62035c319b58f99340de0825105cec2729e3f216a1ff315d721537a16b0cf45f3d96e3435cfa55fb5476fe6a7d3c609e6952d12c28955afff03d363c143b84e4e3532aa17e82f520ea5a961f1af8d4c61fced06812b0b4f8ccc323370f159e6919d561c23c91874bbb06a8124dac5e499852de393522bc9c7421f2d3e34211f9ca782ba22db7b66e1849153fe4ab5d24870b035926f7d6240f41fa8fe1d39ad5f4651ca5ed5e0fee577dbcc88fd5ea8c889296774f1873eb1b9acef96f8b51142a55349aafa9c90f866ffa8f090d6deee15bec1f7afa9abe06b91e01ffd2056e3307b8a8a265eca7c050a46396d7a040dc147d3c7e2cf129e427672f2ef075b4d9b5de2dae490734793011c112775c6134f0be8f5f531750dee354c97213992c3613971d9a67e5b5b1a60c9af40bd99529b8894f321e5940ad7caa648965bfb61fd41b11f2a2a2a193f18c3f5f8e6f7b2f6ce057c8b14881b525cdb90e6f1276d969c3efcf93210ef53f58687fa164bad3c3a315ba226af9f12367fda13c5257bc3ca9e31f68ba3f2e6b9f663a2496cbd992b9c2a88f42fc075100c0ed6120785355d7037e73f7f2dfc7d80d2a11e47ffaa905bbad1602b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h77697698645709e069ec2027deabc004096ab3960a9f7faf11d8019883a58d9470104586cbad656f7de2c6c9d06c0b8ac38e61de0e5bbf07ce28ebc96ffd1de301317cabf5f22e3d78889a5ee0134423ddda6bfe5d9d6ff0ab5bfc236344e360baa5af9fe196fab4d95e365fbe0d769b6b311bdfc3161235fbc7a2765d9de084359e255e85d30cab1cf7c21148f9889cb2e9a712a63b24120a136ae9fba6db1739cd2a0eb8db4bb87e00d520499db5e16ebae6abe18daf0b450b0659cd414a93968dc12b255ed71ef5c112ed1c7563bbd8fbef15ce672fc1280d11129ea694a2b54eae23643f40dfc1c2345a66e035a3825843f296e9924c01d4dea8b09aa95e8207984a78b7aca467b1913f0e99d23b06206dc7d2a24e2b9d2ec1179d9eb7ed21b939c27ebe794bba0990444bb916f1e5f2ab6ad91578a257cb2e1358fecc15914f0174a9de6eb600645c8a8938e48c48eddec25860d31991f149aba01ffaa356c121d5e611f7015f03e308a5d91c968b30ea2f8a67cda2a1a5948d3bb2e4a86b8ca910596589c3b6d77cf8905a67bac08fd02dfac774432f1cee41c87f7712539411434865d7799aa92c73edf49c5ff90701bac02b3bb4579ac8b8163eca5ce01f25bbcadf7d7601505ae14b799302de3f7760dba7fbf95eea31acc639a13fcc5fcde7fcfc51ea81183880adf3480e50e579218d78e93490818335a997bb0519e45b63da75cdec486626b681b1681a01748c93eb54153de315fbb55a0e751e38f97201ddb4229d97945f746c9b82a775ffb440f7a7ca05bc9e85e302965761b6b1f2866a6ff466b281228a47aa8aebc164b9a1a9c99004318a1ac37b8f17c23703d3f058c638bf52ccb9c8a9d067d47cdd341fdb59c9bc2c11e54276edaece776188ee4c23846ce9e860d180ab570f19b3c8e185541b35e5cca2452bce2e3f9a9d1948de4701c95e84595db6d8a701633a9eba9060adb8f9ab4f0353f2433c971878bc30e7d11b31ab3601e54d72cb115c0046a94faf7068288ac70b804136f1248df0e1293e4a3d7c51b88597dce6b56506c077e39640616882834d10f34356821cd425732024c72389456d65c710d18f13bbeccdfff057699c480342721e50bd3b2a81843d85db980a1951af929f8f854ef914f969240cad5d1f635d7f64b57f7014308e2beb0bee3ecabee0c92f1b339c86826e6d62633bef9dbe1a57fbe5908cce7483ce79eb87d4b20f7897b2f238c3b41e00a4e1d02ffa2f06bb5b027029b1c729238e0615eb51f360cd5090b62a94333b47b23d50a9a85fb2ddd0fbcddb047a4294c525ca58b5c25d7ec4fe8c13b99f09917a6f7be6a0742bc19ac1261f4e4ffc5478dc377ce8bcd050192db08096b42149ff25570fcd62f9765c62f9ac95f95282531e3f38338fbfa8073ea0733527add3b64aedd6186fc88a2f3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3984cf33c8056e52f4b15f7f2d8d4fd8a6305350f5b399a39cdca210e968084100cc3f6f79817d6717f9b004d54b11af28e56e572956290cc8cd7a572778d2cc82ff2fcaeda405f6c15c4a8e8dff977023f0a544c20cecd299bbf0d5bb80c73e7231a54a3462c6bbc9a43739afd2ca4cbe077144ffacdc8dce67eb65abdddef8b9cf747657a6d4ee02b6f24b458ed6aca09e9c89a73ec249d12a6e19fcab5772e3efdeb6fc586af6cbe35b0a607b0e2a5523fa633aee5cd6e490ecb0565e8bc77584547edc982adde93b35404fef6286eaadedb6bae09a824a8bf1519ca4975c0191e937627a60bb03a944d71151f41703370fc575f6ebdeedf1b2e60bcca8341b7e018cbeaa2cecd2b8be120bec3995b964395f2c81c472ac4dc04cc4644dd135bccbb298f6b2717a0f7f8ecaf2a5af8a70cd516d69aefe80368157cc8c0cb360054925de44811291148164668f4573ad6d5edfa633cf95ee64c3546f5d8b423cb6fc5e6a87707a09f333dcdd93f4e3fe01e1f4556dffe253cd059c23f3232fcb470ded020c9544563fe850ded344e5ebc23d7830fa4882ec15c76dceed84076a31d96d3c1667783141c1fe8086f9a0054f3ccc18754019b09a6526590a582a71936503996259f3548f670170ad9d71c2b27086d8ad9b63e57346aa5f6586a46306306f8f98ac6429d33ccc39b88694bc401bb6ff3bdcb5be2d0fc939548add9cb0debcb81ef1069fdb89bd15b5cc526754378dce31898180399bacf242a7fdbf05dcb0d198e5679ae29dec5c2b41a9ad71a666dd0f4e7023a36bccb45c5dacf3e121b75487aa2f2eb40819fe256ba7faa08cd820fa004e1b3fe9065587c728e431e26f1dcac3e65ae702d3ef6d939693655fa859ac82facbdffd8f1285d747d4d0c4322b279fc467b0761d9359385e4d3c8f29690fa66d31f135dadad5eba4bf72587f7ea83766eb733a8c2890bb2dcc89b03363a1ee43cae3ca81900a0b4a36144e20054b7ad52235f594664b182d5406b20c3d2d6f52bf7f3591729acd90fe71ff1be1168394c5f6d6b6a3a805a7b46f229f5506a9390664f5ee80d4ce9d9881de24b2754ebc8d7a6dce8f77a9623479a3a9112341017d7512fd76f2a37ff8f21545faff02a3a2c0430b1aa800fc0003dbf41f2cff3322a773d81d758016e5feed6499233551893a124c4f2c1f8892810c8ecc21664d880139a8ceb08622fc8f7047c6d33be6efb7aca711635264e486bb647f02aa5ef8c7a8bb8f0380d96b76b831d556d41edaba0cf6f9791a58af83569d084378cd47341003b9fe5c8c236f9b1f1e8af9d3766f364baf244d24e6ca502366dd4e883677cba0ea75b9e52e144fd95ebc55c2141336a0c34951246dc53aac8260e441c807326737ef9932a28c8f802c344c19633ed980425499b5ef2c0b5a5f8d2f60522fcf9d628f99ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6ba585f04b04e744c0da7d63c19a14645358acf1663b9fec4ceb458c391b852f1936212aad9bea29b848ed3ec585223e3621111092e1b241f85cb9e8ea2b3881a933702ed1ef2e0a4dbb9b09a406d87a68c20994973373034574a734710eaaea54eb8041fef2b83423513c7c797c59b00468cdaf4097b3ee00dc98ac73922ca1557c20b36551398d324df9e46006ce92ba7c418608fd6af806a31334cebabd1c967250dd9b2e012675b895d05ffe02f797ca8e18c7f715dbdfa2a304aec0c8bbce82ee4c741b9ae32dbb022cf546b352170341c9d906fa0a327ab2c346bfe943db0c36a36d5bfaf5ad5156f7fb1ecedfcf5fb14e4db0fd1da1ec3ae52c969418d70b3ebd344cdf6137cfe2bd6e73576eadabd72822a4c5041af0f47461ea6bd2eebcf80c8d6e6c4980194e0f3c7049ed520c4217529bbc45e3021a97ad04e73648cb61a9755d3506aadb792186b91967ecbc10609f219ff2469ef3d9c09e7aa7100867d725248c0ad57732b277b31d8d9100da280cf87f0f52ab38ca7ce13bbb509a2c17e73a75f30d293e1ca16bec24782543fbe792a23d4a0e779c211a94e6c48e2a92b31ce1f405faefcd586644a1fd44d6ae2fa9f793060fd6d861b948b986bb783660b47fa66893ebf612bbb058771c36ad8a8fcd7b5caa48c8b38b83ecaf5c2848f4f01dc1225c39c5749ef851eb18f420006de82ba8f7e1d82a54839608bd6335e8ab177d6c1ef8d733ca4ee3d0906ea1b03b91c340907c50b9413e6701804bb55304fc1975393c0e5cfd607202a9d2bc078c61eb3f7857d3411a58f9b089dd1f4615109b40283b6faac3b59550d6634c3459708e9c997711ff0ee6c0cf8f23d587ff6041bb7e537191e8388f0cf9cf528bcc81b5c087d30aaae5561eb6d93637bdfd61025174e55472404548f9b5755745b26e6d5c10174e298abb6888e0a3b4573b949c311ff23c7cc78b4a4ff410d45c001a456e75dc3bc069bd4eeb8c096afa2f5387e5b190ccefd39ea969ba8fe91cb9c72cb7bedf8791225f88915f8068c7a6206b78d254eda9a3210447a0a95b6f645a00232aa6dde3d8f274cda3ff3b3f4c8a3cd83adfb23559aef3cadd6f9bc81495f699c2ecf90655ac7440ec345dac2c5e86f5d95cc322198b4aaf453c0cbdeab9f77ebf40ad6feefe3cc6e91040920d8effe3b0d2a889a685f2e50a1b58e723bdcabd135e7ff65901489c53b7fc15b2db1ebdf04fcf886170644130d5146adf21ad6a36c6dfb7842f47e0d2e3d4c2778ddbbad8e0807d476817a0a133cb9d848c540422c6d4c88d7da4b1a48a11044ae24adaf504637ccc4f9560bc1aa24f5014e00dbb0600586028aa4b1eb9ddb4ee92b46947ead6a7f50e2a4d056ab3f0d824e149a2891e59495147c17ea04e666cc300c2782499bce400ff764427a1a2e3689ed7d8348f2f1964c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h902591243dfc8f6c391daeb2d9a2fdf4e824be39bf2e05d3fa332bada643f5f32110d83ffe0fd4c136ed6ec97a0f1d8352477b5c88b0d6cc996eb729f792cb5f27386493e1c7ccd21d9827f80aef537d44938840a4ce8aabecc6aca223c4088f854a25c8355cda4eb914a2a59d0ee8771309aa55b7f4fd1543402c58add254ec569b88aa6ed2c724af9572165b0fba8f73d4010da1eb1a80f67db96f52ef90cc33bbd7fad51754f77cdd0f829d9b24ee6234d838e50f7cb43329668784cc2ff3b269eaf52e5f4150f65e6b09e9b580e8ccc1fbd6dd773f05e7ead78c28980f5462a22ede76607a6db7b3bed8594913c129bbb793e23849aad093ec459db677350ec50553b54efed56a6ce76f70ce1c663dfde1e0e68e2dddfc25521ee30bf8a0cdb5fad69982afcf5e7a996f5201046ca1306041067c14f83d4db5597600a9eeba09b0b57511d4bc32fcc2abb0eac83ae0401f1daf3305215d78dfa17828253226df73b9dd01fcc133e4c1c13fc85d36c71cb8578188c642521a09521fc24578fd57906749ae9f611b6149ff52bf97cf4962d815adbf40468378d59c74f21af0629f7805484ab1377492a5be6ad099acdfa58417303f5b5d7d701f90f430b0765618ac17bc02fc0c7a1e554d680bca4e8cddc12c15d29391cc621607406256a581e98fbb92cf80fca29c263ff0d6f8e68c484c0addf7275fc131224ba9e916cfde0acc8bbafd249f0fac16ec6e85b75687c689d1a93d9374d74fe319d944eb85e541748677acd6e0d4acd3b9ed0029216708a813105890ef11b35164cc0e488061a8a07073c4d545a8b290619e2c527cc4448bd27092f35948a519980afb655d0378186a76dcd30cce858630e4807aeef795ba41143c938781da61f46ab36c7307cb72b5bb61b6c16aee1cdfed5fd5ddffec21757d20769f36e91951face41b8f5e1c73542d30b3bb506dc24cc38629e4347c5c7be4d1204f439197e549229ff69730039246b6e0e6ff6a307f9c7e0d84dc07b1b5f080deeddda599f5e4e66b5bc872a12b64ad2a9db7377c6284d73638e746fc80969adba0ad354651cfd2e485f82f92baca6e145027b71a014609638a7c12eb78c101823dc27640b42600a194517be22867a2fc97decf59a8334c18435e1022f5cd8428a2632e5d9699e90ef3a1b1add44f2121a744ff2ba6f58c5685be0fd7c73f9be3a8756800ae7f785f1ab8967dc359feec3998af8ff4fecefae7258961e23b11d5545f433cd6552ee3d44b16152ad3fe3108692b9382791cb822cbc3af5f395766d94a02bc79c67d43c0ab19925ae09aa8e90cad0c410fb87a881c6dc01276adf5694771bca62d1503897ed66479fecce74a1c3ed1895d6101c79916a66c12272926db95260283e9cabc74ea0e717731b100360038aac61d3c44e1271ccc2115ddb8b37bd48f5724e42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbf5d737a0baff2ca3d676b7dbb7870bf34eaae95833669e09b68578c38271362caa94c5174e04eaf60cdabb9a84b08fbf033caa3c1a4bc37b068166495c31405a6f91aab7a413e2ffc3e1c4786f4fc4b974f9d254dce6673aaac8c71e60cc76a4e476284f9829b10fcf11ee359233c6b3eee2f5093468c04939d424ddbc0c2ec1d83adf706806316d3db7b84bc4ccad4e17b353323719eb79c4e8e3b50cd3286a4e39ee4f5e5546540325526cc0696a8ff725cd8eedee13f2a50144f85de911f24eee111d7d9b2e29f5c445f83eb8561ea44f1d7a87aa5db2d29f04e11269ab48353cf7a2f2ec3b475c7e687350a975e5dd8a4babb6896f95a6c1feb864b48438188838f18c0e2873f4c0019f4f1ec96bf62affb3e5a169c41099ba180acaa05ce3a815d10e55a76521decf0aa5965236bb7a29e5f7a2d0fa1b03d205979cda792a370e639c20a094116f4d370dab66049a432299438ee1524c80ecb11f7298f017fc29ecf562bfae6239c2920cb1a24d271b8cf91dcfc03a7a3d254004c012e7586d4ed6cb33338a93be935336b5fd99dc0c6d016b6d088398569c37e98bc91f6e2508f68a47067b5cd25307b1f1f7dbb75acd6589b66769e014ed8f476455ef20ca271cb8ed50afd9b1c9a9f0f9ed021e0a23a27c3e0dd6b4c7e6d5b87cf52b07b9a17873c45ef892e117eae3d0bc9ee6ad9516cfe84a5672fdf3b038158c5857073efec5a49be974f05bc00acbdfcc30fdb72e705ca1e97700b58ef4b90abf71ecbc8ffddeaaaabec811aa68ea4ce70268866afd654c100fd0b0195014f84812339b015c0b0efa35bc64c24cff17815deebdf803fd074e26c4bda42ce9351b7fe37bfe28b4a0ffd84548bc6f2622f418501ba7c62d63a75d1345f89ab531b5f9d9176a3a285f0d830163f6d4d44d91f4b14ea065806fbacb777ef8101b71ec3d42513835ca16a2b9200d12352fd79c50f8d8587c7c0214bb197a842ab1364cbfe9835d45ab0daa8fc7384b9e10e071fe59b6e896679ee0de082f52e19637b39f8ccb0201280489a23072627745bbb191b11d2905c3ef64b9310c2e95a6c80fe1bd2a8db52e83c9eef78fdb6662ece991b554a6b2eb0b5505d1c7806eefb3a0a9703e45ebed4dceee57cf58131b3a84ef8e53c6d43a360ac4f0c24f3b01d245fd3b9451ee3787a78d560409baab7ddfc2f4a7a130758ad8290958c4d940b58fd7e9afa08be1b1d68fcd0bf65e26c833b4d49b5c327988ae09b36530232140147820eee0ab129abf6af99add89e95a3f82eff4c5186bf31d5eda6db195a8d7fd1d3283cb6dca5c7722dd42df65ec417a90c0e9b2fd643284bb5b7a4abad3fa3c1dc9f656d4082ce3bf94c07e75d5f1a621745b0e1ed8829d15bf4645a3b236815dece7df33e84e7bb458c2877a7dca14ae56c2c12cbebceee73179db65a0838;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf6a9173ca4d2b9694b960f7b3bec827c6c0a22c89ebd7aaed4001fb18ef12f26b22ff07faaf3cabe326ab16e1748d6c793b7f33ce3400f80764ee63ad139200d2cdc4da56df37a7d15f1498b8abe4b6a6d5b023ffe1c224fafb3f87ce6c850179638fe614fd74cb12c6043e9927a2accc81da739c72c9361cd16e3ac5021a0c94f567da47f429d656dc4dcd480aeb68e12105ac38a45ab12bb761f5bc8dcf1f278fa03d7fecfcfe3c7e8a3f5d913d1a87e9dae2a66acba3b50863d4a955f21fc5a2ae4ddf9ad456ecf3796d022e3c14d581bb09171152ca54fc3733564b0bca0b591d47b0727a517a11df483746c85c4488f70cd33d942cc2fb10e301185f76b7049dca9cf26589e5493aafd53c6238939a478a389f633fbd282e0e8f2265048cb0aa315c3df1259440bfc014d5a74d088188312e69522e22b5c1f020b11686b18490b04ac12d12d1519fb253102235d96761ce7f283345234626609a3b5a3404682fee020f48660c42251bce058388d3884ff73777cb490d34138ef2d24ccfb569bd40c893b4f5d4527ce994302a4584829ccd8d79c9df77b84d7fc570ba74db965a7ec9023f1025263306d78580aa6ca486c565376bf5d39f6a45cc2a3396ef46ace004ebb88933307621adcb0b3fb05d6aa75fdac4bac6ea535962447b93fdccabdbedda0edc856deab72a03500288999f97c2ea007eda78f9b50f5ad320d524d64973b05fa0e2004d173e09ce8a67a850252b2591e183c3bdfc6829d0309abfbcda379ef8724d4c3b11dd6573a607ae4bbed2706f038f2988a2730dae65f5c8cbb5de76b0df9b7297ac3be4976ffb1f02e5d140db8793bf875cdc96a56b43c10722902bbe4ad8974f70f0caa9f08925c63d3b0eb0477c3c55a32b6d59e9d8bdfe43e3e6b257488c308f15310908634e360527ce79398da302005434b1cec5a91fdbe5c75afbc9d1e696818eeb1f907a42c1a2d8b6e6a47b37664576f5f978d07ca19e73d91f0c4db349314e77bc717152c4b5ab60a4eb4dd120736386d4c55cfd92c17f3f39271a7f3ca4ae0246165244da1b05b54771e49d150e048a187ac3f6626b4378dbc54d4826b709bf96278e2980d4cdd30caae1630acd31abc30282e088492674118f50deb3e79c7a19878259df63331b4f1368223f0e60daf0fb63922c2f2ec6d56aa0e62641b21615301fa3a02457f71e1425e04ea01e0bd5e998af54358f653e4594ed28cb921cc18f28043d22dcf85fb5ea0a1be15fcbfa85e744d9d4a0962a69ed7893cd14fdd9a882ec8bf5060766593de47bcf6ec5981e3d40d7f3e94c73eba1ba1bb87c61d1476fb860e06bd50ae23178ce81d2e60ebaf45756c035eeaf0aa9d243c4d464e79c4dd1f06b436e67cad1295fb48499290fe7174338abf8a80a016900b54e7cf9c26a34a455aae3af4a5154e86326af758;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcf5b41f97f7a38886a638f63e54e58e8db4894f173993bc719ff643ef12db06f17e770aee26be5f44ab0ffc43cae284872e899a4b78fd11effdfe4defb7bde3ceda737d8af01e46925768d7ce12b8d49272c5d2ef5a1c3947cccb598ea1985ffcde0e766c5204cb48e858af473d32347595240d457a49a87bfdbad9bff10449608e65335aa1135453256bb85af9d4adff261aebf6e54629956b1c809a977088d4814932664d254833ba54c8c1d87b1f0c7daecc3037fa5c95b7b9a85734118ea863884d2ebc0ad9ae7077550570dfeb6a6c1b4f8bad7faed997f90c8e99bee3f7fd0e37a3c381758412ee257981d86ceee65fae935eb354e5b4552b405feda97cafc7d931074af6da91e7e96b6a75252a7dc15703b5a7a127b05e537b58742d3902e0953465de87faf51b5c3d10e6bd37151d5789dcbf00612f1be3f30be8bcb02a5594897b224cd7d7002835b86580068fc07c463f19c0b5ca1868d6607e7689f2c352d3d26bb44e2704959c281acbc93ed8b9c152a6b2b44c2d5c9c908ab7a658c935470a7f367674a24bde25498a2488706c85619c6a7934021c99407161ce9636a7dd8a3f2218b209cdfddd2cb58520ea0cbb3e7ce99c39f65e27162eb4e59b99c1f2f410fe58cc68962ae3c5d206e6a27fcb4d2a66836cfe825751eb57cfe5f2c07ceba19580e2825b26febb55a14d415f1cfa0a9a0bedc47445e48aa204712cf2ac23cc40e0d2643b0b641b47cef6ed384cc6c54c0edbdd28727d512f6cf78aa6cf9ed6c31572e758f9eb9311f6f7f586a430d4d5e4e98ed363630605da8463b82baec5e26ce0974f8a86cd4ad675eb40a39754133df65edd7459f7215b727e958b30f567e8777cdb865b8e57a301c72d0c38c1797954d72e8d76daa93c03fc6eede360a729b97134153202bc88f0421d15d7d495953f9684f2b3ce19d1adc5afb4b8333ac0ec19a682f11a80a79a7801def93146b3f5fdbd42bc750fe9202292b1ee94774ca95178ff4bda355d43bd6312190d3cf9c41ddf1b834b1ca25feb8ec220a2b745d767ab370af7ddde352a56685d64f921f9008e31c655c183a35b7b98677a91ec801e9dfc0c56892f584247a457acd282f4904211fab54eee877608bfec7887c3ad498727a18e8a8e5cb02f401183fd29e00e1c670a7f55ac7de741598837dc7c8be10d5315cc51898450330220e72d5e66ffa3b47ab84dc23ab8e8f73b4d63307df08f79ccc15c563a916051bc7f68578082727e6093101afebf5d38e8833e857bb8a7270ed8e9d07a48ea6f6c95d2a8e18aa7918a204d55773441969ea2f900b6c9b7f684844e6586671a8fee5d60faac7bcdd193ac600dc6b85c525d66f0e375e917133e4372aa10a3272897cad043b8bd7aafcff807d614a03de0d92c1cf73a2e4619db54bb4ec2a4bdb0d2587020783b8bde0c50297;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf8bb0a1cf62936c328dd120ed248517dd5c0c300aa542d18f42a824a7fb13bc2dc9f21b2cd6b925015f0d3d319a8e4f179e061771b7e88627fce10ae9ef32281a2fae0c1c6f303d1df0fe76e21570a6e48acff2af320a4d309078c3a3ce67e55ddf09b3b185ea80cf714f5629f5b0d0fbac2835bc051ed5c95e59154b6d3425c8c4ef2f1433068617f6ac0a274dae165836791beaad62e33b63ca12a52da9183235652e342ee59e641fa6575b70aa5d39306827e657b7d2a98226278273bf7133a6c16a88bfddb520387e3f0e34ae56ed5952f0d07a078676c00b390baec7ab754c02f0a73292577c7d8b8a5e49fe1db94553f58f7afa9ea9d23df3356dc34f0f680931589bd8a5257958c3750a0f99e2321e2778c622303c40925978354958afca9b07cecbf0bfcd812773a45df30eea979813de72cb2e23b4ea96b6713f212c91a6343ccff7d20eb3cdba390b3ecd29a4110025bd53c8d9fc8da04916a87d81552f70cdc2860fe3f94d8e7f88f2ba0fd884fac529f3efd1b515a6b402a93db66de0c8434e4272e02c0adeafdd9a58598907014a8b0a7a857aa161bb5c01bed4f3b079f3f4bf7705beeab120a4f9510f66b499133eadfb0eb453061676de7f2d9b5b997a4ce5d3a4d1cfd2e6ea13b2cbed286014f51f283feba4af7662576ae97f31ed1fb8f7563e4f6c51f3ae03fa53ebf0ac9f775e8bc737c48236ad4ca14ef0fb6ef299a7ea9ff58f27e34a39e2aa15f100890f89ba76d172f2a3090b194767e76918caccf8348236ecc46df58605cab7a65141271cf56844ad5c7b420ab61da3df0b7407558939b07bfea4e6d5810ec51663ec2dae5ee6b4345150768348cdf696a10b7644ddd6debce7439f0c2af449058f956a62fc1271814abbdd2a4ad69d40b4d721051afdbf63d92372cfe2ab7e48cb9a4e5aad8f71434e09eda8621864998d8855e74e2bd239b095a2259d5402abe7f408ca3e74810796a1779b1ce62f3fda93578678d45feb8836da59586df25884424eb284c4b285824d93199153cf7c980d85823c2563701e264fa06c79230eb5129b263f2baa288eba158a898d88a1467fdc67e04956f40a9ad2bb15296f1b6afe11c68e96d0490a36db02dfa0171d3bc34f9fa3460e7071e4dce93ddf87a32841e49ae8e87f168ab90338510a47cbdeb070f268641e008132a66644da6d05c6d68c4f6c1aedf1d47faa0fd3d5bbc1457a51d5c51a3f3fec2e8ad3480d03218f173df8a63da37831a33dc4c6420d75d99dc82b7b598be9ef01e89af1622c970d5083312319991014cd9d6354229c6701aa7487eeeeb84bd9d5e411cf26c0834c1757e0957f5980c53549ef6e58037b3c70e08a29b257d7e6f4fbb9556758b213af849c169be07e2353e6c94e88de8cac1bb87d929440570ed831393c4b58192dde895fc38e88a6072982ab4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc9c6ed12b60b29dd1f05580f70616b0d304ba029a8ddb9f45d405d990b1ad383bbc839908097dcf7ca1dc602b7ea1b989b8e1fbfc79c7095c9605c94d6e18826c06e8f586ed56e93526f4ed99b195b006828a87035ee7ca86cc35231457c76775f16bb3832f460cb0b519e15ee4005396ce90991e9291cdbe3c38bda88b410b754fb33c0fa0200271371454de104a68c49fe457867e1c2eb6a718b9bdb4394742211201c71611244acf3b90ac379586b11696e50217c1759758e7b5f2215c50a59c488662112382b1a38742bd0af4f00af6433d4b60b7a7565f53ff398d08d2799f9405aeb99a227a5bd70e44024f26715a570e2a33a2a835000b0cc4bdb6d288ad7fe83ea950c37afd8c31feba2a532e22925c85dd048546af9467ced813b2bcfffb6a8ac30462d4fc07e2566d7b481814ddd1100fc64dcdb4136d1a3152678d797f84749d9a9894732132dce0a0ede2bf166ed882c1b6120d0969f2cb55add2892f0ccdc5d34d22b11f80b2de4c2fa3a56a9013e60a13554f5c91f683c9b382c26e811c3d9afe3ab944823526d4ef11b2c3324cb687f31b1f363045b8ddce0a15594890368a893aa4106e804dfa52549d3e523567e3ac94609647cdfdf32169bfdf7e007a4bcc5c0b857743415356051ccf12088202b44aa75381672817d33dddc74397b5bc723e87456ed7d0019f1085c3cdd9d18540cb14afe529ff4a73bff6ade920a8c9f2fcffc14687bdf8a95018d0c6f5223908ff6a760d110d728c658b14de195a7db07b8fed51599634c9d6e5478b0eeb96ccaeecec32c10675c387d69d69f8ddfaa1df854f63a8cec2939ba66e26b8acb550d0e5ea3cf19822a894762932ce43e8675d8d3cbe0a97dd9f7311d27ff6ba92f8b491b4181ce3aea52d5d1eddca0936f0cc434694cfea76fc27ad0e5da79fbf32f413aed399e7b17da8fc94a105e9ffcfc65bdee92b3842c9697368522b7b0edd581a86c6a1a0c032274cf426bd48d01ee35515ff0b87578f9da8938ff8541ca69e719c54f2ceab5adbf299ee4156fbd51fee6329ce69131117119a7726681b1d1ede39b79e1f9670215ea65e79bb71acca0015881be2173dd229cf61431675ad4af76da4898f3c640e90d9e1d897d3a4340b662bb29c67a8ad333a5a4952557ad711f68a3c072de9a3b0c0ffcc4987ee590e3189948ef5e78e3840604b7aff6073aa739db8ee37bb3592cdda6b496ca5618470fdccf72dcd8175de7fbd6c3a6a13e0639de5b8398534efc3d11e289f52bb58b5fae291ae95c1cda1de235d6b9f9538b9a8fb3fe2f9e82d707d6c02f48552be4dc0fdf0e300fe63552147f6c9383eb71e1766f240a6ecb8c6c8d899066b117ba8112d30b03ece3cd656cae8296f2f05b17274426d973fbc1731fe16f11e50db3f0e273c302692120e8ca1076a0d4923def36a2d056f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0a46d73b78a819fc9266db16a565e99ca7cdabe2e02645ffb1220c6bf8c2683d8eef3c9ed2931b16796873fcf6faf90c005a445a9701b56739d221a14704bbf5f008b092f854336e731a7f04a7e319309fdb370d195740154782782d00ecc45a8b88b3402f3c10f3fb3a48a12f724dfcf8fd728fb9e896d525e3adf2a95c99d12fc71d45fabc70c78d0eb2c36c1ed306e5d8853dddcd69788889b2ca6ec8a87fdd9d41952208b45218afac472eb18ef16a3c354aa407c04dc710fb9927d4c3db12226b7b815f2ada89454ba3ee320ca7beb373dee4be29f5adb02b2b9059d67c54e4dfa5eab9847d5365ef611565e781986342167723e954f8704d802469d0892a550417ecadd6ac5609ac5ca79b0ff6eb32b3e24fb1d2e2751672260d3b9f7d2cbf3d4119ea1f78966ddc458348481007aaa216483b265803c0fde19958204050b5dfa1086ecd00ea4ba84670d10a5661990888c9106454bcc55f383a17b29da7190dfb5f840b5f2db6d8fa57cf87b4547c326611be21e27c37146ea727ba8defa360aa6714f621efb6e0c9dad61012e9b94571da583eeb514658c05d9b5c4f1e082320a6050de9a48e39154262d821a235ada9b966b5aec2f0ca7262f672b0d4685db72e79e566962ab29a11b4346eb2ec600f1f28d39949a38531bca5f4bc991d7831a5b7866fa521b41aca78730a9ce91b3dc2ddd362041e8edce196a4dc531e1a01591c5b61e6b8aeddc59bc1df4ee16b3caf7cdecff8497d715da9a285c70651b7b3c2012b7b8be942820d46a9a19c56383f89f86c24dbc7cffbb575d64150e9c0b9ab96766c4e36b6640b747421192d88366d228bdb62f57499762c419a8134bd24b1cbac72b8e601f3a6edfdb742bb6c03207fd129f1e128b9c0153f97acb8f9b1084d1a35f74463b5642236a4518b89fd271da5dba26f3335d9db16051d00ca5bc81d41d7839eeff8bcb7a77dc5fae54d80ee91c1c6f281fd05d87865de2f8f2c2fdcc3c323b88fe82f47f9223381f8d37054d5d7a5f6b09e4419ff19a2161b144a27f45c94811b8a6be20b4f683e249a4a0ae69958ff6f7dca5d73ce981e83c6a1d337504c18beb888c67a703d3196c64ed21806b3eb90336636c48f77b649cc40c23aed38099264ec28f9e94e12b75c8d4314ee530ef8a8bd64b11c03f25bb07e93f782a8b2586ab0a2e27749bc250fea310a41aa600535d9aa925631bfeef9d38306edc20f814a476017ee5285d8b4a2c1329aa5575d59e428e7a92c3b3a2e6171fa4a60a1b2a3eb3b9fc81ef4c4f254e2cbbdad187d093c6419da607c22ee471b04d6a03a0992366d1db67a787aec76b3882929d709b68775ed3f9736517f046cf26ee9c2b0d920d5d8a1e7d2efdd41410a6cd506098c1bc9860a483d0ecc980af69e19e980acab8240e36b480dcedae85c21364e104d3bbab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd6c4e8c248031417decb3a9a18190a86634ad9c98c77327d15e3ccd2c5966a40cf8ab210473fedc612d05cad13a5cfc444b9844237d9e733876c744056a0f4ff78d6a9978ad0ca56830249a9157be08cd18333c8e5cd65dec61edb9cf99b145be17ad1fd236bcb50a9ee85d68e7b848bf2ac897b5ea4109537066f35bcb32056ee5b8425a17f4bdf8b79b4561128e70dee6f7481b95fe0489d24335e42eb53e4bb7da8ed0d114f2d1ae120e5401bc51ac8c7eaf1e862e81e97557bd23a62ce93f53dea72f451d4148c50652fe192d8a031ac1f0bca961e297d9196fab5cf76663fc948aa69a41c88d6b220e928bfbb55d65a219ed794897fb19b5a4232d3fa7753e8d76136deee06c0632ab74631de609e2d5af8909f03c8f39a9cd19fcca63a6dbc08e42fdcbb1458a6c1671919caf96541f8ed9b4aff6fd58f4b19ba9dc2a1e48af9746e173e75ca40ec450d6d4450fa26e3e88bc76946cc807620f5d13438a334b8e4ee5af94c9e5ffbb4b9e34b132783665f612ec2ffde74987f9fc90d93edca3d54971cb759b58caebe317d43cc58926b186aec048211f31b73da5622b14fc86ade174342b3a6b85632473e3a51a0ac22441aee7b5a98b37c8862588a5ecd76da24c35c7b99569fd41df59b2de0a486a1cb879bce0467af55ea3872919af59e795d33b90b8113e3a14de138d361f18e9d83b6488cb2616d470d8f7e00a58635533cf843a8c30f47bc32b72a808a2e33a8778ee1c5d319e4ce0ada6a67569027188214c9621d0cbed57461844dba2b0b2d93094198b788ab8d92fbedcaaedf3796a0778f3bd5c4933348e375585426811a800375f82c969ea8ae180ac14646ad7c9d5ca26879914be6e8d9c25c0aea657b52b1df6d76ff1f60d6b770b8263449de2d4ae34adde1bae45acfd0713c96e50302443b6ba3fc48e1bc01965139a7bb98431ae537cd03474d173f892ac54844658d6291f0527e32c239528a59f87af76b5248f74c9ac4a9bb1d2761d2e9c605cc9415f99b67ed4d29daa0cc03a53573a3170e1dd990845b393ca4bd4b82525816e8b6414ec748ab52c11d48f531acc841d6fac1c1022938a2daed52d5d22ca243f50842291bbbdf9e7c3ff97702471aa6f11efffb18f1681faa4bb66530af7a7ecfa87ddfa680fc5a88e1ef0f347f642210a04234813e02a341ef61a35b6879e28e4191c4c122bf3893291a90bd21b8a41e2f6757a238151b200cb5d65dab1f1e8147a6ee4f055155547db9c2a6c04b4965ba2868148e344bef9b078b9156acc98c621e2e063334d221f49371b43a8187303720a85d459aa926b6461f712514b49fb7a8f5562474b21f594e2dd44cd27d7768329d198dd455a31ebf8705df918f9a2dbe74511d0861b3f426805735c91338b07c010f596a9d6ce9b9571c1b9c48b68192247d24625e40ec3d8a1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f0803b77f98736bffe3f26eb160cb020f4ffebc4ae475633ea58b5991be198d316511b9b71e8e6240b090ddf48a63802884f40fe5275d8611ef0579b28b1552a48bb80c4261ab53f9ff7c65b53ae6eb7194f45dd1470aa1651bdb298f41ce88de56501ea9a6729b46c3040c8fc9060861c1493a237b3e07da4c8188453c5514d1407ea037534629eb4ed86c82ae73b180bac317109e020caad14effb460c88d8792100415fa193f8a19efb2413b7dddbf53c15ee273d6b516d52d059bd9c04709db5b09e71241df7f0b18730d1b1edcdc8f6b1291ad923a1e706665ec983e3874a4c14752070804ed28a820474e54c75320e860233fa7649786774a38c79f33d1f9b291c25428803f46e8295be883b8ad488c68c28a4d1e6144f9e96ed8fd401c3113fecb98c459b0b16225b33960063e099baa99020cd5718a22741e621f0f65eb84c8345f6ca1ae8622d9ca92a3bf9c820c135eee32f443597173100227cf0ce12a052bb73b9d70f247e740606d3f2d3ae46d8212c09c1b8a5056365c0a9f7c29ef016d07bd2271572259f6ce1c6d43730a898cfb5a8660cac45af507a7ce4b781e81d58d1136f6de2d2b1dffe68350834b63c1bc4ffed09734ae902420dda877a5e84e93797db9600b19efbd1d27ed1100fd6a69e1d5807f26241c81ce45556171fe6a81276d20792b02792b36d1a70c0106e5ceca7265b004f1c119cc1a56cde9ae71b9458a1b492c5be9149f57ce71dfe267295bcf9394546950f3280e18f5373041f545b504c1ef8d1008339a633301f24069d995eaa21bf2f8b0a89d41618634c4bdd1c03a335a1ee2a2102a431c067bf04bc25a9b886ee8b6a5e4b29236e406feca7707c628b8f022a49fc84d91687fd65f9a6c280b0578c5a6b0d2a5bb7020743414c2ae9be118f010ee0f5dd6c8314c1d8d2b993a352ed1e5ba862ff801f20d4e35ff0460c85b920dab33e1152bae6d4e81e6e0aab0ecebe6f68eba5c8ea7a2cabdb9aae6239a2c7da0bd45b36711e181a89c9f44c4a669055ecddb872494748c599eb2a3f2b25cfe882f2f324741058804e4fd50171ced277d2da250ee55947838788306a54e1c4fa60aa2c125bf0384be6c57b1318163a6ff18efeb07f8b6197af7a40d82ec297e8abd63673e24bbfcd3d2112e3a21088ad9d40aeded46931b093552a90ebe07e0bda9a70c3d4e0d7407a8b5f7e59c073e9a253bbdb1dfbcbdb747b68778451ed4f735c17011e02b503351e8332cdd6920129a6dfa3215455db1d7d2eb02a25f232ec10bd59cebaee98749fe6f3a9dabae7ad71821371408850cb27c5eadf8889d51f693322280a4d03e5c82cda03bfb4b12732228bd34ead4633c67b95a2dc61ca1fcb9d212415de760acb500a2c1d28244c2a179779b97c42ff1ca8b48334c389b92401378a75038824ecfc335a4cf706360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had8c3c39a29c82e73cc44f226a58c467137ea64fcd21c5ebed33f13f5f1ae5d39b0df231cba5649e2f6cc8977ff0c2a601865253ba27b51b9b54c21f0d4544892197d58eb084d275126d3eb6c04661543ce9dbe045219800a1649586d8d3980f8a18b8e0aaa1bd1ea6df35a622b2bb820a7a738d60d2d9239e5e704f9b6522d994232f540f7ae963d2510957fba8010229ae939bd086a9c6c4d6c365b4e4392c3082e45dea2a4deb667033fd72af099a3aa06daeae944e80f5304489888aa3770580d8f1839696cf5a9f2f8e86b3e021ff65fc411a818bb2ddd8bab9a74fbae31f94b7dabf5c0eb63272edf1a68689df9901f81e440ecb13d36bd278d7e2459cc022ddb3cfc19d9f22577b83d1b7c434f6dd6b143c0b19deee64154fde78022a83416451dde3424ed6c8abd5f13584d2bcec00effc9ef2c41271792108335b9a099b8c9d275a06283c58e2d9aaef28dc9f0bc7fbccdcf76bff24f52d78ecad2d46f73ed6a5bf066f402ab55ec542c7ab51c4be199b7dad48bcad38478509fa83b4e6680e744830e8d442996f08c80acfefaf9a8e3e85c84aa4cfd5175063215126498944fb04a255196cb0e559e7446a47f441a9472cdfe01b19b63c90b684123e1c91c52a849c0763b5740deb58023cae956cb1974dddc915d19a617240b4d6e4b08d6a4aa6b7100d8c9717d831f88c7bb62f7b3c9b8e5cc0a3ea8ad5473299a0933a68e624c94b7312c6ca3ef1cea4fd30c0ef008eced3bd7e12f38321192cb8aabf035a16a81bd2fa866e8c2bca76fca000a91ed21679943f3120fb9201022f4fa6be19635a2ccfd46800dd54d1f79c7e541fd7dbe9100c41d95d9be936d719b76264ad97ad71308dfce9a12b4dbc3c474f82e03f5094277f2bba004c7386c3e9938dcfc8283f139800d4259e6a44e03844e83a690d7513365459f624182c064d790225b3b26a8549029bf88a1b938cc8ea6a07535e318df360621e56c492b07074383a17bdaf7c7ba1ff7ec509dc58f56023f7ab5db6313c83dcf38b4461c8edaa8f429c9ad306796ea2d520ea360580f3805016d2d310a06dd9dce198d3799f7e8f32100ca52a6462bb081930389f4f24c08aa3f55e4f03339e4171c83478d2313a84e7d06295aefdf895a6b765f8a5c9cf70511cdfc42ac92ff810a19aee1566b31a1ea05c6427a7094371de7c12a5b3aceaacd31f5e37ee193aba5b5abf9ba35a3fd104d85d0dcc4ef03aae9014d90f3ff0b32e016c473f772a85edb29ac008dfdcac83012d1a70c3eaf601f668a7783da748cbf9e1938d3ee5fb9db507a559425a26fe207c896069670adfd4a51ec2e579d7c21072e8bcd1dec60b76c046f7fe3591f5e0be6baef0956424b1760ecfadd02ce8536d27ea7d4316db3c7d4bc65d1f869aa8ac2ebec23abe847f3d6e9819dda7c2e9448efe6be755a68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8aec06f8ecea2f0b71890ef02a3efcaa851ac7e1d59fd97a999cb8416202e26f32fdf3ef91f9f7ab2886d21ec2415d7f5dc17ea68f47e7637da377623c5b9e38acffe7cba40530eb9d6b1c063bdd55273e2dedc988c437829a25a5dd5d69bc7ef836b3f5382cce9b740760ae5d0442e639a68d2da48daac89879c53b8a2fc857d57a1eaa2f0f55e1f76b066e125a289f9bc9d5c4a88b9aa8f34654c9be72743733f474cc4b1de09d1080557ccc0bbc24178367e4b9a7784d8ddae5b93798634ddb73246e5030ca7d88378e18898c59d255d7b8bbf67501690774c1c19bd4a6bc5ccf688defc7da72565bbd0baea58ad9620136947e28ff9754835305ce21c671f8059aded2467f57e0e75503e13c180db2edcb876d5e9d3788e086d7767404ce08a120cdc5cf95825f140f138ac82c7d73a929c54e89c88edf4232bacece861db82c6c36c16952d602fc32b4fbbb2771b2e775721cc1e99b0df696c9a417da1078da0100d4227c2a0beeb77a825848091fd65a4afa7ef4ef079065f6f20ac0b79d944acfe84c017331f6528445c3e801c624c36383616fb4670b175862b806b09e0d7c8b4820867776966d4a8f1d2f8dbe510c5680777421aa61d95a8901988dd6481a361384f1790d5db95bf6c78eadd91d1f8da3a9ed28bd8794e6c305380dd2630ef6f3b287344d6dfc27e50f149b1bfd9c93bf8d054abc7deb293237db8defc2bc16fb5b32afc65d635079243cd58d7d943339f28c5aae2d7ef72e53344b3c4c6bf843e8a839804b65b1b54803689a753671f3c4c9dc86241603179124ff64d295a2c5490cdad8fab87030817761486eeb0a9996478e939b57c4101bcfd98e2f33262372262db18ab3e51c81339607dc016b2e0deb6711796454dd2c648327546302615d802e77fc9f2e0e64f4b4efb8d13470510a2dfc2517dcd119428c62950ee01a29c4220de3411181e3be44c7239d137fb575748d562557d6975ef0c86091ea94a1fddc6b709807b6a24b67cb0b17ddecc0199fb4335c1c8bad35ac206d5232450f5e46a31dcdca2021acd5ac7ef639e577ebff3d644b91bc9cba4cb65cd9d8ef77e55e64f9ddc2574a74e4258407175bf949ee01b0a0267070e55ec3ab955beb25c0d7c46137c724bb9b08567f276f33fce41a4b4335d66514d6edb9b46fa68a4508c5f9caad65e7403206c3f4a321bcecd7f21efb70415b9f66f55ca724d2a6db92a4d4f682d87b756b131f7d82c3521000d1c9b96f57fb2699136dda112625857cf62dc5813be98887994a49aae4c4ceae6041c77fa66c8b5ef9246171e2b208ddaa017a74c9485dc0c73d791e33b72fd3b6b77a4dda68c7b3439adf222f22450da6969dac0c676e3ae4f2fa4b0144d61b57d4d0ad76558f81a79ff30fd6504e290f6ae197a84f63ef976c968d9198e931dae5b0b18bc04658e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7348ea1a195a894c034d99e6b86d2b8a37278db032500edebc517d84f9d9464fbdd1f543a37a8f5cc82995a3272331f4e08e746ae746e89ff1c37266161db1c4216fbb49e44c7bb21c1192f341337bd9f29a809db55aa340cd3be77f16ecc18989bb1fc7281d4e51a20f17be849b5b80ea0349ca47eb129a52c1b0ba7e5c66e7c25a94195f50e9e58a450ffe5eb7a18b26b2636dc66013a97db37eaf5a145631f3f282669c7aec9bb240b0998afc57f18fd4a97d2f74aee797eb5cf4af5181f7472733626feca1a574f45e51ce62ea945f2de78de739ee7aae961b960ba6645f167ce8e47b504a181c43128460a592fe1e1cb5715f7667a2e7d7add949ddb4528a63b426224a6e1fcb1109e6079089c7303ecfd0cd8262fc14344489857dabc6c9f720ff8df5a8104c30fff708afccca40b2250ba26b1c47b1f67523f4890d5ce556460158462ad2a7d9250fd754c7867722df4af06fd4fded4365502e5e6802faa5f9f66a82ded1f991f487e9f28a1af9026b91428c21ea1f899205a5246f617ac7853fdfa29431f3ee2636b0302e31d0b3cfde6298cac61933264f88b4089f6f3cab5515e20a051240a8d11f6cfd648281f3d7eed82228aed2880b1e496d000e4a78a04288e7183cdc4f0657c243d98ceb46f76f4d3bffdedd0ffb0418c6a7da1f6a2841931370f641c62e0d91e63503229570c47fb7b8093b24781ba2074290b97237380dc88d404f6d0232cbe5c62fa91a83753732eb1fcc28196f278dfcf872c8c08152ba383bd5d699dd107ab8fd5f2bcb24da30f8ac1737d7ddd767d435786eb2d448fdda77ea246ef7b6d20392c682cc4712c75a9118c7211ea1274793c1cd91963194283ee2c10ef145b728e553314cb8347d372b9b2f53d59631ff491b16d08f4177d045b606273e085193c94ebe40f9e663148d889991f3622ad86080bf2c0c49d12b8a5e979cd06a488678ba4fbe3a1a5fe0effe03c9d890deb5a61f14019d99f46f0f24a66f4f488150a1048d3879a20222e98ad021207814904d12b9cc95f793ed5afbc4f0aa2a908e5f09ac02189041d7cc0b324f08b359755338584e384e52978fac2fff7d226a3b19bab77ed6c87900fd0faa4f8507b0acbf01b8bcac867a7c59d84fc3ea7e871637eac8b9c912a99ab4361074a841316ea191e30d8e05b297117860f4e7298c2f704ba3e6deaa121ead79b8afd99474eb164c8fe236f880954abeebbf14eda9bd14e39a9d41afe86923bbddd2dedbdbf8ee89876033ebb0237ff3c6a7ee1cb81b8ebd52522998f1d2bfc1bd66b183b5edcf7c8788fdfc6c3bd66f1ebce09dc31afe918659fd28ecd3b19fc68f8436792e10ba58a35a923a27d87355b221d9dd61fd059d1e697222e1d26613c179412f8c51e1105f374382e8331b92bb70839f96ed2fdc7dc85b3c217cfb021b4c55eb1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3bf3308f47e9fb78f168c99fd56ffb8bd09e620f6b025e6482d9cacfeb8a4ddc24a06c51681babdb45a0d1bef79a4d4e1ece53502f3a415ac5ce15f41a822e5bea26b8c0370d26eebd55cb917765d89046d524fb29306baf14bca2ffc4337302f4cc7c7deb8e263c6dbb1821ea8ab79c35376f70a4e6ff89b7a2c0bd18513878928eae407f90b4792924ab343971ba948c505a094f473d4f9293337393744ede221ac71a543edc227ec3369f72f84ce625d44c5b45847e688fc5f271e7975e0ab089a5eeb848204b4abb2238b087829c5e34e6895a8152f366a836d59b87235a093b9a2f92390a4bb97803b8472f7d806442a107b72dcdcf140c63921490ecf1843e6825f3435c3efb7e94f482042fc9bcec9f821a7fc6cfad52b7696eb5f22eb5de7ca0287983d899cc83d1c2dfc59043e7af35ba61c2344032f5899f20ba85d38fb65e08f0c954158c12193876924e4ff7cc4f22d7b17d2d934e4ddb42adee12a9fab6651dd335055e9f80c427dfee71a5a583de1fd2449ad7709848c1d1c582fc76afa067a770a5b6e566f9281ff30711c06a8f65850b2fb7bc4dc01287874754910ac8b0cfbb76a194067edcee57d975f60ac1e4d7fc6a85ae92194a6856b853c8ce0386306e42f2201a1f04fe0fd6fc94b465d6af4584b831055ec1127a5f9733263fe65db4e2bb9b52b8454aecf9b59b1ec5fb9d9441e5569f3a075caebdd6f7c6df83d196543666c6ab4b5efefd44f009882f51e5e256f450eff597d6eae18b482a6eac858f40de8cbfebaaf17972e66d5c17ff1fd18f55ff5dc153d99e98946700c6dee2c6f18940d1f3a2233a9ac21001fc8de39b460a2715a81b12c99f6818d5c758d1cb971fba027aaf1e9c46f6f8b35bf4a58058126d70cfbfd44b8a6e542056ba4f8f10973a47256413521ef49950e5adbb81a6570a23aff6db78d44dfd380c8a2ecc38bbd34d25338459501fa932fdd26d59011db5391f31087fb4b705948ba452d70d8f58ee63c08e5927ca83d02fcab99d3dc2537ea434424d6e3351740f55bb688bf7c564c6a489c3a550fb3caba58cef54033493869c8e2ad7de1231aabd333eb9cde351f7491a1ef1eb8ae75fd7e62b3d3ba617ebdce63ae1c1646f281e77dda49a712334e87ae822df457a4d5ce496aec300b85f5c0301a52cca5f25209c0e23d20ba76f6e0fac23658a6de00ade2ae73bca7226de002fc1a4dcff5f8d36713f84258da8077a7e1ea7743f641c37c82e2024ee6319c1c494a51582dfe9dea6567a6547c25dd4e0915bc79974caf7ede75e320bcf9f5ef08fa481ff809c5ef47eae44a5ab0b3bf284c43679196bf60e68f785178978ed6eb3fb8686f7e7d6485feeda9255ee81d0d125cb17fe4abb6a5de5ad5b794ca5e9f036750c8445f64e3b067f444bcd860485ea401a7dcfffda4b4450d5891bfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ce4ec05a0edc183039c18b8abb08dce3f5b0d46ca062e601985bd0a902bb7ac0a667b0c5e2dd8d777976979e4b36ead7930e9c1331a88081962998c65c6d3c14dc1a9194b7f2b356cd1031f593eecc0a9f80e13797f08ef0e8f134ad26fd26c883fadf667c72a1b24432ac56342eb521bbbd90f12220d5ea968e97f160aa1bbcbc11aee37c18a77ef559f67590b428741d277abd9e7f6368b489b963fe36db5a6613fc374e5723f3c7f0b3ab4cf4a4630436ac4bb31463d401bafa9093b160e1e60380d1833e5e483668d7db0ee3cb7a689c25ab57ca16a4be13ba7ed54de040d97d9911d1e6a965b78ee3c0b9d1ca49bf4fd6fbb7fef748bd2ee391f152a422cf526ecefaf3a4ab13ca97c2d97bcacdc51c0a23f92dc8307b5e2b6d6b146db662617044dccb7d07effc7dfa84358b5e88c5c83b82bff5134716b50a68b87f8c7fb0be7d457224427abb484360d2272b9389ded9ba288987cfb9cf48590c331670faba6b09eddac59e897fdfc667c971e320cf6609dedfed2379958ed6648a563fa5859e33c9287bec50da8f507f280b5f6b0837bd6846cdc55033cc62ca3f3198dd890d938c87af1297386504fc084501800f82b34a888245f50b0d2da2b54d5206dd7a8669d9470164c1d03a795092dab49861ccf60865f9fca838b312c303727aff451b3a0b3e639502e67d6756ba089969ac6957e47cbfed09a700bdd743cb46c3afcc43d5a7cb2d15d97c82e31f9d037e4bee03eeb7daef0507b62ab7874bf01cfc9b6c1edcec6699c20238b8960028e9c3cbb946c1c0327b16c7ead22c765b57c3904d089c01b0d4da292f24ac781751f3a35224c7393e67a9c1f36ea4cc0db20502b5aceb9ab58e4abc7850b2885d97da8dac2e92522735b03eca861ba0dfd98dad186479abdf04c632b48b660115fd0535924be38f201b7ea4d7c55b5537230340f03de4d243ff7baed09118eb0bfb987b718d23307b12b65db46f07d74aaf4d945d8b81c093204e7107aee5bcbcc7f11de57302409ea532d9f6e47a5f3efbc719a3c2ae08c354ce0c1dbefb5ca1a9a317e219c82abfc4e229c0c3c9db739f48e3dcf6b331f3336b6c05d76eba0da2317a8e7fa29d2bb7623f0332121aa8d52a28e0fb83602b7700ce51d03613856e5e9b49ccb191f41d3ab7720553e4bea446c125309f10ebb5917b5931fa7eeb0c808e46bdb66c455e4b5cac3afdab9e364656b3cbbf89f5dc6c08dbf651dd4afac5e7197234099ab2e7835e3bc47aaf00051c31d49dfcf9c662f902313204cc23b84a20f75a05d48d8a0793309678634d37144aa5d412db3a899b6dda9e5b603ad71879a981e98d286a84ac5f94b4defaaefeade5946ffa03fd571b48934ecae221f8c4a56d50baf54d2c4fe67b59452f0ea244c3f07fbd4a554568fd20e7f4757b65c25def4266a73a8f6761a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfbace3f67893f78f6e632cea8227b04e641be2436dc066acb22429ee67b239e8a1072719f3d3606eff2a4f1e66fbf5bdea9c85b42a92c16a724c5d1ff43a8341abbef487a2c256bc171ac18648da5b8404823db9ce6b2c0617396506c8ef234ed956b9bea7f3fdb192b746a1403e47807e7d5988bfbf73fcf71c78f7c8ebdcb3fff12b8082e45d7d176d62d1b534b3f5b66bd6bda8e166e0cb7e7a550235c1a534accb953e508e60e8a3907f214952e7dc94d88038bfd6a7ae31ec57415a1d42ae7a461e071dba0211c53fae14b57da974f29a240c579cd00861bb3bd7153a0b7343c54fa2f7c35d3719c62e4370c28c202a33fabbb97fd78ac89305f87a18dba8ad6ee7a990af232696ec6764f3c20176357e24d948dea16db8a6e7475fb4b18a9fe72b2cae9f7a6ce7e96453dc9e33afca0e7e20d83cc594ef75d9e3f5b430364cce76e882905639af8d7cd6e12a096da0243b2ab726040ec045601e7c7d97771fbaf8a41f2bee3252b8f231af14433cb64a3a105a4210754738aa12d7f2eae3465e74abefedd1016a162606d157a084a0bd052652d87de06ed5979d7ff3cc473c2035a08401b59d6f6f95ca8b1535015ef241a6a980c7b18fa0416a7e5bfa5add84506298e320fac5ebdb5eb32570415b5e519ac71e37b3b95b13aded28ede9b26eeea13da9fa450ba33b7f62581bbbad76ae26034ae8a8722f0ee712e61e7ccd14142e2a70912cb9cbc1558df14093c5bdeaccede788edaa66c9391454aea297a5d3d04ae2daba5f51903367cb36e7c6a239759858f3800c0088c92f7d31b00f05bb9c47edfc9469ce16719d922b643521a257e780109aae256ce69ba6e4f2c4d3c154aaf2df0599ad5031b1286e552946020a6d27c051f947af88d3611ac29cef9c78e836e1134b0422aafc844d25d0f9a3b85a9bafe44eb8189cbcaab323057678d91206c88f77976e66c50c84cce5f506505fa6cd6589617ad4bd4b31977b40a986492475932f29d0ad4cf6c107d7a316f5cb4c9962df3ffb5873e3797e77ddba9fb9be8dc8a5eab7bd33c485cd9d297a7f033fb63d729d7f8ad0c9eb97e71ae435a2b772d70fb4ab09d476d34915596b56db38327b0889641cb81d6eaa1373fc6f35445d281faa5ba281a55daac0b7c36c0de6faf5625f776e5769b85d34641cecde6edd67f625a008a61f44f062a05190db26ff617fcc3106c87460b88b52788682baf2c2ea2e09f570f0153544c2bc40fa5a7d6f0544ac2ebbb070e614d1f56aafc5b4c7988a0851987c505c4f1bab566b80d0d25f5896603e2c85855f7087f0f05ee2c6595cadae4a0f191830386d6685d30b4b4ad7c61388745eb0ac3b35e4dfbe3d7860530ba69628bc429426db55e26c03135acc6624b00c40a99c6e83b3b719046daebf9f3e72fc1ea2c2e7a0039e503b24d3e8cb0fb98970;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbd4ff2326cb87bf6577618646686e0b1029171ef7e3fb3c109626d883cffa1abd562d8bd7db0673f801be35b1cbf76214e76257e9493812b4964fa1f50d694ead7c47647195660306eca811e2706c78404e05d85b2c9658bd280c0e0b14e321df2f68c64d97199ae2cd4d861f17a4c12425338977dacb90f96cc0d635427f8cd7b2d9e91ccdb97874f5c448bcbc193a853edf09bc9ee9ee6f3d9f33d5aef33b50e1818823b2bcdd92ae84dd1fd1b0613833ffb523a55bac7a33d3a5b520909083021a12140da94fd31340e327d713f827cbe3dbe8fb78338ec72ea63c448c488a329fc46a2586abbc9a50f8979fb1e1698c4f2a2c9e7346d911a64228a79f0ff3f89e876ecf8ee010b02120df7ed459a29722e029a30965a7e1a7e9a26d162b441858008e0cfb0f8f6aeed15a09abc3978ed05a02c18fe69f53e75af8b1fb11cf0de0ad34097cd090c01b5be38240e0ef1f4bead22b1b05134492815476cd92dfd5e7cb6fd6f1ba55a693517adc4689efb03158c69bc57f7ea513fd28c10a7721449dc7492e2d53a749dd0985c63d02185ddf57e52e5c40b8e3069c5e0ff67b63ac05776a68aab2aa869991e9bb46fe4bc52d725a39dfcdd156d43e08b6ef1a421e49ed9fcf0be3595b1d6300ab375a6b0bfda8a6573d6ac9742ed4e96a8a953d331ba996a04dfe9740583ae000ac6a1c3a2597ec4601e57f6549665b5a26d8ad6d0b66e17aa78ad80576aba97ce5f8e3e4e3907aebe0671a92320427f97d0c406204e1b2e182306710cf91c6ec9a28b097e0ae950b63c419d0a8e8f629b9105ebd59e2ac4d29bcaba5d820654a84667664ba89ee3319ea6f0d03a9dd65f399a76e228ad230c8ffc6858c71ef94be54e4d44a88c0f823669b19eba7719e3e74bb585baa2b1ad64e79b8d1b7e1d1033fda06d2a15fe39fa94a2d5333d3b22f0a776e51577e96f0f5c3316fe3cf1581763ad2e45794fc583839aae468b6540c56e75b41495208d33c9d91e778a09a912072399bbc0486a887c11062764d9c805e997bf55e448bd4f190b14d98e10ee24ee612a05b7d6b869aad3654994e0f7b1a72b976f38f15c5a7169653df142c2c5b0c1128ee4f7a43bd4943aa524ff47f981c3b320e825c0dfe4f7bf9848113587e4057003b8351456456a40518227c144108f317195629f9e8bad0f4ec4de6c481a42eadfad784574d1720cf9fffa53be482d82982bc67bd1ab84c8e4918c8fc43bb165c2c140adf2b63fce754ac1841c3af597cca1f90b97ee16369854a6129a78e598e6473c648dde0d110abeb20499cde26538970c43ba27fd6d0e78055bebe812c2228808191ecc213360af6ad5534ec9a2f0225776316952ad018c793a5fbeddc21b6d8d1d1fa376ff8f5a9e95b9ed6219a7990356573e1c951b5dd479edb7c0bde36009d49a2773f642aa070a1584;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hde1bead32e5473922bb21a75ba419c2a3382d1123f80ba1e04408b3df94d71489184ffc11e92de1606825f7bd1e88ee05e3272ef169bb0bab517f7a52baf423e87401efd65667359b7cca4d63e1cbc0af5ed4394b5abdd33ff4eb57ae17a3d224766c7fad6771bfa3f2448c053169a5990d983841cd3c0cb2788afc69af6f29327aba51ed42168fe8a4aaeecaeb9f1188677bd7a7b7bbad56957b648bc9f6a13223dd4101658f724c53a51e08343f912c10362a359136c60c9a232acdf09c8f666338c6cf96d04fb1c7192d1fd9c242e5ebcf3363b0ed4baa9468019f61cde3bc88a36eb2021c6db4615d416affcc39ae43def24f8b7486a4c4b18d64cb6ddaea1ce6d0b92a0042cdd4999083691a5dc577bf856735377cb6c4ab784dd4f5aa68f5750a392b9d7ce9bb7aa050a35b316c9a1bb0c28ba658d88ccc9d5021fe6894800acc08dc202fc5fa93727b9ff111cb62f6a70f96ea37f3d3a4816297a7b9612b78dd29c094cb1099eb4960d8c43ccbe27c802fdb6ba19a04dbdbc6c1e5a51ece4ff458ab2bdcb99e605c2350d31f8580915c54900a5fae99a3b318a2a11085ed0b7bce86baddcbef3076a51171005576e80eec0ed0056ab0a9b00be3f709f09a5c861dd27e82b7b33f7e62f07b638237d9ce2571383d1293740f74f62ecc4a20a4e68176dfbce05b144c4f03ca39ad4a6571a80cd73f1388494278c4cab79501d648a0d4b4479077a3d2caf31894d6a78019249a8ca1bc7254a8919b2111e51a9f0967ebda3f2b09afcee7068bca31e541ecf79d723de235606c20928429e70ae569ec4b900043166b7d2c74f880d1aad3b78d08869309edc5443e677d146f9daabdbca6391be19300310b38861d1e7287469d1df1b2a042bdb195dbadf9302ce76f7cd3c03ee5ee8c38e1e73ce24a78be1fec8807c41c0c6a28ad3b0f0a13cabffb458dba65e81c385074d67eaedc8919c252a008625348b33000e631a62cee1e4e6700816f7bee30d193e48fe7d85217c587c0d0620d669a10f51d91bbb0a96cde19721240d8d38f0c9c7b064e10c8c2b0ea3ae803474c6bfe368cdccdb2ccbd332a95e3460b36f6fd15a5ecc64dd3432a89c9d839766cfe28a335f144922d609158f8b1cfbb54f77c68950cf0663d3888195202ed4a28c64552aa30ac6db735017567dc61da027a9cd7210376f710c86e074b688b96b7481b6f90a2b6a5d67b739be83da4f3e1736155b8fc5acc9cde20e18ef49c97d02caed98af623b4b11a3fbbf7f8aab02ae3a15dba10d204c0111d386e8255c6babcb007ccae20484653849bac15f982a83b7a9202c9d1a3d6b426ead47faff374f452311085b9583458613b1c29d01e59920f86fb497ee40cd8682d96272c5fa28b86a8ff31270a2737452cfb16c72b5e0164e21c6bd3df8bb4085b245e44889ef1aa71cef94c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4bac9b8d46290b9b785d7cb9db55946be7ed8815f5391ebddf979184351f36656909eef36f168e2b9da20edc4e2fcf3017b4bbae56d35b6d7443eb687ad5454b70b72e0ceb540b364afacc506c5d0bf9d2ddfb0e0cb0be9906c5318f5ea2421fd9f970f0993370380e8303aaf4a0eb9804f5c470647724579b29368894bf1e401f7aaa5f62919e7cc166dd5ec8b6bd4b60eceff021fc67051bdcb936df487840fc33a4be47a989a2e15ceac4136d8df0ab4d1be1a134a56efbbad0e8c3c72b234cdbdb29f583a25828a4430489a345752e1bb9883f9765a3f87f1a117d1fbf0fcec7a443df2972bd936849b704f2d45383a0faeea3c8d5a876d0bdd3447242a249c8f75b79e9d7d0fc410280d02c382c8b62da80b75829cfeb0ad077b4d11a77691a51e8fb0fa135535e210b66e6ace5f99a8fd6cb3ac285ab17cdf4594a039e7d7450d7087021fd5af8fe5b3f9d8848cdf90e47e56eebe7759b47525c6c7a638b5f68b0d7ebfd9992ef792e0336c1010cbb5ba638871ac1ca17fa273550a464e19b3874e755e298b9056de4b70d353248ed44c7fc406d25886521cb5c66ef620b8d47fbbd2f6b70d040cb3ff557d67c39586162125ae6f55008d8f88f742bf5747f61c048d66c9e70e73bc6b4bd103450491f9597144b837f887c6225aed30183cd383bd34ed983394f56db0f1d8b3f6a6f2df19328a46d08e3aa21a6e90050bb3e7001fe8bdff133bca0b70fd18b17573fd7e9178beafcbd3ef5c8fa3fcf039eef2a7cc98aa013701e1cdb37590fad9c5aea4c1eb1561c0c9d42db2000354aa2b8096839bf89fe703944d31cc5200aa7a520ea86850f98681f3671a2073b5549264acd325f81ec1926f2dba8ba5eefe1a68ddde3dab875972214e27fc5a1dd5b3efcc59216a08aceb14d0395917df3d9a20173d69828a61ac053533195e65aa0d5dbe33595b049652c6a31fcbb1c22e436ae7f3e5931723166af0f030acd87f30ae6c1bcb0dcc02f62c32a1e18dd762f26ac903001ef8acaf60cf7e630cb4f8b6918ff1ef01981e09ec2a17cfe362cdcb374f48a54ba687afa338f9426fc42067fa86ceca2e9705bb7a7f2d1f6945976ec31d4468a520316f31c94a1163dc26238a8f1d9310ad2914d9f2db760bf305e81378d5a4e073f5e09262c2fe24c70d94aaf3337a9af46d535516fb319e495df37e0db06c80920d4b6e34fd44a65eef0d33d552462e4b78a1c7f2459dc4b28a2abaf45d36836972dce43e5c07994afa877a01ac5ac3da62b091357e7de006a9d11fe0f58307c4dc51c1371ac5fe08482a90f573090f50103ae63dd564692bf9b0cc6cc92e98b2b67f17af800797ee2c7b2a1c7a7e840dd46fa8d777edbd5998e230dd0cab33fc5bae1f08eb5165776bcd9dce2a1b13ffa56d7d0ac1d2aa73ce59664e262e5e8a4599bea9203a7e159;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he8fe077b041fa2e9a7894b6e41738eed5d832339f0a68f61d5f00101a85921506f4be185b9d9aac340ad204b47e0b2ec71ee2ae0595f9e26468ac2164e50a742c19b749c9928c62ab24bf94d3c6f4848dd294f50333900338b718e11aafd3334026c1d5b138891a52b6c7ca921490d6cdfc8c542317a7cf4820320b3b44d6f2f2d54bfee26be5c93d1c345bd3146d2f1d68b43d6c66617be17e68d6eaeb9a120b827b8fd346c955a73594238772085ce5504ae635d481b025e356ff503258a722915e30cfdaee64c4c0070cef6d17f6a7b7b3ef00f7ce43b18d91d2da0de4a04f1c92308ec907d400a9b41c4cb700710da7333a364ab8d3efdd9d664cfe34260fdf2482067a6d457f7bcef10116e004742686228340e0ec86ad9757a0ab8a527f908088000c39358ad8accf66653775c880b1da621023b9162954e357ad6bcdb562bc841301c0ef3c47d5065ac48ad54c690e238fce7ab3dbb36c886ca9a2c63f8a57855a0a4b9d3e3679e59d513a0ce9f837c4b0c62f8acee1efc8796b5197d44e64c670b05151d11f26593b1865e9431746fa967cc4a1b1ce7d4eb2b5c05f92607c6de54b1404ca29fdb83c8bedf1dd18f70657af7f3b952cd1617a4bbdfb196fec36ae48d9d1ad03aaf3f110cb6e9a31e2800c4cc6c9454b5b2aeab8f772959e2701ea3bcac1f9f214c5b42b3dce4c4f8dc41caab255eac2ed0985a7f26489b67e42b4c9b46e69181ddfef8b28ff822302fa6d8d52701382d2dd2a6da7fdc91d3291c6ecc5ea3d110a2b6e31f900a93bf225a6ec343832caaa91ac4e62d4ef6dbea654d625264f3ea82047cebafd05d290c1b0c8960165a5ce193f824f1953f08a1107b78b34736d85e340ccd1855e946bb586556bdcb998f6ef1383cb4a2c21c1dcf652a42ad738f577f0cb2bb2bac17606e84ba1aa69e7114e98ab237405484a17eb1fe76309114d979b0483a7d81472a87ee85941b455c50f313a6389e50b0010a63be6b71a586eed6a492a729e355f2482b673de48869f8da0f48f2aa1de111012101b5c3f4221182fc4e3e8c012f883c83e04cee315324fc22616a63904fa4a31a2c85d77c4d6f5a4f580635c4b06d048a78e49d8f5627cfcda22e5cf3d9b5282d7b003ddcb089471a87373d1b52fd8ac80a580b24fea74150986a9063ee6b083e61f8feb0cd8fcac48ae45be8d473eb107bd606efafb2d451e56cf3121abfc84007f39414daf646784c7dbb9bddf4245f22c98a8ff45a5e4d28812ed485d3ab340e95583ccbebe35e918b96dbdd6831f09f606aaa04847db1757a7c0d52d9408b6a41522dd2e76cfee8feee68a417410bab0804299277cc4ee02a2006389662f20430f647586d90bc95b2bebd9656cfad07a22bdc58c943be4c9cdc4bede9b644e16cf5ebca6fff3f96425d789fb38949713317b40f320a23a91134;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h92759d0c9232e462e3257d142a445ff05d03f151ad9062db8f62a53765122e34ef422ce8b4074495aa5916ee9418e05d1247baa88cd260064b61d379d1c057a2244f274b117cb942f6ab8c11744e477f1cfa497f989e07e315867e343aacb90dabbf6cc35bee4b1f779cbfde859e047f0b1b4621b1f2714480d84d2cc47c8e82fc720a6afe1dc1c8c26bd8e6707c2c5fdc20439c30a9f36df1f40d8faaa340c840961ea53e6ebdb66ed2e5233a4e248bdade1684f2487c2fbe591505cf34154488a02222d4cf9807d5c401cfdc4310cb365cf1e05f5c4d7b585f7ed8ca39aadf002a1946ea259b78c59c3d926c44829b87a568feefee4cefb7176c2fa744da755f4a03bafe937114f7a7ade7acf40f0ff8d0b238b94760be9803cb7a290a17aa0ce1eade98c6ab2b42cb5dc760749037c023159aca1a06b0dbace6ba1456eba8b147b1d69747e0fd06c7630674f28b31567f6033923493aa6ce671faa21b799d59397fe0fba511ec70bcc81059a3554f2d78475b956b00aafc2a157b49d9359b162a71582b912bbd37034233a4cd9e7d3ff3bf0aff290ddb59f8cf29f00b2f87d552df922950ce40f0cafad12cd004221eb5ff6ed28a1dd106236aace288fd0d8476b7bed10d2f8f5b8120e5c7f23d45e9fdd1b34c449caadbd70bd7bb99941498d5f76f2e40454c108cd5ae753484e0514743bde53feae295fc76b5da439d6f791793c465e5addfe752d682fde0c5df88bffffffc5a2dd6c0947d75a6d16098bc754cbb7067481ba12069a8197f4ec6bb56929e4ce4c03c4cb508ed954bc8c1c7df095f3925440317f7d8b62872e250d3cfe37b3044a8c67a3a25b91d2f72852cd550e0497e3b255d99fb8d6665590a5b2362d053b8618246ee9a064cae73c196587eb44ead46f35fc57e4c78314a302c42b9c801ec9606ac7da571aeee95e54bb2ecaf1156a3686b4763a164d00e7ce11b11ef582ebe42efe4fd03fe85dc605f85cd5196b27570c1c394b825fd7848bda05382e1036b485fe9ac1a249efc23d4cd9f3f1a746c50a902dba392a58227638095af81cfd05a6fa2c58e9e0970c4e244cb9b09c25976a5b80ae2ab7165969c84c654ef33308f1fcc7a60d53a872133769ffb6eebb8949690828bbbb68904ef69cdfd58383f4e46f28aa49a50ee7f6ef0e335880eddc4370f784ea88f729bad06c4f89f42138e14a1ae9886cde7c3f9c2f152c23c5dc7f5d4e672476c15ce0391ad65a08e8897d0e4a1fa3e7e0c24142e4bda267cc868f9df202a87b52ffebe6547253eadb4f9ce31d58e1be6cbfd2433616b672b3bb9ef7c1d0cfb574efe6715e350567cf782c0a70a88e21a2d8e96ab42d84c1df1cb6f4ca637c3383d2513225595a6eec0e220318f99ac806ac83c19b78da7d5aa0344fcfd8c8a4f746c73dc84bf11be40aaf3f5c751a7f6dedb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bde1b6bf332334cc9899eeb810f1890edcbb3a94b828d98fc50caa9e31ff10578a87898a4e2da19bb35b4e3a8141fb3bc6e00653a1d7ea80d6accb0a7506bdf3560efcb7988c863b49e5ef4ceb8b410e9cc29d5e88ae5f6a04930780f575c2819750f3e75c36c1cf80bf80c10ebed7ed98284332c9ebef91e65758c0b51754a92120100e7d830825a68d7b519ba5dddd28b4ce28a02c26000bb579b564550b8f3b158655ddf60f0ac708a7c39ed7f2d1ecb81feb284e98d4cf2e26f15fb0c489c2563a21897be755e9f68ddd1ac4b405a79c56739340c16b09736dac7e5c5a0f67c7e505dd9cf7611c1cdffc2276c558a246bd4a903661a092697bfe0b56265a00f3e799667b6269e156082ef4a3ee7e4cf93f8bcbea1b8a0180bbd03dc1624900d07060e4f416d4762a35e09549951c31a17fc889253be107a420ae024f6fffe0f7973328d08e959ce514dd76c2cfbcdb734df8b4c4cecc16d9af84881e5f9547282461dcfc695cf03c5d8ed249d1bf17ecc92aab1ecf89e20fd853a0808550d8758ff77cacb714a461ae6441409c334d459a16f7c0b75eb1cdf07089981529bbcc0d701453365e9356547c46d9d4bd1587df81eb85b17e096e64df53c8445e8e8a8b51ae828f95c681e0baf8f3d04b1927cf51f6bdcf2535bfd4c6c8d56868d00f6f7c4edf7c53870587d9e548920a8f14a4a8832d07c7901ba982bf6bb7f17fd54108e28b02bf5f78a474ee66a4cfe58f0bbccfa3e59552d9e6da8ee85c07cb445bc0c1b7437cd8649740fc84f587d1354ba961031c03e636983c998992289c8730292c4c7899395d1a585780ac8824df09de69631def758841aa725f634e899990608e44e0885698d630138c72f47a60b6c0fd4eb19c184568dab8967251b92261c4cfc61a5726cd7788ab818f5071be7d36662bd31aad92367e9b9eaa7df4c2e1aec6462f97d5d5c973cdc2ff508bded547a515864ecc47b0b3ff31f112d712e6b8d47891bcbdfd1ec3f020a75d51fa5492d699a8dea1f4136c416cceeea27969d84a14a67cfc7222fff6371b57121cccc4a76dd1ad66693f954c67bea49a34391bdab07cf79808d263cd7abe7c38af253dc45b52e1f9a7d636f569230d8a57cee27736de5ea25ebae51038ec8a2ece49f7ed149ad59444fb60f4779fce83dc5d8f5949c02c4ebf49d4df244e9c773b39aecea7b5af94003ff828b372c93033ae2aa64a8f88b7ed8848988a680c61b8fb206ac7a69de7a9e67fb639004349efe67753a633975ca1858f6fe9ee972cae993cb1265e46cbc3471b30c04a682dde640e342b31237348d60221cd47582120c7ea6d6c9cea5b68d959c27c11a08b9a2d12b4d763983c9d24b2c2b58f7708f8d5066ab9e3c7966b6678addf724c7532b2e2c7073e534b9ec6154e19339ddaeb3ec41f077076ff119976c602486;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha18752ef67cc70dc220a189b189c58c36ae2ca75e212d91e30929b6b3a8b2c2be96002f82150d75e3807acfa36d46446ca08eb6fef06729c54bb017d4363851dc258aef9ee2825f586198dcdc0df442eb8828c58b3b570aec0d41bcfb9ccfe8b457150a0ec1a52690ace9f30c37bd504d5bf71d0f25f71f7bd13e952c1231eac5d79bc0e068486ff5c656aca55e18582a670a342b918c752e4c471d26904dd247eeb91c3def9da16d36f935870d9646466645ae4122029bf073b47f6d6b2c887607697507984b93e2d6fb446686c13afda8a281ccb0690345f30da92d9ac9910b00825fbdc8bfae566aa916ca46d858a118199338a344436d61a720ba320de908182d3f4fd786d0acb33111d53102ec551ee6a8c035e4ab7e14f22df54e207b36e33525fb37d91a88670cc4c3272b2317f830f48a529c62c15449c006ac86004cd272267743c657afba64c6236dd23803ff4a2bd5a3bd0877cbde8d66fdeec28386eaca3f00a2ca912b475e70bb7fed9a33038f98e69e537be923b5eace622d727de89cb3980c72cecb80cfdab9a1073e4d4b93d9f29e454f1cd2213fc96bd309d7014eec97c4f79faa355a8edc554de5c70ba0076d89af73cfe4d6871df81055ea0deed9b09a06821b9fad76f032ec1846ac344edddd2f12c985110238215066782065fefec4b18bd2016d05584c55371105ddda9eb8b59fdd70e8e52f4682a59cf7ee4040b36718e1bad459f51d42d57a644ea50fc46b0eb56241fd089e2261b55d67a86328888196c2455ccedf990a104a3f2522e5acdc4d308d2c18f3a6b21e84f2668721a9a21c2d74919676039b76e6cd65722216a9586e6dc6cbf2c0af9b045f8dbae8f3e7d2d7cd076e6f62068151f75f50e5bd67fdcce3103bb463a5d5b01d419969db9b639197727ce6e8a21ec7c8d97677f063c9fa1d52202172c8d04d6e9388d5452aa2dbadde56f87ce6767ad4ef74cb49bc3119aba415dc919129367301bef04d317185bfd365b3a6c3b3b9fca6f0752c0c7ce7f391fb3fae4748af70933e2773ffbb71114378eaf1c702df9cfffdd11998d0dd094aeba913be1e6578d1928cd49207545a6e5c6a0087c79a633d079260431a6519eb144fa80da9f6c8bb37dc7a84b4efdf4da268c6f6cc39a96e1670f97bba9192165c115a634f33b776933b45e9030c0bb09ca866cfff48a9f45bd4a887c5f26d5be53f555295c1e42ff5d7ff2cedb4f30ab0c611ca37472a2c6ce537db33dcac3676be8bb44cd6c330fad662d40bc3e86309d235cfd0d7008d88b2bcd39c66b27c89d03c204a27441f1d93771b0e0a2b492d2ddd11a297be42d721e8411357a239ad3c0c968e82bc400410576b257cecfbf107cfc87cc6ec7a36191912aad53eea09d21dcae4aa127a1f0f369096b1ade97f4ab4468120f77e108c54fbad902dc19b4824a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7156cd1f3d2b542aea8651415a019111c2b0e60362ebca94597687fb0b3a91883c4fb893d2e1b41637032f8a7b275ba7ac71212e60109b96a490e7838d587d90bed93c9d419148c22e61bbc7031152c9661a775286c41178a1cc3b409df7286c9dadeb43010bbd76b3c0415ab030fb9266f2d6a7cf7a283205107ed4d04af9b62975b045ea88841625c09dd6f24c26b0c150fa16b9088580e63fae0abfb91632a274ab9b661f12f09aad304fc68a1dac6c665633e9f460baf3454f33bccd177bf7d8876644d20d2c08c20ad16830397cbc5aa9d80c4bd0cb7691a60257afe9fea5eb175b4d4915703e560e81a39cb0bc88b2114d313961aea167e1aec137e1b3ded36b08ee3cb8399a3aa6ceb4d20bead69c2caafcab03fe2b8deeef133803c40b98a3e2f4fe2f7b97c3e028adfcf05b4788dc8977ff8d76bf3b26d032eb7e3bc03b378267bde2e7fa346f14f5e7d25075c41262f0fb2330b7d20f41c61aa3a7ab701b7d6c665ed70280398731db518f25d79081967738334eedacde38ef0b550cb6aba432d08c022e4964dfcdc34746a7de3568b89e5878e05bec11899daa39430c5f89669d91c4484d879aa0c37ed002ee45461576e7669a6713d039f35485a0ff8287fa94349fca6e6ad470927c761fe94fce039196f39d5525e464c1423429c92003121ad55568de3148e9f5cd9110c0790caa10d6e8b45c81578c197024f3edf7e931a3ddcf3dd7cbe873f33c17b1c94887cdd886a9aea28afbf571c3a7152dc334b4b0de5602373ad4533cf822c71b6bf4ad59fdf26b76f4813c1a7ef4ad178d8eb1f6ab25c595d7978a36a6917c5f903d117133b0fde4b871065c53e5c022d32d610fb69e7cd9bc0503248904bcc835da558d9144b8de0452d5990925074e4fd26a4fd84c75d70d81e8eef7b6af0c87fdda9262a23c4d661726baf66af364091e472622dd714c0ecaa01a311876c308d817cea9319b1d48ffdc1c120aee7dedde749a8e6d295a1c2ca4ae4f63de662465e980d8f0dd235c7631b4ae053c18aa2d008770594bfd2bb4d046169d4bdaed8311ab4d9df578d75246aff3e1ecca83a23bd5db445040d8d56a25880a342461e4b264fe31ddb5d8b5038bde2e18847adb2e7f58e40ccbc83a681963776b42860aaff27b181dd1789092044eedeadf09f915c1da524404a8876b66306327b17f78dff95203e5fc3880b63359ca2fb009c70e4fea76b80e2f9e530a514a77c128e8b85e9bbe08777d52da7d69e386d55bbf9c2d62ae4ae597c5300aeea86a91552fee8fc27a487a806d20fbe00d7f2b38f87ef0a193f6651f390e7df415eb654fa51f3952f78096f21df268c35002b6fbf3d9269c7792ec1ef156d4becf230941109b6cad0f3301ef46fa5c6273a49c1b06a7ef4a3d7b738cc5db35072b41c547e98fbda447575cf69772d71365;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bec7c72e87fdc6f8b6156704b601d2927beb45ff59b0b904e41ad611f7ff7a076b02bc34401e92ac5be2cea1b2cc377419b894bad84dabe6271942a8ef56b8c9216f295975ff4ea40186fadfda9b0c9adaaa1b224915deaea96051fbee14a0194e42f35e9d0822b0674935dffe07f944bfec2f8ce87dbad9f2c66b394d1c0e74c9f161229e6645dbf8919d5f5ed5aa1f3d953e77c7ae2340db9dc76b2055566da731d69867c70c06a48fc2f56dd6f1c3b61268e7fa8fd9285e1bc80c7f1670e471acf92252c9e5ae8b5d8a10038a333178d532c9d5ed42597e8206ac01010cd7453687c5c5d3adde5d468afef84f6ac92a7fe51c92c40065fce74a5b943faf0f48ad6180f3454e3ed75f3e15d948a38bd2665fed4a84e181ef1663a112fbdc01f40f1a18f01976fc41e81af532f1aee5e23b87862deae5e4d012beceb9a6790fd04233818f1aab975d4bf81321e19c8a1e15d4db4ddf120cef19f676a1fff89f48abdb2387ddf99922a94092808dcec8e80aa60f08a30560080df149f1ed5b2204340d55c0e774d088b913c5f8203c1d22f88a058166dd84c9427dced1b7d0355932ca8abfe8526c66f84543ed03bca92240555155bcf8b54569384835960052d56bae184c60ff31837819dd8ebdfed6d9f7e33e73633709e582ca11211da167fbcc6ea2bf373f1c898f1b2b3c2cf2a3fe57ad6fbffd80348f8db4113b89cb188565950385b0245bc5338993ef502f3cc039732e5b67d7c6c511590d067cc6887830a962642cbdd3097d4392518a4bdda8bcd43cabfb43094c3bfc546882d24ff184168a78e91aa4eb52e0dac2943ab9a506841a06b4850d289dc8140b85f25c3a40275f63f8798005e5cb74eacbb0a6b4ba5156c4ec87962abec0721407cab8520ccae0a98b2e0a646a34fddf884baf89fc0edc5826bbc5d609e030572e737989c6d5cde387cae9d25dcfd954d9cee15092788b6654ef66b06b0a9984bf41beb25cc21c1b177a148856ebb77094558b354ad693883d9848e7972b5161e8a22b7bde78fd2290efa3727e3038df1683969e2c2637891914edf746bf724b0acc0641c56115f6602808443a315928f047a737e366736cda2200f2bc6158513efdbded70e4b665e355bb021fd9cc506495c177e4a038bfcdbd63aa5956e277fae7307ea5e791b1c73c857367e75a3ee8ff2b7415cdb31ff9ca5fde1cf70b83b562e122987f40218fd46e56bb10bb27fb140194c2518c5acdd711f1a6c35bb00fb1743a90cd65ae0c8862abed4e32feb4559e45851a1c0206998e35bbdf8351c0c8672845de35fcaae70b7556fcc51be20d5ad7c2a195b36a3d828898ef3a3bb7c1fc00f54bab460c8484e6de1674b8168a98978bd71fe715e4007afe92a89f930192f4a3ce2a320a41b2b2f2f289143f99a50391439e00ada40d87556e616a95595;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3be63764c6f3fee5b08d361e93da2ba61b26ee1283ebf0f80482b3f60c2fdd9ec56bf0c8b108018212a42b23207a302f48db54ccf18a3512d3fbcd72f94dae5e56c7588ac276293e7aca622947875e15db61e9dff8a8526d7e0af027a5f56c1423027e01350b0f6f4ed9961581ea0657410879302d004d98512f8ca4b720c8c73f82249f34b64bd71e67c5f76e17e0c941d64bc313cb88b23fd45623f75802d55305bd4d69f50ad06eaeadf9a4dcfd94721397a50744c64006e4e9283a977dbc8fdd05c94aa4efe2110a5152914109568f1ae76dff43aa28f1720b6473815805c8066bff96e9aacad222f38052a0c9930ccd3f51a5ce0d6c9b2329a9360a0085f0472e4dc992c755039ee04e50a878cba363bd695f36827ec772cf5f1792e873e5ad94c047d83dd33856e2a76039772be252ce82ac5af3f1c507ecc0002ddf71ac2212698e4c098a2ef3b18b7f99a2929323a8baba106a603f2cb2936d1ed3082463247e89ab0cbbbd1b1850d2c30fe5be3c3c77ece444b8de9673549702b2827b739ef193f3ab678c3bd349a6b69f97ac3c28ef5e8a7be5d5aa793c08bcd2aa6a1c68bdf765f104274954a8cfb9f479668ec15cbad4605c950c3a89baba7d3b43d91794d9db46d4a60b8a673ffc81f38cac9f97239a127622868b85829873cf6c829e1ae876434a650181b03d575b600ee4788bebd4e9e84fcbc21faa01d2081f78a7998cd1141b2ad380b039c9a5ac01be5f9823ddc3a1aefe4b6365cdc0d1ac2775e98dd7088c4236f8390ec70ead7365ba39cb615893e7e0e6fa20618d11d29351b2398e77e501035fea88ff7a62c6931693c63585d9664fbd0fc174ea36f4540c05e2dc6f93e7a9652001c2ba0889c2fe385a44c8f839ba02597a6360090bda8c4c8fcc1c64f1201631173e06e592906d8112702831fa224a82f8ba49589ea31c0f0637b102e18b9e172210e143fe0875bf9131746be6988dbd91b383a0b2911cccde4f17549f180672c540dd333b660db9670b6e8e03dd990e7f130f5947a3e1f04ab4d3ba5671869ffdba21ee17a30b57e06e260b8068cbefa071f878814128592cad84840edeb6a7c0a1f38c8879cc4af426342fbc605558f4b75118ff65b4dfb2fb526348e680be0dc44a1ba5a83976a5cd92c877b1ff96a249d6f344e4f676ad4b3aabc08f6cb11b4895b339a612524e4978a6a87e4874d547f07d7478729e06c5a234cde57f1989d48bb11d19890263bc1b42e089629d3a1b303f05e828bb8eab01ffd3cacb992ffb0a2347b56a6e8f6603a8087c52f2b36af4ea2f7dd378310b5e84978ab40284386e79344a3d4e853e7715181ded561fccf0c1ec8f6fdf4d74283ca1320f31897b17a4f9550435f25ed012cef9d387b2f7c55cf9425de8176d8e94050ac8e073929adb572208a36eaa104eb9ce424dc3915d24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd5c7b19acf9b072b933ae69537941586cdb31547204a5c882e280b17f61ad0b313a71a3ee21fede8ce6eae32fa4e904398e991401fd34f2360935ef741450f8da954c5e5bee92a7a6dfbe8c8979053868ce4dee8fe528e7528506f23fb7c03e26d064d6312c43d165b463f388dd0b181cb2be16c35c86c26acd45f3648e1d9d1fa8bc447eade28c99d3c110a36681f2fcfb9a2fb6f2aff039e121110f35cf70af761fcc831eff7dd6e033c026ecbe97ff8c90112704cf30157131d788b9253952f7e1ebe95f530c25e0d7845a6a5c0130ae3b3333899130671b155843f2209f0631dcc5481d7acb5d87bc36e6526a522787650509ca88caeb77acb89b0cced69bb6bbf2b0b614ed33c07d8357d04d33ee916d52b6ab94a084c5abc33cb60fd2be3bd657cb1298f618065ccc06a41a35fa8500bba5348e46ce72dbf9a4b78b6e91f3b9b8a8fa5dddb4d5e42f5428d3ceb35a75deee2894bc6fed4022721fee1481cab2845271dbc4905655b4c6004b15b428b1b0671c747d762031f90e47e92bda4a50bd45f6a10274d3c35e4127717ec0102d70a90a037f1c81bd328e30d034877f930c9445bd594e368c9dfc41761085b4a77b48efee1b08a50e709c4f795e0a676be5fb9da9f1694727044b23980c02bf4476a245a54490e0f5f83c08188200461cae5a311a4c88d55138013ef8eb22cd928a5efbaaaa5e41dce13f396da043d5230098082ff94b610d32b1a25aa9286138f4716a9da0e3b4c4c65153b82dbc8f5ac1022085124ec51911765bafe5cc29a4089fc39f2a260a0095834f434c759f2c8a194184f8b9ef3e60f30a778095599180e7c9f1bdebd7aa8dc073ea631bdf107cecef7be62cdbbcc74b4c8855ef8f7c13b91a7bf65f4265a86a62db7c02fae06cb380e758e893c4416543cb39efb0ed7f5c61fb2ce5f65cd196d1f5939baa40a72ffa39f8cfc81179bab0fb71a3e5682d0cbb5388315a3959baf0038ba798cba340c12250972f67af9f18ad7571ba3831dc8a6c62e0b8e5e9d46761460ea83c17353b1153d6c430335b81fae224af8277731bee2b5c7986e41f90f76ef837a0c2b8c45983a9c05c75f0b6fb0437c896e3c135aa615487165f43d375ad82dad8a89562b1107a9f6e0e020fc079b8330ca97030980fd10958248f1a733cecbb0b3df4ebe4af428713f2bbe05463d71796401ff872ff78cc8188706b3aeb805f319ec6239d6cbd3921349e05fd00a66eb2687e6815ba1f4bdfb16e53a10aa23954ce868867ca2af425e7d897d6f598d8882410d6b6cf60a1848dcf49b0fc6678560978775f190cf47b58e4996206b62ff4422bfc93c37a7374d72c93a02382b8a3799cac5cefb1f4bc7fbca4bd5a5802d0d1e288ff56455665f5948d80e2706e01eb5f3b3517f933c5ea0ee21fb17fdd42cfdec29088b64fe37c904d7146c;
        #1
        $finish();
    end
endmodule
