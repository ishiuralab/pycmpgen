module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    compressor2_1_162_16 compressor2_1_162_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_162_16(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    rowadder2_1_23 rowadder2_1inst(
        .src0({comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [0:0] dst22);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [32:0] stage1_0;
   wire [47:0] stage1_1;
   wire [63:0] stage1_2;
   wire [91:0] stage1_3;
   wire [74:0] stage1_4;
   wire [70:0] stage1_5;
   wire [59:0] stage1_6;
   wire [53:0] stage1_7;
   wire [89:0] stage1_8;
   wire [82:0] stage1_9;
   wire [60:0] stage1_10;
   wire [57:0] stage1_11;
   wire [72:0] stage1_12;
   wire [77:0] stage1_13;
   wire [77:0] stage1_14;
   wire [53:0] stage1_15;
   wire [48:0] stage1_16;
   wire [27:0] stage1_17;
   wire [10:0] stage2_0;
   wire [29:0] stage2_1;
   wire [15:0] stage2_2;
   wire [36:0] stage2_3;
   wire [29:0] stage2_4;
   wire [29:0] stage2_5;
   wire [29:0] stage2_6;
   wire [38:0] stage2_7;
   wire [29:0] stage2_8;
   wire [51:0] stage2_9;
   wire [25:0] stage2_10;
   wire [28:0] stage2_11;
   wire [33:0] stage2_12;
   wire [26:0] stage2_13;
   wire [29:0] stage2_14;
   wire [50:0] stage2_15;
   wire [17:0] stage2_16;
   wire [34:0] stage2_17;
   wire [8:0] stage2_18;
   wire [0:0] stage2_19;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [18:0] stage3_2;
   wire [13:0] stage3_3;
   wire [14:0] stage3_4;
   wire [11:0] stage3_5;
   wire [10:0] stage3_6;
   wire [13:0] stage3_7;
   wire [16:0] stage3_8;
   wire [19:0] stage3_9;
   wire [14:0] stage3_10;
   wire [12:0] stage3_11;
   wire [15:0] stage3_12;
   wire [15:0] stage3_13;
   wire [9:0] stage3_14;
   wire [17:0] stage3_15;
   wire [14:0] stage3_16;
   wire [10:0] stage3_17;
   wire [10:0] stage3_18;
   wire [7:0] stage3_19;
   wire [0:0] stage3_20;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [10:0] stage4_2;
   wire [5:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [6:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [6:0] stage4_9;
   wire [9:0] stage4_10;
   wire [11:0] stage4_11;
   wire [6:0] stage4_12;
   wire [5:0] stage4_13;
   wire [7:0] stage4_14;
   wire [5:0] stage4_15;
   wire [5:0] stage4_16;
   wire [9:0] stage4_17;
   wire [3:0] stage4_18;
   wire [4:0] stage4_19;
   wire [3:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [4:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [2:0] stage5_8;
   wire [4:0] stage5_9;
   wire [3:0] stage5_10;
   wire [3:0] stage5_11;
   wire [5:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [2:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [5:0] stage5_18;
   wire [5:0] stage5_19;
   wire [3:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[8]},
      {stage0_3[16]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[9]},
      {stage0_3[17]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[10]},
      {stage0_3[18]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[11]},
      {stage0_3[19]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[12]},
      {stage0_3[20]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[13]},
      {stage0_3[21]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27]},
      {stage1_5[0],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[1],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[2],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[3],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[4],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[5],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[6],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[7],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[8],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[9],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[10],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[11],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[12],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[13],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[14],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[15],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[16],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[17],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc606_5 gpc49 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[18],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc606_5 gpc50 (
      {stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[19],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc606_5 gpc51 (
      {stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[20],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc606_5 gpc52 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[21],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc606_5 gpc53 (
      {stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[22],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[6],stage1_5[23],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[7],stage1_5[24],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[8],stage1_5[25],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[9],stage1_5[26],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[10],stage1_5[27],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[11],stage1_5[28],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[12],stage1_5[29],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[13],stage1_5[30],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[14],stage1_5[31],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[15],stage1_5[32],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[16],stage1_5[33],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[17],stage1_5[34],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[18],stage1_5[35],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[19],stage1_5[36],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[20],stage1_5[37],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[21],stage1_5[38],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[22],stage1_5[39],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[23],stage1_5[40],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[24],stage1_5[41],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[25],stage1_5[42],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[20],stage1_6[26],stage1_5[43],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[21],stage1_7[21],stage1_6[27],stage1_5[44]}
   );
   gpc606_5 gpc76 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[22],stage1_7[22],stage1_6[28],stage1_5[45]}
   );
   gpc606_5 gpc77 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[23],stage1_7[23],stage1_6[29],stage1_5[46]}
   );
   gpc606_5 gpc78 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[24],stage1_7[24],stage1_6[30],stage1_5[47]}
   );
   gpc606_5 gpc79 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[25],stage1_7[25],stage1_6[31],stage1_5[48]}
   );
   gpc606_5 gpc80 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[26],stage1_7[26],stage1_6[32],stage1_5[49]}
   );
   gpc606_5 gpc81 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[27],stage1_7[27],stage1_6[33],stage1_5[50]}
   );
   gpc606_5 gpc82 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[28],stage1_7[28],stage1_6[34],stage1_5[51]}
   );
   gpc606_5 gpc83 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[29],stage1_7[29],stage1_6[35],stage1_5[52]}
   );
   gpc606_5 gpc84 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[30],stage1_7[30],stage1_6[36],stage1_5[53]}
   );
   gpc606_5 gpc85 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[31],stage1_7[31],stage1_6[37],stage1_5[54]}
   );
   gpc606_5 gpc86 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[32],stage1_7[32],stage1_6[38],stage1_5[55]}
   );
   gpc606_5 gpc87 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[33],stage1_7[33],stage1_6[39],stage1_5[56]}
   );
   gpc606_5 gpc88 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[34],stage1_7[34],stage1_6[40],stage1_5[57]}
   );
   gpc606_5 gpc89 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[35],stage1_7[35],stage1_6[41],stage1_5[58]}
   );
   gpc606_5 gpc90 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[36],stage1_7[36],stage1_6[42],stage1_5[59]}
   );
   gpc606_5 gpc91 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[37],stage1_7[37],stage1_6[43],stage1_5[60]}
   );
   gpc606_5 gpc92 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[38],stage1_7[38],stage1_6[44],stage1_5[61]}
   );
   gpc606_5 gpc93 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[39],stage1_7[39],stage1_6[45],stage1_5[62]}
   );
   gpc606_5 gpc94 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[40],stage1_7[40],stage1_6[46],stage1_5[63]}
   );
   gpc606_5 gpc95 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[41],stage1_7[41],stage1_6[47],stage1_5[64]}
   );
   gpc606_5 gpc96 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[42],stage1_7[42],stage1_6[48],stage1_5[65]}
   );
   gpc606_5 gpc97 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[43],stage1_7[43],stage1_6[49],stage1_5[66]}
   );
   gpc606_5 gpc98 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[44],stage1_7[44],stage1_6[50],stage1_5[67]}
   );
   gpc606_5 gpc99 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[45],stage1_7[45],stage1_6[51],stage1_5[68]}
   );
   gpc606_5 gpc100 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[46],stage1_7[46],stage1_6[52],stage1_5[69]}
   );
   gpc606_5 gpc101 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[47],stage1_7[47],stage1_6[53],stage1_5[70]}
   );
   gpc606_5 gpc102 (
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[48],stage1_7[48],stage1_6[54]}
   );
   gpc606_5 gpc103 (
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[49],stage1_7[49],stage1_6[55]}
   );
   gpc606_5 gpc104 (
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[50],stage1_7[50],stage1_6[56]}
   );
   gpc606_5 gpc105 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[51],stage1_7[51],stage1_6[57]}
   );
   gpc606_5 gpc106 (
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[52],stage1_7[52],stage1_6[58]}
   );
   gpc606_5 gpc107 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[53],stage1_7[53],stage1_6[59]}
   );
   gpc606_5 gpc108 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[6],stage1_9[33],stage1_8[54]}
   );
   gpc606_5 gpc109 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[7],stage1_9[34],stage1_8[55]}
   );
   gpc606_5 gpc110 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[8],stage1_9[35],stage1_8[56]}
   );
   gpc606_5 gpc111 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[9],stage1_9[36],stage1_8[57]}
   );
   gpc606_5 gpc112 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[10],stage1_9[37],stage1_8[58]}
   );
   gpc606_5 gpc113 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[11],stage1_9[38],stage1_8[59]}
   );
   gpc615_5 gpc114 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_9[0]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[12],stage1_9[39],stage1_8[60]}
   );
   gpc615_5 gpc115 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_9[1]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[13],stage1_9[40],stage1_8[61]}
   );
   gpc615_5 gpc116 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86]},
      {stage0_9[2]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[14],stage1_9[41],stage1_8[62]}
   );
   gpc615_5 gpc117 (
      {stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_9[3]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[15],stage1_9[42],stage1_8[63]}
   );
   gpc615_5 gpc118 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_9[4]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[16],stage1_9[43],stage1_8[64]}
   );
   gpc615_5 gpc119 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_9[5]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[17],stage1_9[44],stage1_8[65]}
   );
   gpc615_5 gpc120 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_9[6]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[18],stage1_9[45],stage1_8[66]}
   );
   gpc615_5 gpc121 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_9[7]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[19],stage1_9[46],stage1_8[67]}
   );
   gpc615_5 gpc122 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_9[8]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[20],stage1_9[47],stage1_8[68]}
   );
   gpc615_5 gpc123 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_9[9]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[21],stage1_9[48],stage1_8[69]}
   );
   gpc615_5 gpc124 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_9[10]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[22],stage1_9[49],stage1_8[70]}
   );
   gpc615_5 gpc125 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_9[11]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[23],stage1_9[50],stage1_8[71]}
   );
   gpc615_5 gpc126 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_9[12]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[24],stage1_9[51],stage1_8[72]}
   );
   gpc615_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_9[13]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[25],stage1_9[52],stage1_8[73]}
   );
   gpc615_5 gpc128 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_9[14]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[26],stage1_9[53],stage1_8[74]}
   );
   gpc606_5 gpc129 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[27],stage1_9[54]}
   );
   gpc606_5 gpc130 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[28],stage1_9[55]}
   );
   gpc606_5 gpc131 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[29],stage1_9[56]}
   );
   gpc606_5 gpc132 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[30],stage1_9[57]}
   );
   gpc606_5 gpc133 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[31],stage1_9[58]}
   );
   gpc606_5 gpc134 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[32],stage1_9[59]}
   );
   gpc606_5 gpc135 (
      {stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[33],stage1_9[60]}
   );
   gpc606_5 gpc136 (
      {stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[34],stage1_9[61]}
   );
   gpc606_5 gpc137 (
      {stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[35],stage1_9[62]}
   );
   gpc606_5 gpc138 (
      {stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[36],stage1_9[63]}
   );
   gpc606_5 gpc139 (
      {stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[37],stage1_9[64]}
   );
   gpc606_5 gpc140 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[38],stage1_9[65]}
   );
   gpc606_5 gpc141 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[39],stage1_9[66]}
   );
   gpc606_5 gpc142 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[40],stage1_9[67]}
   );
   gpc606_5 gpc143 (
      {stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[41],stage1_9[68]}
   );
   gpc606_5 gpc144 (
      {stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[42],stage1_9[69]}
   );
   gpc606_5 gpc145 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[43],stage1_9[70]}
   );
   gpc606_5 gpc146 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[44],stage1_9[71]}
   );
   gpc606_5 gpc147 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[45],stage1_9[72]}
   );
   gpc606_5 gpc148 (
      {stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[46],stage1_9[73]}
   );
   gpc606_5 gpc149 (
      {stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[47],stage1_9[74]}
   );
   gpc606_5 gpc150 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[42],stage1_11[42],stage1_10[48],stage1_9[75]}
   );
   gpc615_5 gpc151 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[126]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[43],stage1_11[43],stage1_10[49],stage1_9[76]}
   );
   gpc615_5 gpc152 (
      {stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_10[127]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[44],stage1_11[44],stage1_10[50],stage1_9[77]}
   );
   gpc615_5 gpc153 (
      {stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131], stage0_10[132]},
      {stage0_11[144]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[24],stage1_12[45],stage1_11[45],stage1_10[51]}
   );
   gpc615_5 gpc154 (
      {stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage0_11[145]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[25],stage1_12[46],stage1_11[46],stage1_10[52]}
   );
   gpc615_5 gpc155 (
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142]},
      {stage0_11[146]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[26],stage1_12[47],stage1_11[47],stage1_10[53]}
   );
   gpc615_5 gpc156 (
      {stage0_10[143], stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147]},
      {stage0_11[147]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[27],stage1_12[48],stage1_11[48],stage1_10[54]}
   );
   gpc615_5 gpc157 (
      {stage0_10[148], stage0_10[149], stage0_10[150], stage0_10[151], stage0_10[152]},
      {stage0_11[148]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[28],stage1_12[49],stage1_11[49],stage1_10[55]}
   );
   gpc615_5 gpc158 (
      {stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_11[149]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[29],stage1_12[50],stage1_11[50],stage1_10[56]}
   );
   gpc606_5 gpc159 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[30],stage1_12[51],stage1_11[51]}
   );
   gpc606_5 gpc160 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[7],stage1_13[31],stage1_12[52]}
   );
   gpc606_5 gpc161 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[8],stage1_13[32],stage1_12[53]}
   );
   gpc606_5 gpc162 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[9],stage1_13[33],stage1_12[54]}
   );
   gpc606_5 gpc163 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[10],stage1_13[34],stage1_12[55]}
   );
   gpc606_5 gpc164 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[11],stage1_13[35],stage1_12[56]}
   );
   gpc606_5 gpc165 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[12],stage1_13[36],stage1_12[57]}
   );
   gpc606_5 gpc166 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[13],stage1_13[37],stage1_12[58]}
   );
   gpc606_5 gpc167 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[14],stage1_13[38],stage1_12[59]}
   );
   gpc606_5 gpc168 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[15],stage1_13[39],stage1_12[60]}
   );
   gpc606_5 gpc169 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[10],stage1_14[16],stage1_13[40],stage1_12[61]}
   );
   gpc606_5 gpc170 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[11],stage1_14[17],stage1_13[41],stage1_12[62]}
   );
   gpc606_5 gpc171 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[12],stage1_14[18],stage1_13[42],stage1_12[63]}
   );
   gpc606_5 gpc172 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[13],stage1_14[19],stage1_13[43],stage1_12[64]}
   );
   gpc606_5 gpc173 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[14],stage1_14[20],stage1_13[44],stage1_12[65]}
   );
   gpc606_5 gpc174 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[15],stage1_14[21],stage1_13[45],stage1_12[66]}
   );
   gpc606_5 gpc175 (
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[16],stage1_14[22],stage1_13[46],stage1_12[67]}
   );
   gpc606_5 gpc176 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[17],stage1_14[23],stage1_13[47],stage1_12[68]}
   );
   gpc606_5 gpc177 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[18],stage1_14[24],stage1_13[48],stage1_12[69]}
   );
   gpc606_5 gpc178 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[19],stage1_14[25],stage1_13[49],stage1_12[70]}
   );
   gpc606_5 gpc179 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[20],stage1_14[26],stage1_13[50],stage1_12[71]}
   );
   gpc606_5 gpc180 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[21],stage1_14[27],stage1_13[51],stage1_12[72]}
   );
   gpc606_5 gpc181 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[21],stage1_15[22],stage1_14[28],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[22],stage1_15[23],stage1_14[29],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[23],stage1_15[24],stage1_14[30],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[24],stage1_15[25],stage1_14[31],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[25],stage1_15[26],stage1_14[32],stage1_13[56]}
   );
   gpc606_5 gpc186 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[26],stage1_15[27],stage1_14[33],stage1_13[57]}
   );
   gpc606_5 gpc187 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[27],stage1_15[28],stage1_14[34],stage1_13[58]}
   );
   gpc606_5 gpc188 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[28],stage1_15[29],stage1_14[35],stage1_13[59]}
   );
   gpc606_5 gpc189 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[29],stage1_15[30],stage1_14[36],stage1_13[60]}
   );
   gpc606_5 gpc190 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[30],stage1_15[31],stage1_14[37],stage1_13[61]}
   );
   gpc606_5 gpc191 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[31],stage1_15[32],stage1_14[38],stage1_13[62]}
   );
   gpc606_5 gpc192 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[32],stage1_15[33],stage1_14[39],stage1_13[63]}
   );
   gpc606_5 gpc193 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[33],stage1_15[34],stage1_14[40],stage1_13[64]}
   );
   gpc606_5 gpc194 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[34],stage1_15[35],stage1_14[41],stage1_13[65]}
   );
   gpc606_5 gpc195 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[35],stage1_15[36],stage1_14[42],stage1_13[66]}
   );
   gpc606_5 gpc196 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[36],stage1_15[37],stage1_14[43],stage1_13[67]}
   );
   gpc606_5 gpc197 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[37],stage1_15[38],stage1_14[44],stage1_13[68]}
   );
   gpc606_5 gpc198 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[38],stage1_15[39],stage1_14[45],stage1_13[69]}
   );
   gpc606_5 gpc199 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[39],stage1_15[40],stage1_14[46],stage1_13[70]}
   );
   gpc606_5 gpc200 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[40],stage1_15[41],stage1_14[47],stage1_13[71]}
   );
   gpc606_5 gpc201 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[41],stage1_15[42],stage1_14[48],stage1_13[72]}
   );
   gpc606_5 gpc202 (
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[42],stage1_15[43],stage1_14[49],stage1_13[73]}
   );
   gpc606_5 gpc203 (
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[43],stage1_15[44],stage1_14[50],stage1_13[74]}
   );
   gpc606_5 gpc204 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[44],stage1_15[45],stage1_14[51],stage1_13[75]}
   );
   gpc606_5 gpc205 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[45],stage1_15[46],stage1_14[52],stage1_13[76]}
   );
   gpc606_5 gpc206 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[46],stage1_15[47],stage1_14[53],stage1_13[77]}
   );
   gpc117_4 gpc207 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[156]},
      {1'b0},
      {stage1_17[26],stage1_16[47],stage1_15[48],stage1_14[54]}
   );
   gpc117_4 gpc208 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage0_15[157]},
      {1'b0},
      {stage1_17[27],stage1_16[48],stage1_15[49],stage1_14[55]}
   );
   gpc1_1 gpc209 (
      {stage0_0[160]},
      {stage1_0[31]}
   );
   gpc1_1 gpc210 (
      {stage0_0[161]},
      {stage1_0[32]}
   );
   gpc1_1 gpc211 (
      {stage0_2[152]},
      {stage1_2[54]}
   );
   gpc1_1 gpc212 (
      {stage0_2[153]},
      {stage1_2[55]}
   );
   gpc1_1 gpc213 (
      {stage0_2[154]},
      {stage1_2[56]}
   );
   gpc1_1 gpc214 (
      {stage0_2[155]},
      {stage1_2[57]}
   );
   gpc1_1 gpc215 (
      {stage0_2[156]},
      {stage1_2[58]}
   );
   gpc1_1 gpc216 (
      {stage0_2[157]},
      {stage1_2[59]}
   );
   gpc1_1 gpc217 (
      {stage0_2[158]},
      {stage1_2[60]}
   );
   gpc1_1 gpc218 (
      {stage0_2[159]},
      {stage1_2[61]}
   );
   gpc1_1 gpc219 (
      {stage0_2[160]},
      {stage1_2[62]}
   );
   gpc1_1 gpc220 (
      {stage0_2[161]},
      {stage1_2[63]}
   );
   gpc1_1 gpc221 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc222 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc223 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc224 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc225 (
      {stage0_3[128]},
      {stage1_3[58]}
   );
   gpc1_1 gpc226 (
      {stage0_3[129]},
      {stage1_3[59]}
   );
   gpc1_1 gpc227 (
      {stage0_3[130]},
      {stage1_3[60]}
   );
   gpc1_1 gpc228 (
      {stage0_3[131]},
      {stage1_3[61]}
   );
   gpc1_1 gpc229 (
      {stage0_3[132]},
      {stage1_3[62]}
   );
   gpc1_1 gpc230 (
      {stage0_3[133]},
      {stage1_3[63]}
   );
   gpc1_1 gpc231 (
      {stage0_3[134]},
      {stage1_3[64]}
   );
   gpc1_1 gpc232 (
      {stage0_3[135]},
      {stage1_3[65]}
   );
   gpc1_1 gpc233 (
      {stage0_3[136]},
      {stage1_3[66]}
   );
   gpc1_1 gpc234 (
      {stage0_3[137]},
      {stage1_3[67]}
   );
   gpc1_1 gpc235 (
      {stage0_3[138]},
      {stage1_3[68]}
   );
   gpc1_1 gpc236 (
      {stage0_3[139]},
      {stage1_3[69]}
   );
   gpc1_1 gpc237 (
      {stage0_3[140]},
      {stage1_3[70]}
   );
   gpc1_1 gpc238 (
      {stage0_3[141]},
      {stage1_3[71]}
   );
   gpc1_1 gpc239 (
      {stage0_3[142]},
      {stage1_3[72]}
   );
   gpc1_1 gpc240 (
      {stage0_3[143]},
      {stage1_3[73]}
   );
   gpc1_1 gpc241 (
      {stage0_3[144]},
      {stage1_3[74]}
   );
   gpc1_1 gpc242 (
      {stage0_3[145]},
      {stage1_3[75]}
   );
   gpc1_1 gpc243 (
      {stage0_3[146]},
      {stage1_3[76]}
   );
   gpc1_1 gpc244 (
      {stage0_3[147]},
      {stage1_3[77]}
   );
   gpc1_1 gpc245 (
      {stage0_3[148]},
      {stage1_3[78]}
   );
   gpc1_1 gpc246 (
      {stage0_3[149]},
      {stage1_3[79]}
   );
   gpc1_1 gpc247 (
      {stage0_3[150]},
      {stage1_3[80]}
   );
   gpc1_1 gpc248 (
      {stage0_3[151]},
      {stage1_3[81]}
   );
   gpc1_1 gpc249 (
      {stage0_3[152]},
      {stage1_3[82]}
   );
   gpc1_1 gpc250 (
      {stage0_3[153]},
      {stage1_3[83]}
   );
   gpc1_1 gpc251 (
      {stage0_3[154]},
      {stage1_3[84]}
   );
   gpc1_1 gpc252 (
      {stage0_3[155]},
      {stage1_3[85]}
   );
   gpc1_1 gpc253 (
      {stage0_3[156]},
      {stage1_3[86]}
   );
   gpc1_1 gpc254 (
      {stage0_3[157]},
      {stage1_3[87]}
   );
   gpc1_1 gpc255 (
      {stage0_3[158]},
      {stage1_3[88]}
   );
   gpc1_1 gpc256 (
      {stage0_3[159]},
      {stage1_3[89]}
   );
   gpc1_1 gpc257 (
      {stage0_3[160]},
      {stage1_3[90]}
   );
   gpc1_1 gpc258 (
      {stage0_3[161]},
      {stage1_3[91]}
   );
   gpc1_1 gpc259 (
      {stage0_8[147]},
      {stage1_8[75]}
   );
   gpc1_1 gpc260 (
      {stage0_8[148]},
      {stage1_8[76]}
   );
   gpc1_1 gpc261 (
      {stage0_8[149]},
      {stage1_8[77]}
   );
   gpc1_1 gpc262 (
      {stage0_8[150]},
      {stage1_8[78]}
   );
   gpc1_1 gpc263 (
      {stage0_8[151]},
      {stage1_8[79]}
   );
   gpc1_1 gpc264 (
      {stage0_8[152]},
      {stage1_8[80]}
   );
   gpc1_1 gpc265 (
      {stage0_8[153]},
      {stage1_8[81]}
   );
   gpc1_1 gpc266 (
      {stage0_8[154]},
      {stage1_8[82]}
   );
   gpc1_1 gpc267 (
      {stage0_8[155]},
      {stage1_8[83]}
   );
   gpc1_1 gpc268 (
      {stage0_8[156]},
      {stage1_8[84]}
   );
   gpc1_1 gpc269 (
      {stage0_8[157]},
      {stage1_8[85]}
   );
   gpc1_1 gpc270 (
      {stage0_8[158]},
      {stage1_8[86]}
   );
   gpc1_1 gpc271 (
      {stage0_8[159]},
      {stage1_8[87]}
   );
   gpc1_1 gpc272 (
      {stage0_8[160]},
      {stage1_8[88]}
   );
   gpc1_1 gpc273 (
      {stage0_8[161]},
      {stage1_8[89]}
   );
   gpc1_1 gpc274 (
      {stage0_9[157]},
      {stage1_9[78]}
   );
   gpc1_1 gpc275 (
      {stage0_9[158]},
      {stage1_9[79]}
   );
   gpc1_1 gpc276 (
      {stage0_9[159]},
      {stage1_9[80]}
   );
   gpc1_1 gpc277 (
      {stage0_9[160]},
      {stage1_9[81]}
   );
   gpc1_1 gpc278 (
      {stage0_9[161]},
      {stage1_9[82]}
   );
   gpc1_1 gpc279 (
      {stage0_10[158]},
      {stage1_10[57]}
   );
   gpc1_1 gpc280 (
      {stage0_10[159]},
      {stage1_10[58]}
   );
   gpc1_1 gpc281 (
      {stage0_10[160]},
      {stage1_10[59]}
   );
   gpc1_1 gpc282 (
      {stage0_10[161]},
      {stage1_10[60]}
   );
   gpc1_1 gpc283 (
      {stage0_11[156]},
      {stage1_11[52]}
   );
   gpc1_1 gpc284 (
      {stage0_11[157]},
      {stage1_11[53]}
   );
   gpc1_1 gpc285 (
      {stage0_11[158]},
      {stage1_11[54]}
   );
   gpc1_1 gpc286 (
      {stage0_11[159]},
      {stage1_11[55]}
   );
   gpc1_1 gpc287 (
      {stage0_11[160]},
      {stage1_11[56]}
   );
   gpc1_1 gpc288 (
      {stage0_11[161]},
      {stage1_11[57]}
   );
   gpc1_1 gpc289 (
      {stage0_14[140]},
      {stage1_14[56]}
   );
   gpc1_1 gpc290 (
      {stage0_14[141]},
      {stage1_14[57]}
   );
   gpc1_1 gpc291 (
      {stage0_14[142]},
      {stage1_14[58]}
   );
   gpc1_1 gpc292 (
      {stage0_14[143]},
      {stage1_14[59]}
   );
   gpc1_1 gpc293 (
      {stage0_14[144]},
      {stage1_14[60]}
   );
   gpc1_1 gpc294 (
      {stage0_14[145]},
      {stage1_14[61]}
   );
   gpc1_1 gpc295 (
      {stage0_14[146]},
      {stage1_14[62]}
   );
   gpc1_1 gpc296 (
      {stage0_14[147]},
      {stage1_14[63]}
   );
   gpc1_1 gpc297 (
      {stage0_14[148]},
      {stage1_14[64]}
   );
   gpc1_1 gpc298 (
      {stage0_14[149]},
      {stage1_14[65]}
   );
   gpc1_1 gpc299 (
      {stage0_14[150]},
      {stage1_14[66]}
   );
   gpc1_1 gpc300 (
      {stage0_14[151]},
      {stage1_14[67]}
   );
   gpc1_1 gpc301 (
      {stage0_14[152]},
      {stage1_14[68]}
   );
   gpc1_1 gpc302 (
      {stage0_14[153]},
      {stage1_14[69]}
   );
   gpc1_1 gpc303 (
      {stage0_14[154]},
      {stage1_14[70]}
   );
   gpc1_1 gpc304 (
      {stage0_14[155]},
      {stage1_14[71]}
   );
   gpc1_1 gpc305 (
      {stage0_14[156]},
      {stage1_14[72]}
   );
   gpc1_1 gpc306 (
      {stage0_14[157]},
      {stage1_14[73]}
   );
   gpc1_1 gpc307 (
      {stage0_14[158]},
      {stage1_14[74]}
   );
   gpc1_1 gpc308 (
      {stage0_14[159]},
      {stage1_14[75]}
   );
   gpc1_1 gpc309 (
      {stage0_14[160]},
      {stage1_14[76]}
   );
   gpc1_1 gpc310 (
      {stage0_14[161]},
      {stage1_14[77]}
   );
   gpc1_1 gpc311 (
      {stage0_15[158]},
      {stage1_15[50]}
   );
   gpc1_1 gpc312 (
      {stage0_15[159]},
      {stage1_15[51]}
   );
   gpc1_1 gpc313 (
      {stage0_15[160]},
      {stage1_15[52]}
   );
   gpc1_1 gpc314 (
      {stage0_15[161]},
      {stage1_15[53]}
   );
   gpc606_5 gpc315 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc316 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc317 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[0]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc318 (
      {stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21]},
      {stage1_1[1]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc319 (
      {stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[2]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc320 (
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc321 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc322 (
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc323 (
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc615_5 gpc324 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34]},
      {stage1_3[24]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc325 (
      {stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage1_3[25]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc326 (
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage1_3[26]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc327 (
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_3[27]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc328 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage1_3[28]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc329 (
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_3[29]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc330 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], 1'b0},
      {stage1_3[30]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc331 (
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc332 (
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc333 (
      {stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc334 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc335 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc336 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[16],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc337 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[17],stage2_4[22],stage2_3[22]}
   );
   gpc615_5 gpc338 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[49]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[14],stage2_5[18],stage2_4[23],stage2_3[23]}
   );
   gpc615_5 gpc339 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[50]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[15],stage2_5[19],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc340 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[51]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[16],stage2_5[20],stage2_4[25],stage2_3[25]}
   );
   gpc606_5 gpc341 (
      {stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[10],stage2_6[17],stage2_5[21],stage2_4[26]}
   );
   gpc606_5 gpc342 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[11],stage2_6[18],stage2_5[22],stage2_4[27]}
   );
   gpc606_5 gpc343 (
      {stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[12],stage2_6[19],stage2_5[23],stage2_4[28]}
   );
   gpc615_5 gpc344 (
      {stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_5[60]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[13],stage2_6[20],stage2_5[24],stage2_4[29]}
   );
   gpc606_5 gpc345 (
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[14],stage2_6[21],stage2_5[25]}
   );
   gpc606_5 gpc346 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[5],stage2_7[15],stage2_6[22]}
   );
   gpc606_5 gpc347 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[6],stage2_7[16],stage2_6[23]}
   );
   gpc606_5 gpc348 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[7],stage2_7[17],stage2_6[24]}
   );
   gpc606_5 gpc349 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[4],stage2_8[8],stage2_7[18],stage2_6[25]}
   );
   gpc615_5 gpc350 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52]},
      {stage1_7[6]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[5],stage2_8[9],stage2_7[19],stage2_6[26]}
   );
   gpc615_5 gpc351 (
      {stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57]},
      {stage1_7[7]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[6],stage2_8[10],stage2_7[20],stage2_6[27]}
   );
   gpc615_5 gpc352 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[7],stage2_8[11],stage2_7[21]}
   );
   gpc615_5 gpc353 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[8],stage2_8[12],stage2_7[22]}
   );
   gpc615_5 gpc354 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[9],stage2_8[13],stage2_7[23]}
   );
   gpc615_5 gpc355 (
      {stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[10],stage2_8[14],stage2_7[24]}
   );
   gpc615_5 gpc356 (
      {stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32]},
      {stage1_8[40]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[10],stage2_9[11],stage2_8[15],stage2_7[25]}
   );
   gpc615_5 gpc357 (
      {stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage1_8[41]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[11],stage2_9[12],stage2_8[16],stage2_7[26]}
   );
   gpc615_5 gpc358 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage1_8[42]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[12],stage2_9[13],stage2_8[17],stage2_7[27]}
   );
   gpc606_5 gpc359 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[7],stage2_10[13],stage2_9[14],stage2_8[18]}
   );
   gpc606_5 gpc360 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[8],stage2_10[14],stage2_9[15],stage2_8[19]}
   );
   gpc606_5 gpc361 (
      {stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[9],stage2_10[15],stage2_9[16],stage2_8[20]}
   );
   gpc606_5 gpc362 (
      {stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[10],stage2_10[16],stage2_9[17],stage2_8[21]}
   );
   gpc606_5 gpc363 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[11],stage2_10[17],stage2_9[18],stage2_8[22]}
   );
   gpc606_5 gpc364 (
      {stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[12],stage2_10[18],stage2_9[19],stage2_8[23]}
   );
   gpc606_5 gpc365 (
      {stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[13],stage2_10[19],stage2_9[20],stage2_8[24]}
   );
   gpc606_5 gpc366 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[7],stage2_11[14],stage2_10[20],stage2_9[21]}
   );
   gpc606_5 gpc367 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[8],stage2_11[15],stage2_10[21],stage2_9[22]}
   );
   gpc615_5 gpc368 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46]},
      {stage1_11[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[9],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc369 (
      {stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51]},
      {stage1_11[13]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[10],stage2_11[17],stage2_10[23]}
   );
   gpc615_5 gpc370 (
      {stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_11[14]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[11],stage2_11[18],stage2_10[24]}
   );
   gpc615_5 gpc371 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], 1'b0},
      {stage1_11[15]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[5],stage2_12[12],stage2_11[19],stage2_10[25]}
   );
   gpc1343_5 gpc372 (
      {stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27]},
      {stage1_13[0], stage1_13[1], stage1_13[2]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[4],stage2_13[6],stage2_12[13],stage2_11[20]}
   );
   gpc615_5 gpc373 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage1_12[28]},
      {stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage2_15[1],stage2_14[5],stage2_13[7],stage2_12[14],stage2_11[21]}
   );
   gpc615_5 gpc374 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[29]},
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage2_15[2],stage2_14[6],stage2_13[8],stage2_12[15],stage2_11[22]}
   );
   gpc615_5 gpc375 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[30]},
      {stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20]},
      {stage2_15[3],stage2_14[7],stage2_13[9],stage2_12[16],stage2_11[23]}
   );
   gpc615_5 gpc376 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[31]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[4],stage2_14[8],stage2_13[10],stage2_12[17],stage2_11[24]}
   );
   gpc615_5 gpc377 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[32]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[5],stage2_14[9],stage2_13[11],stage2_12[18],stage2_11[25]}
   );
   gpc615_5 gpc378 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[33]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[6],stage2_14[10],stage2_13[12],stage2_12[19],stage2_11[26]}
   );
   gpc615_5 gpc379 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[34]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[7],stage2_14[11],stage2_13[13],stage2_12[20],stage2_11[27]}
   );
   gpc615_5 gpc380 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], 1'b0},
      {stage1_12[35]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[8],stage2_14[12],stage2_13[14],stage2_12[21],stage2_11[28]}
   );
   gpc606_5 gpc381 (
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[9],stage2_14[13],stage2_13[15],stage2_12[22]}
   );
   gpc606_5 gpc382 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[10],stage2_14[14],stage2_13[16],stage2_12[23]}
   );
   gpc606_5 gpc383 (
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[11],stage2_14[15],stage2_13[17],stage2_12[24]}
   );
   gpc606_5 gpc384 (
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[12],stage2_14[16],stage2_13[18],stage2_12[25]}
   );
   gpc606_5 gpc385 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[13],stage2_14[17],stage2_13[19],stage2_12[26]}
   );
   gpc606_5 gpc386 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[18],stage2_13[20]}
   );
   gpc606_5 gpc387 (
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[19],stage2_13[21]}
   );
   gpc606_5 gpc388 (
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[20],stage2_13[22]}
   );
   gpc606_5 gpc389 (
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[21],stage2_13[23]}
   );
   gpc606_5 gpc390 (
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[22]}
   );
   gpc606_5 gpc391 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[23]}
   );
   gpc606_5 gpc392 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[24]}
   );
   gpc606_5 gpc393 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[25]}
   );
   gpc606_5 gpc394 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[26]}
   );
   gpc606_5 gpc395 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23],stage2_14[27]}
   );
   gpc606_5 gpc396 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24],stage2_14[28]}
   );
   gpc615_5 gpc397 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[24]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[11],stage2_16[16],stage2_15[25],stage2_14[29]}
   );
   gpc615_5 gpc398 (
      {stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[48]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[8],stage2_17[12],stage2_16[17],stage2_15[26]}
   );
   gpc1_1 gpc399 (
      {stage1_0[27]},
      {stage2_0[5]}
   );
   gpc1_1 gpc400 (
      {stage1_0[28]},
      {stage2_0[6]}
   );
   gpc1_1 gpc401 (
      {stage1_0[29]},
      {stage2_0[7]}
   );
   gpc1_1 gpc402 (
      {stage1_0[30]},
      {stage2_0[8]}
   );
   gpc1_1 gpc403 (
      {stage1_0[31]},
      {stage2_0[9]}
   );
   gpc1_1 gpc404 (
      {stage1_0[32]},
      {stage2_0[10]}
   );
   gpc1_1 gpc405 (
      {stage1_1[27]},
      {stage2_1[9]}
   );
   gpc1_1 gpc406 (
      {stage1_1[28]},
      {stage2_1[10]}
   );
   gpc1_1 gpc407 (
      {stage1_1[29]},
      {stage2_1[11]}
   );
   gpc1_1 gpc408 (
      {stage1_1[30]},
      {stage2_1[12]}
   );
   gpc1_1 gpc409 (
      {stage1_1[31]},
      {stage2_1[13]}
   );
   gpc1_1 gpc410 (
      {stage1_1[32]},
      {stage2_1[14]}
   );
   gpc1_1 gpc411 (
      {stage1_1[33]},
      {stage2_1[15]}
   );
   gpc1_1 gpc412 (
      {stage1_1[34]},
      {stage2_1[16]}
   );
   gpc1_1 gpc413 (
      {stage1_1[35]},
      {stage2_1[17]}
   );
   gpc1_1 gpc414 (
      {stage1_1[36]},
      {stage2_1[18]}
   );
   gpc1_1 gpc415 (
      {stage1_1[37]},
      {stage2_1[19]}
   );
   gpc1_1 gpc416 (
      {stage1_1[38]},
      {stage2_1[20]}
   );
   gpc1_1 gpc417 (
      {stage1_1[39]},
      {stage2_1[21]}
   );
   gpc1_1 gpc418 (
      {stage1_1[40]},
      {stage2_1[22]}
   );
   gpc1_1 gpc419 (
      {stage1_1[41]},
      {stage2_1[23]}
   );
   gpc1_1 gpc420 (
      {stage1_1[42]},
      {stage2_1[24]}
   );
   gpc1_1 gpc421 (
      {stage1_1[43]},
      {stage2_1[25]}
   );
   gpc1_1 gpc422 (
      {stage1_1[44]},
      {stage2_1[26]}
   );
   gpc1_1 gpc423 (
      {stage1_1[45]},
      {stage2_1[27]}
   );
   gpc1_1 gpc424 (
      {stage1_1[46]},
      {stage2_1[28]}
   );
   gpc1_1 gpc425 (
      {stage1_1[47]},
      {stage2_1[29]}
   );
   gpc1_1 gpc426 (
      {stage1_3[81]},
      {stage2_3[26]}
   );
   gpc1_1 gpc427 (
      {stage1_3[82]},
      {stage2_3[27]}
   );
   gpc1_1 gpc428 (
      {stage1_3[83]},
      {stage2_3[28]}
   );
   gpc1_1 gpc429 (
      {stage1_3[84]},
      {stage2_3[29]}
   );
   gpc1_1 gpc430 (
      {stage1_3[85]},
      {stage2_3[30]}
   );
   gpc1_1 gpc431 (
      {stage1_3[86]},
      {stage2_3[31]}
   );
   gpc1_1 gpc432 (
      {stage1_3[87]},
      {stage2_3[32]}
   );
   gpc1_1 gpc433 (
      {stage1_3[88]},
      {stage2_3[33]}
   );
   gpc1_1 gpc434 (
      {stage1_3[89]},
      {stage2_3[34]}
   );
   gpc1_1 gpc435 (
      {stage1_3[90]},
      {stage2_3[35]}
   );
   gpc1_1 gpc436 (
      {stage1_3[91]},
      {stage2_3[36]}
   );
   gpc1_1 gpc437 (
      {stage1_5[67]},
      {stage2_5[26]}
   );
   gpc1_1 gpc438 (
      {stage1_5[68]},
      {stage2_5[27]}
   );
   gpc1_1 gpc439 (
      {stage1_5[69]},
      {stage2_5[28]}
   );
   gpc1_1 gpc440 (
      {stage1_5[70]},
      {stage2_5[29]}
   );
   gpc1_1 gpc441 (
      {stage1_6[58]},
      {stage2_6[28]}
   );
   gpc1_1 gpc442 (
      {stage1_6[59]},
      {stage2_6[29]}
   );
   gpc1_1 gpc443 (
      {stage1_7[43]},
      {stage2_7[28]}
   );
   gpc1_1 gpc444 (
      {stage1_7[44]},
      {stage2_7[29]}
   );
   gpc1_1 gpc445 (
      {stage1_7[45]},
      {stage2_7[30]}
   );
   gpc1_1 gpc446 (
      {stage1_7[46]},
      {stage2_7[31]}
   );
   gpc1_1 gpc447 (
      {stage1_7[47]},
      {stage2_7[32]}
   );
   gpc1_1 gpc448 (
      {stage1_7[48]},
      {stage2_7[33]}
   );
   gpc1_1 gpc449 (
      {stage1_7[49]},
      {stage2_7[34]}
   );
   gpc1_1 gpc450 (
      {stage1_7[50]},
      {stage2_7[35]}
   );
   gpc1_1 gpc451 (
      {stage1_7[51]},
      {stage2_7[36]}
   );
   gpc1_1 gpc452 (
      {stage1_7[52]},
      {stage2_7[37]}
   );
   gpc1_1 gpc453 (
      {stage1_7[53]},
      {stage2_7[38]}
   );
   gpc1_1 gpc454 (
      {stage1_8[85]},
      {stage2_8[25]}
   );
   gpc1_1 gpc455 (
      {stage1_8[86]},
      {stage2_8[26]}
   );
   gpc1_1 gpc456 (
      {stage1_8[87]},
      {stage2_8[27]}
   );
   gpc1_1 gpc457 (
      {stage1_8[88]},
      {stage2_8[28]}
   );
   gpc1_1 gpc458 (
      {stage1_8[89]},
      {stage2_8[29]}
   );
   gpc1_1 gpc459 (
      {stage1_9[54]},
      {stage2_9[23]}
   );
   gpc1_1 gpc460 (
      {stage1_9[55]},
      {stage2_9[24]}
   );
   gpc1_1 gpc461 (
      {stage1_9[56]},
      {stage2_9[25]}
   );
   gpc1_1 gpc462 (
      {stage1_9[57]},
      {stage2_9[26]}
   );
   gpc1_1 gpc463 (
      {stage1_9[58]},
      {stage2_9[27]}
   );
   gpc1_1 gpc464 (
      {stage1_9[59]},
      {stage2_9[28]}
   );
   gpc1_1 gpc465 (
      {stage1_9[60]},
      {stage2_9[29]}
   );
   gpc1_1 gpc466 (
      {stage1_9[61]},
      {stage2_9[30]}
   );
   gpc1_1 gpc467 (
      {stage1_9[62]},
      {stage2_9[31]}
   );
   gpc1_1 gpc468 (
      {stage1_9[63]},
      {stage2_9[32]}
   );
   gpc1_1 gpc469 (
      {stage1_9[64]},
      {stage2_9[33]}
   );
   gpc1_1 gpc470 (
      {stage1_9[65]},
      {stage2_9[34]}
   );
   gpc1_1 gpc471 (
      {stage1_9[66]},
      {stage2_9[35]}
   );
   gpc1_1 gpc472 (
      {stage1_9[67]},
      {stage2_9[36]}
   );
   gpc1_1 gpc473 (
      {stage1_9[68]},
      {stage2_9[37]}
   );
   gpc1_1 gpc474 (
      {stage1_9[69]},
      {stage2_9[38]}
   );
   gpc1_1 gpc475 (
      {stage1_9[70]},
      {stage2_9[39]}
   );
   gpc1_1 gpc476 (
      {stage1_9[71]},
      {stage2_9[40]}
   );
   gpc1_1 gpc477 (
      {stage1_9[72]},
      {stage2_9[41]}
   );
   gpc1_1 gpc478 (
      {stage1_9[73]},
      {stage2_9[42]}
   );
   gpc1_1 gpc479 (
      {stage1_9[74]},
      {stage2_9[43]}
   );
   gpc1_1 gpc480 (
      {stage1_9[75]},
      {stage2_9[44]}
   );
   gpc1_1 gpc481 (
      {stage1_9[76]},
      {stage2_9[45]}
   );
   gpc1_1 gpc482 (
      {stage1_9[77]},
      {stage2_9[46]}
   );
   gpc1_1 gpc483 (
      {stage1_9[78]},
      {stage2_9[47]}
   );
   gpc1_1 gpc484 (
      {stage1_9[79]},
      {stage2_9[48]}
   );
   gpc1_1 gpc485 (
      {stage1_9[80]},
      {stage2_9[49]}
   );
   gpc1_1 gpc486 (
      {stage1_9[81]},
      {stage2_9[50]}
   );
   gpc1_1 gpc487 (
      {stage1_9[82]},
      {stage2_9[51]}
   );
   gpc1_1 gpc488 (
      {stage1_12[66]},
      {stage2_12[27]}
   );
   gpc1_1 gpc489 (
      {stage1_12[67]},
      {stage2_12[28]}
   );
   gpc1_1 gpc490 (
      {stage1_12[68]},
      {stage2_12[29]}
   );
   gpc1_1 gpc491 (
      {stage1_12[69]},
      {stage2_12[30]}
   );
   gpc1_1 gpc492 (
      {stage1_12[70]},
      {stage2_12[31]}
   );
   gpc1_1 gpc493 (
      {stage1_12[71]},
      {stage2_12[32]}
   );
   gpc1_1 gpc494 (
      {stage1_12[72]},
      {stage2_12[33]}
   );
   gpc1_1 gpc495 (
      {stage1_13[75]},
      {stage2_13[24]}
   );
   gpc1_1 gpc496 (
      {stage1_13[76]},
      {stage2_13[25]}
   );
   gpc1_1 gpc497 (
      {stage1_13[77]},
      {stage2_13[26]}
   );
   gpc1_1 gpc498 (
      {stage1_15[30]},
      {stage2_15[27]}
   );
   gpc1_1 gpc499 (
      {stage1_15[31]},
      {stage2_15[28]}
   );
   gpc1_1 gpc500 (
      {stage1_15[32]},
      {stage2_15[29]}
   );
   gpc1_1 gpc501 (
      {stage1_15[33]},
      {stage2_15[30]}
   );
   gpc1_1 gpc502 (
      {stage1_15[34]},
      {stage2_15[31]}
   );
   gpc1_1 gpc503 (
      {stage1_15[35]},
      {stage2_15[32]}
   );
   gpc1_1 gpc504 (
      {stage1_15[36]},
      {stage2_15[33]}
   );
   gpc1_1 gpc505 (
      {stage1_15[37]},
      {stage2_15[34]}
   );
   gpc1_1 gpc506 (
      {stage1_15[38]},
      {stage2_15[35]}
   );
   gpc1_1 gpc507 (
      {stage1_15[39]},
      {stage2_15[36]}
   );
   gpc1_1 gpc508 (
      {stage1_15[40]},
      {stage2_15[37]}
   );
   gpc1_1 gpc509 (
      {stage1_15[41]},
      {stage2_15[38]}
   );
   gpc1_1 gpc510 (
      {stage1_15[42]},
      {stage2_15[39]}
   );
   gpc1_1 gpc511 (
      {stage1_15[43]},
      {stage2_15[40]}
   );
   gpc1_1 gpc512 (
      {stage1_15[44]},
      {stage2_15[41]}
   );
   gpc1_1 gpc513 (
      {stage1_15[45]},
      {stage2_15[42]}
   );
   gpc1_1 gpc514 (
      {stage1_15[46]},
      {stage2_15[43]}
   );
   gpc1_1 gpc515 (
      {stage1_15[47]},
      {stage2_15[44]}
   );
   gpc1_1 gpc516 (
      {stage1_15[48]},
      {stage2_15[45]}
   );
   gpc1_1 gpc517 (
      {stage1_15[49]},
      {stage2_15[46]}
   );
   gpc1_1 gpc518 (
      {stage1_15[50]},
      {stage2_15[47]}
   );
   gpc1_1 gpc519 (
      {stage1_15[51]},
      {stage2_15[48]}
   );
   gpc1_1 gpc520 (
      {stage1_15[52]},
      {stage2_15[49]}
   );
   gpc1_1 gpc521 (
      {stage1_15[53]},
      {stage2_15[50]}
   );
   gpc1_1 gpc522 (
      {stage1_17[6]},
      {stage2_17[13]}
   );
   gpc1_1 gpc523 (
      {stage1_17[7]},
      {stage2_17[14]}
   );
   gpc1_1 gpc524 (
      {stage1_17[8]},
      {stage2_17[15]}
   );
   gpc1_1 gpc525 (
      {stage1_17[9]},
      {stage2_17[16]}
   );
   gpc1_1 gpc526 (
      {stage1_17[10]},
      {stage2_17[17]}
   );
   gpc1_1 gpc527 (
      {stage1_17[11]},
      {stage2_17[18]}
   );
   gpc1_1 gpc528 (
      {stage1_17[12]},
      {stage2_17[19]}
   );
   gpc1_1 gpc529 (
      {stage1_17[13]},
      {stage2_17[20]}
   );
   gpc1_1 gpc530 (
      {stage1_17[14]},
      {stage2_17[21]}
   );
   gpc1_1 gpc531 (
      {stage1_17[15]},
      {stage2_17[22]}
   );
   gpc1_1 gpc532 (
      {stage1_17[16]},
      {stage2_17[23]}
   );
   gpc1_1 gpc533 (
      {stage1_17[17]},
      {stage2_17[24]}
   );
   gpc1_1 gpc534 (
      {stage1_17[18]},
      {stage2_17[25]}
   );
   gpc1_1 gpc535 (
      {stage1_17[19]},
      {stage2_17[26]}
   );
   gpc1_1 gpc536 (
      {stage1_17[20]},
      {stage2_17[27]}
   );
   gpc1_1 gpc537 (
      {stage1_17[21]},
      {stage2_17[28]}
   );
   gpc1_1 gpc538 (
      {stage1_17[22]},
      {stage2_17[29]}
   );
   gpc1_1 gpc539 (
      {stage1_17[23]},
      {stage2_17[30]}
   );
   gpc1_1 gpc540 (
      {stage1_17[24]},
      {stage2_17[31]}
   );
   gpc1_1 gpc541 (
      {stage1_17[25]},
      {stage2_17[32]}
   );
   gpc1_1 gpc542 (
      {stage1_17[26]},
      {stage2_17[33]}
   );
   gpc1_1 gpc543 (
      {stage1_17[27]},
      {stage2_17[34]}
   );
   gpc1163_5 gpc544 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc545 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc546 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc547 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc548 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc615_5 gpc549 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc550 (
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage2_4[1]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc606_5 gpc551 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc552 (
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc553 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[4],stage3_6[4],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc554 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[5],stage3_6[5],stage3_5[8],stage3_4[10]}
   );
   gpc606_5 gpc555 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[4],stage3_7[6],stage3_6[6],stage3_5[9]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[5],stage3_7[7],stage3_6[7],stage3_5[10]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[6],stage3_7[8],stage3_6[8],stage3_5[11]}
   );
   gpc615_5 gpc558 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28]},
      {stage2_7[18]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[7],stage3_7[9],stage3_6[9]}
   );
   gpc615_5 gpc559 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[4],stage3_8[8],stage3_7[10]}
   );
   gpc615_5 gpc560 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[5],stage3_8[9],stage3_7[11]}
   );
   gpc615_5 gpc561 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[6],stage3_8[10],stage3_7[12]}
   );
   gpc615_5 gpc562 (
      {stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[7],stage3_8[11],stage3_7[13]}
   );
   gpc606_5 gpc563 (
      {stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[8],stage3_8[12]}
   );
   gpc606_5 gpc564 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[9],stage3_8[13]}
   );
   gpc606_5 gpc565 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[10],stage3_8[14]}
   );
   gpc606_5 gpc566 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[11]}
   );
   gpc606_5 gpc567 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[12]}
   );
   gpc606_5 gpc568 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[13]}
   );
   gpc615_5 gpc569 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46]},
      {stage2_10[18]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[6],stage3_11[10],stage3_10[11],stage3_9[14]}
   );
   gpc615_5 gpc570 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[7],stage3_11[11],stage3_10[12]}
   );
   gpc615_5 gpc571 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], 1'b0},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[5],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc572 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[6],stage3_12[9]}
   );
   gpc606_5 gpc573 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[2],stage3_14[3],stage3_13[7],stage3_12[10]}
   );
   gpc606_5 gpc574 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[3],stage3_14[4],stage3_13[8],stage3_12[11]}
   );
   gpc606_5 gpc575 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[4],stage3_14[5],stage3_13[9],stage3_12[12]}
   );
   gpc606_5 gpc576 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[5],stage3_14[6],stage3_13[10]}
   );
   gpc606_5 gpc577 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[5],stage3_15[6],stage3_14[7],stage3_13[11]}
   );
   gpc606_5 gpc578 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[6],stage3_15[7],stage3_14[8],stage3_13[12]}
   );
   gpc606_5 gpc579 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[7],stage3_15[8],stage3_14[9]}
   );
   gpc615_5 gpc580 (
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[8],stage3_15[9]}
   );
   gpc615_5 gpc581 (
      {stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[9],stage3_15[10]}
   );
   gpc615_5 gpc582 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[6],stage3_16[10],stage3_15[11]}
   );
   gpc615_5 gpc583 (
      {stage2_15[33], stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[7],stage3_16[11],stage3_15[12]}
   );
   gpc615_5 gpc584 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[8],stage3_16[12],stage3_15[13]}
   );
   gpc615_5 gpc585 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[11]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], 1'b0},
      {stage3_19[5],stage3_18[6],stage3_17[9],stage3_16[13],stage3_15[14]}
   );
   gpc606_5 gpc586 (
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[6],stage3_18[7],stage3_17[10],stage3_16[14]}
   );
   gpc1_1 gpc587 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc588 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc589 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc590 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc591 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc592 (
      {stage2_2[2]},
      {stage3_2[5]}
   );
   gpc1_1 gpc593 (
      {stage2_2[3]},
      {stage3_2[6]}
   );
   gpc1_1 gpc594 (
      {stage2_2[4]},
      {stage3_2[7]}
   );
   gpc1_1 gpc595 (
      {stage2_2[5]},
      {stage3_2[8]}
   );
   gpc1_1 gpc596 (
      {stage2_2[6]},
      {stage3_2[9]}
   );
   gpc1_1 gpc597 (
      {stage2_2[7]},
      {stage3_2[10]}
   );
   gpc1_1 gpc598 (
      {stage2_2[8]},
      {stage3_2[11]}
   );
   gpc1_1 gpc599 (
      {stage2_2[9]},
      {stage3_2[12]}
   );
   gpc1_1 gpc600 (
      {stage2_2[10]},
      {stage3_2[13]}
   );
   gpc1_1 gpc601 (
      {stage2_2[11]},
      {stage3_2[14]}
   );
   gpc1_1 gpc602 (
      {stage2_2[12]},
      {stage3_2[15]}
   );
   gpc1_1 gpc603 (
      {stage2_2[13]},
      {stage3_2[16]}
   );
   gpc1_1 gpc604 (
      {stage2_2[14]},
      {stage3_2[17]}
   );
   gpc1_1 gpc605 (
      {stage2_2[15]},
      {stage3_2[18]}
   );
   gpc1_1 gpc606 (
      {stage2_3[30]},
      {stage3_3[7]}
   );
   gpc1_1 gpc607 (
      {stage2_3[31]},
      {stage3_3[8]}
   );
   gpc1_1 gpc608 (
      {stage2_3[32]},
      {stage3_3[9]}
   );
   gpc1_1 gpc609 (
      {stage2_3[33]},
      {stage3_3[10]}
   );
   gpc1_1 gpc610 (
      {stage2_3[34]},
      {stage3_3[11]}
   );
   gpc1_1 gpc611 (
      {stage2_3[35]},
      {stage3_3[12]}
   );
   gpc1_1 gpc612 (
      {stage2_3[36]},
      {stage3_3[13]}
   );
   gpc1_1 gpc613 (
      {stage2_4[26]},
      {stage3_4[11]}
   );
   gpc1_1 gpc614 (
      {stage2_4[27]},
      {stage3_4[12]}
   );
   gpc1_1 gpc615 (
      {stage2_4[28]},
      {stage3_4[13]}
   );
   gpc1_1 gpc616 (
      {stage2_4[29]},
      {stage3_4[14]}
   );
   gpc1_1 gpc617 (
      {stage2_6[29]},
      {stage3_6[10]}
   );
   gpc1_1 gpc618 (
      {stage2_8[28]},
      {stage3_8[15]}
   );
   gpc1_1 gpc619 (
      {stage2_8[29]},
      {stage3_8[16]}
   );
   gpc1_1 gpc620 (
      {stage2_9[47]},
      {stage3_9[15]}
   );
   gpc1_1 gpc621 (
      {stage2_9[48]},
      {stage3_9[16]}
   );
   gpc1_1 gpc622 (
      {stage2_9[49]},
      {stage3_9[17]}
   );
   gpc1_1 gpc623 (
      {stage2_9[50]},
      {stage3_9[18]}
   );
   gpc1_1 gpc624 (
      {stage2_9[51]},
      {stage3_9[19]}
   );
   gpc1_1 gpc625 (
      {stage2_10[24]},
      {stage3_10[13]}
   );
   gpc1_1 gpc626 (
      {stage2_10[25]},
      {stage3_10[14]}
   );
   gpc1_1 gpc627 (
      {stage2_12[31]},
      {stage3_12[13]}
   );
   gpc1_1 gpc628 (
      {stage2_12[32]},
      {stage3_12[14]}
   );
   gpc1_1 gpc629 (
      {stage2_12[33]},
      {stage3_12[15]}
   );
   gpc1_1 gpc630 (
      {stage2_13[24]},
      {stage3_13[13]}
   );
   gpc1_1 gpc631 (
      {stage2_13[25]},
      {stage3_13[14]}
   );
   gpc1_1 gpc632 (
      {stage2_13[26]},
      {stage3_13[15]}
   );
   gpc1_1 gpc633 (
      {stage2_15[48]},
      {stage3_15[15]}
   );
   gpc1_1 gpc634 (
      {stage2_15[49]},
      {stage3_15[16]}
   );
   gpc1_1 gpc635 (
      {stage2_15[50]},
      {stage3_15[17]}
   );
   gpc1_1 gpc636 (
      {stage2_18[6]},
      {stage3_18[8]}
   );
   gpc1_1 gpc637 (
      {stage2_18[7]},
      {stage3_18[9]}
   );
   gpc1_1 gpc638 (
      {stage2_18[8]},
      {stage3_18[10]}
   );
   gpc1_1 gpc639 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc615_5 gpc640 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc641 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[1]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc615_5 gpc642 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[2],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc643 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[3],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc644 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[2],stage4_6[4]}
   );
   gpc615_5 gpc645 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[3],stage4_6[5]}
   );
   gpc615_5 gpc646 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage3_8[12]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[4]}
   );
   gpc615_5 gpc647 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[13]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc648 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc649 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3],stage4_10[5]}
   );
   gpc606_5 gpc650 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4],stage4_10[6]}
   );
   gpc1406_5 gpc651 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc615_5 gpc652 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[0]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[1],stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[4]}
   );
   gpc615_5 gpc653 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[1]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[2],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[5]}
   );
   gpc606_5 gpc654 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage4_18[0],stage4_17[3],stage4_16[3],stage4_15[3],stage4_14[5]}
   );
   gpc615_5 gpc655 (
      {stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[4],stage4_16[4]}
   );
   gpc623_5 gpc656 (
      {stage3_16[12], stage3_16[13], stage3_16[14]},
      {stage3_17[1], stage3_17[2]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], 1'b0},
      {stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[5],stage4_16[5]}
   );
   gpc615_5 gpc657 (
      {stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[2],stage4_18[3],stage4_17[6]}
   );
   gpc1_1 gpc658 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc659 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc660 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc661 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc662 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc663 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc664 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc665 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc666 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc667 (
      {stage3_1[2]},
      {stage4_1[2]}
   );
   gpc1_1 gpc668 (
      {stage3_1[3]},
      {stage4_1[3]}
   );
   gpc1_1 gpc669 (
      {stage3_1[4]},
      {stage4_1[4]}
   );
   gpc1_1 gpc670 (
      {stage3_2[10]},
      {stage4_2[2]}
   );
   gpc1_1 gpc671 (
      {stage3_2[11]},
      {stage4_2[3]}
   );
   gpc1_1 gpc672 (
      {stage3_2[12]},
      {stage4_2[4]}
   );
   gpc1_1 gpc673 (
      {stage3_2[13]},
      {stage4_2[5]}
   );
   gpc1_1 gpc674 (
      {stage3_2[14]},
      {stage4_2[6]}
   );
   gpc1_1 gpc675 (
      {stage3_2[15]},
      {stage4_2[7]}
   );
   gpc1_1 gpc676 (
      {stage3_2[16]},
      {stage4_2[8]}
   );
   gpc1_1 gpc677 (
      {stage3_2[17]},
      {stage4_2[9]}
   );
   gpc1_1 gpc678 (
      {stage3_2[18]},
      {stage4_2[10]}
   );
   gpc1_1 gpc679 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc680 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc681 (
      {stage3_4[14]},
      {stage4_4[4]}
   );
   gpc1_1 gpc682 (
      {stage3_6[10]},
      {stage4_6[6]}
   );
   gpc1_1 gpc683 (
      {stage3_7[12]},
      {stage4_7[6]}
   );
   gpc1_1 gpc684 (
      {stage3_7[13]},
      {stage4_7[7]}
   );
   gpc1_1 gpc685 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc686 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc687 (
      {stage3_8[16]},
      {stage4_8[6]}
   );
   gpc1_1 gpc688 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc689 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc690 (
      {stage3_10[12]},
      {stage4_10[7]}
   );
   gpc1_1 gpc691 (
      {stage3_10[13]},
      {stage4_10[8]}
   );
   gpc1_1 gpc692 (
      {stage3_10[14]},
      {stage4_10[9]}
   );
   gpc1_1 gpc693 (
      {stage3_11[6]},
      {stage4_11[5]}
   );
   gpc1_1 gpc694 (
      {stage3_11[7]},
      {stage4_11[6]}
   );
   gpc1_1 gpc695 (
      {stage3_11[8]},
      {stage4_11[7]}
   );
   gpc1_1 gpc696 (
      {stage3_11[9]},
      {stage4_11[8]}
   );
   gpc1_1 gpc697 (
      {stage3_11[10]},
      {stage4_11[9]}
   );
   gpc1_1 gpc698 (
      {stage3_11[11]},
      {stage4_11[10]}
   );
   gpc1_1 gpc699 (
      {stage3_11[12]},
      {stage4_11[11]}
   );
   gpc1_1 gpc700 (
      {stage3_12[12]},
      {stage4_12[3]}
   );
   gpc1_1 gpc701 (
      {stage3_12[13]},
      {stage4_12[4]}
   );
   gpc1_1 gpc702 (
      {stage3_12[14]},
      {stage4_12[5]}
   );
   gpc1_1 gpc703 (
      {stage3_12[15]},
      {stage4_12[6]}
   );
   gpc1_1 gpc704 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc705 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc706 (
      {stage3_15[16]},
      {stage4_15[4]}
   );
   gpc1_1 gpc707 (
      {stage3_15[17]},
      {stage4_15[5]}
   );
   gpc1_1 gpc708 (
      {stage3_17[8]},
      {stage4_17[7]}
   );
   gpc1_1 gpc709 (
      {stage3_17[9]},
      {stage4_17[8]}
   );
   gpc1_1 gpc710 (
      {stage3_17[10]},
      {stage4_17[9]}
   );
   gpc1_1 gpc711 (
      {stage3_19[6]},
      {stage4_19[3]}
   );
   gpc1_1 gpc712 (
      {stage3_19[7]},
      {stage4_19[4]}
   );
   gpc1_1 gpc713 (
      {stage3_20[0]},
      {stage4_20[3]}
   );
   gpc606_5 gpc714 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc615_5 gpc715 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1343_5 gpc716 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0], stage4_8[1], stage4_8[2]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0]}
   );
   gpc1343_5 gpc717 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc1343_5 gpc718 (
      {stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc7_3 gpc719 (
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], 1'b0},
      {stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc1343_5 gpc720 (
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc207_4 gpc721 (
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], 1'b0},
      {stage4_13[3], stage4_13[4]},
      {stage5_14[1],stage5_13[2],stage5_12[3],stage5_11[3]}
   );
   gpc615_5 gpc722 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc615_5 gpc723 (
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {1'b0},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1],stage5_15[2]}
   );
   gpc1_1 gpc724 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc725 (
      {stage4_2[7]},
      {stage5_2[2]}
   );
   gpc1_1 gpc726 (
      {stage4_2[8]},
      {stage5_2[3]}
   );
   gpc1_1 gpc727 (
      {stage4_2[9]},
      {stage5_2[4]}
   );
   gpc1_1 gpc728 (
      {stage4_2[10]},
      {stage5_2[5]}
   );
   gpc1_1 gpc729 (
      {stage4_4[0]},
      {stage5_4[2]}
   );
   gpc1_1 gpc730 (
      {stage4_4[1]},
      {stage5_4[3]}
   );
   gpc1_1 gpc731 (
      {stage4_4[2]},
      {stage5_4[4]}
   );
   gpc1_1 gpc732 (
      {stage4_4[3]},
      {stage5_4[5]}
   );
   gpc1_1 gpc733 (
      {stage4_4[4]},
      {stage5_4[6]}
   );
   gpc1_1 gpc734 (
      {stage4_5[0]},
      {stage5_5[1]}
   );
   gpc1_1 gpc735 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc736 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc737 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc738 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc739 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc740 (
      {stage4_9[5]},
      {stage5_9[3]}
   );
   gpc1_1 gpc741 (
      {stage4_9[6]},
      {stage5_9[4]}
   );
   gpc1_1 gpc742 (
      {stage4_12[5]},
      {stage5_12[4]}
   );
   gpc1_1 gpc743 (
      {stage4_12[6]},
      {stage5_12[5]}
   );
   gpc1_1 gpc744 (
      {stage4_13[5]},
      {stage5_13[3]}
   );
   gpc1_1 gpc745 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc746 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc747 (
      {stage4_17[6]},
      {stage5_17[2]}
   );
   gpc1_1 gpc748 (
      {stage4_17[7]},
      {stage5_17[3]}
   );
   gpc1_1 gpc749 (
      {stage4_17[8]},
      {stage5_17[4]}
   );
   gpc1_1 gpc750 (
      {stage4_17[9]},
      {stage5_17[5]}
   );
   gpc1_1 gpc751 (
      {stage4_18[0]},
      {stage5_18[2]}
   );
   gpc1_1 gpc752 (
      {stage4_18[1]},
      {stage5_18[3]}
   );
   gpc1_1 gpc753 (
      {stage4_18[2]},
      {stage5_18[4]}
   );
   gpc1_1 gpc754 (
      {stage4_18[3]},
      {stage5_18[5]}
   );
   gpc1_1 gpc755 (
      {stage4_19[0]},
      {stage5_19[1]}
   );
   gpc1_1 gpc756 (
      {stage4_19[1]},
      {stage5_19[2]}
   );
   gpc1_1 gpc757 (
      {stage4_19[2]},
      {stage5_19[3]}
   );
   gpc1_1 gpc758 (
      {stage4_19[3]},
      {stage5_19[4]}
   );
   gpc1_1 gpc759 (
      {stage4_19[4]},
      {stage5_19[5]}
   );
   gpc1_1 gpc760 (
      {stage4_20[0]},
      {stage5_20[0]}
   );
   gpc1_1 gpc761 (
      {stage4_20[1]},
      {stage5_20[1]}
   );
   gpc1_1 gpc762 (
      {stage4_20[2]},
      {stage5_20[2]}
   );
   gpc1_1 gpc763 (
      {stage4_20[3]},
      {stage5_20[3]}
   );
   gpc1_1 gpc764 (
      {stage4_21[0]},
      {stage5_21[0]}
   );
   gpc615_5 gpc765 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc766 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0]},
      {stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc767 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc1163_5 gpc768 (
      {stage5_11[1], stage5_11[2], stage5_11[3]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_13[0]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1343_5 gpc769 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc770 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1]}
   );
   gpc1406_5 gpc771 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[1]}
   );
   gpc1_1 gpc772 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc773 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc774 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc775 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc776 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc777 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc778 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc779 (
      {stage5_7[1]},
      {stage6_7[1]}
   );
   gpc1_1 gpc780 (
      {stage5_9[4]},
      {stage6_9[1]}
   );
   gpc1_1 gpc781 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc782 (
      {stage5_16[1]},
      {stage6_16[1]}
   );
endmodule
module rowadder2_1_23(input [22:0] src0, input [22:0] src1, output [23:0] dst0);
    wire [22:0] gene;
    wire [22:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[22:20]}),
        .S({1'h0, prop[22:20]})
    );
    assign dst0 = {carryout[22], out[22:0]};
endmodule


module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor2_1_162_16 compressor2_1_162_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h37f4bab07de726bb65b36f4c21de4fa373af28aa8dd6468859d1f6c9573a3d2cf68387f88fc0fc7552f2f4d600a50cc6fd43720ec15a7fd4849e244ae33f25ba6e88315f1f9ea7694a11e49e8ce6610105ddfd8fb36abefb289f132f19e9ae10b7750bfd3b3fb9b4fdf054e1dddb7002be0f2750184d431d5d9028fecd9cba5e1690a7241ef68063fc206fcc2d120180fd854ad11038325d770c3251a82089947842ca46ac070737f4608a5ed6e5a520c603098b26df9c2fefa59c623efc5545cc7244084d80873489eec9f56a5c42283730d80ff52e973fc49791dceb2dfa6822199536a4c48e84bd9703a560a87776f88139f5705876285178f5092258c33d827b87c8ba9feb47ba9216fad1b26b418a69cb2ea4a0bd6179b43129edb64ae6e574e79237f558e551a7b6ea366e202afa00e34cfff2cd4e48b94b7e1056c89ded2e6087;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h503ac7a2b6a202aeeaff477912b8b3a8741cdd0bca49419997bede402470d9a87818b713bb2d07dd47ac271e36aab5b7dc0943910b37c16d6b4381242884f9ac4b16f8514d294d61ac03f8f8190dc3aad6f059104c930a6114cef228c900c496799a7408fc693829cd9e1fb86a22a4158f491c4874e1b3c686509db02284687e968100548b9879bf67194e8461498041ee77213a69b7ad7fdfc9af03071fe5fe1a405e32569d88439f557f736c641762faaa6737bf3e9218c3b7cd31f0362106f0321f490c4aacdb631f3fe8b2fa8c86dda2cf79e3176b51b499010caa4a1df62809067fef6777d91026ed95f657621b6c400bbd6a007a080df7d50510a2d6cd49f3941865063ad4f37b0028ed38a5e6aadb9d5150f5374b588a76cf62bab85a6c03f2cf97871d252c08ad33ecd19bc68b38e15e5c2cf9d8592d88272428bcddcf01a272;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4846a2c2c0bd6c270347cd42bc33464b226b7f6ed604d6629cc56cfa9672323bae53e9ded675b390b3aeecf609791758f62105c5dd0943408d6e7a7212aaeb07890818cb39bee03da12b9fa532db6b34f00dcdcb61612d45215d2105b3a8df15e60cfca3c47208bcf62f03b3333524c63cda033ee79f3488a8ce22f7c0b5aa34351ca7ef220d9355e44161a18dc6249516d5ef22c0d6d12fe2110cca43ef1215f3b6c855c01d85873fd3eda9b4c90108c36dbd92448744f9155046dc890cb85a3adbcef68bad0cd329debae24f22fb1c56de8e6949d268560a7c3b0d9bea80028b346e2f2bf2000a869f5d52a39c0ffe948400ad55b286fd6dd152fb87f2eff806412595be423a8153338dbde24e8e483554815f3e5ed3e8ff2da5ab62c7898a6040b5c31a3e41840145c937b74231eaffef744bf3a742eba5c6bfe264a60b411565421b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hed1faa6987eac4f1de1b030822fbabee60e13390839360d28e981748db370e75a73773252e31003fe4e2c9d447200e04013124e93336421616d956a16a81df512afe576e36749639b96b51f39496ba1a9155a47e48b9fc038a93eda75df5a9d64f305b0222ad228595e1af54ef1b8d35de104b4ba671328891940f75c73519b8a98f158e05f78459429c0afb1f09992a1a9dcf9051ca624d585063ea4727b6e75d1e7464aa4b346109285eb66d7cbc7abebc55cfd03fc4254c6e09a14b1874d2b9632c2826e998eb96000f93d4b643533c52555c529ce11d3a5f60a9ba375e20792aac82f040c3379ac571c83fe8f8314fedaaa5ba817853f3d0fc701b16f90d53484c616fa3ba3b8bed1b4369d7b89a95b05e2b74cc9a0f97f2b26b1cdd62a5d41f2c951399310c4b3c74aafcb1c49746ed0c41679592b5cc58c713329d6e98093c10cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1dfcf4cec936c495a4fc10c05c277b20265fd987a842e8ce7b698aadedc78d822080bba664933d8f68a7dd2376fb52ffb05524d4a1205483049b294aee1f3cfc90c4a2d57ca6835a3263b0ebc7b5a5e4f1e58fb0fde0232a74ea3fd3a1bbdbc5a096d684802425560cbb64e7cfdb2a30054dd56d0ef0e6684b2446a1212b3d0b7a7e5d7b3a1e15f7223c740ddfce9a04a06960b0f0cea8dbbd48087016b548fa4cc11ec7598540f9600687b8055a9e1c8f85bf5ec55489979c15bd248c160f65ac2cd3caa1a2dac5a819c92228f19001ffd556de52bd47d72cdcf1f4f76c2b3504126f060462333a13be449c443344f07f7693444eb64a9fbb719145fbf786d1b71dc6f78e8e8f58973b210981d637325fffe8b2c626f6be65be111254dbb86840f513152b26ffa0de259bd2e4ea523c8b316884ea3daad1a953485232b111577b2c96e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hce82479280e3eeadac076bbabaeaadfe81c6133ab6b37495acf8ea0a205f3f5ebf52cf5e47d4adb149b58b4e452ce12a3c865e4338b3427100612416119d05db4c472a2cb4a5fecb03e39bc613e50fce61ff98055a8f873e6b80dc0a625de24d0bc500279ba7ba8a07573ffed97c00397fd234e1a8c634c846caa9caa436628abbcaabf2284aceeeec95a8ac979ea4a1e9a90e75ae6b7e4eaa18a4d7c76af1f4d676e21e74ea0483586d71c740a586cefc01d45a748a8691bd9d5edd85052d098fd7d9090ac4aa5cc7c1fc433eb0bc2a6885a195c70f9b3c482b9d446116e198774d411e7f0dd84a8e158faa02bc5acfb508e76f73e7e56c2521ef54879344a88a72009e496c2a26eae2d4f4b441b8fffa84960f2f58704973a27a327eae13a9fff0f8ed8f7ad180cb27475722ba872d6de1ddbb97b90859b526e1f8a9fabc40d795d72d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hbb0f49516e866c96a90f735a914c3a42ced29ed0e2851c74c4fbb586e460d1d32424c7cbd9a5a3de86b6df656c11f643eb769230daaac25ec7fcd43726acdded90c45707d032795de2406174b93a884d7375eb93882852b75e81d4d4f74503b8b22a78d51da7fda5064130cfc4f3a5445da68038a53b602562658c7228a10808fce2d20cc8479b49fc71b401053c0378e08a80db6fc236167e3f680977ded1443123a094b02bad7a39d9777941aae83417f0260010fb29d494bd043701a936ca2dce4dd302ed4045483c8f5709720e2bb8fcf89366d81dc20d3b36bbdf6c36e1a76a1c6999c704aa1f54524c25fad731e6f84204c2988c20ef2b16027e9bb91dc90caa4aec33f51200f181302e7153e9c5ebc416244f5b6c5f157c9dd0dfcd37c35efc40245117937e0bca3d0ccc12de660f1c169762cea60c4e5fffdbd5126543b23a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5d0108d75affba07a9a8aa62917287da581a3724ee752af068f3c3b1a03f77f2cf9fcfc3eeca37c18bd65da4a39214f33195da5e7d4fb12bcaaa50b2b12db755d2ddb9162e40ef9428fead35f22e38c09c24701bcb01bac534723a860fb10e6a4e93131ef63d4e7e76cb71001fab6ece87abd26218a544a3f94ed222bb1f6f21543675e35beba776a5cc554567b93d0313745dcd57fb6f770fe7bec182fd66532caf8023d4a4332c5ab00741937b4a784a4e098635b0c7c37907bd061aef431895a92b61e91da662d795b644d92af799dd93ff55c0ad1104926b76a3c089b8a1884f92c4bf76226f67a1f52644cf5a91cd4dd10e2ce992871b4666ec2fc67765a0307982df89d097e34facd88d327b9548f09a63fd242ce618f97d474d94f1e9ffbbd4616114619394e55c5edc5e9d7b844089afb3a50f37f043624900f6cd604d0e233d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hcaa13c2b5ccedb7a124536cfb4b40019f972e8cfceae1262f7ee61cad66bef0276d1153e1b5b21e39676ca19237930aac3f872598f89aaf98777188e9c16fa52f8a0d448026413a29ca8f93777112595363f18cd39ac95920de856775d37cc4f729872a3a2f836b1cece60ae4fc5d44f64a7e18c23b8ca8ff8b087db93f789175814c90022ca23f17fbe341d421d4835753988bf70e52712bf1e866b31bbb15ccb46d15fd90cdf470079e16fb18c48fa2ddffcb73c4077865f3394fd10fa64066e3556f8aff249762636575f7679f4adc12f2bc5ed344aa69b1d79deeeb16e87b35d6cb439fc2e57b43bb0ac7e372e8364edba38c334d52416223776f1fe0856152947c853a660c93c57e2aee36e0335c67f52cb1e6714fb94aaecb3e7bd0177eb75865e28d5582586f5f71bb7e652daa5bfda754735a16c9abbd5643d2d92631fe3015e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8064c6f1cab7919b2868eee351e8ccd7a348dc63678c5b399a6d40e274f3d5ec80a442e49793fa047e282a7a9d001ae6bddf2e02a7adde98767655ab2b970b452d27e392a0c416508b6aa2147e6a4ab6f0a72b726f0d10e36a3eb494519fde299102d2349b82983ccfc59d6a11c46c966028e29070999668bed810b6bf5500241443853634cdd3520c7f0d60f4899b32752c118cd954996f4fb8525b4a6fe956fc0293747753b1b26dab51bf1ea6fb0779d0b2c620fbd486ae4a72faa1198aafee93faf851ad37916aebcbdf7f44d671a507611551e66e0193ea5b0a9cb5fe3b5fc950f90e25213a2dff7fb59dbda2432eeed8b25429c01e81d952d0cdf5b1df6874cf8bcc38c7cf1319bc91adf9d1279a4fea0774623aac7dd62133087c4ff1d8da86dd19b73c75ff2e84d71afa6d3bc6370f90ef66a887aa0bde5beca0cecb2b6ee385;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h86cd799b2c9855bc8c02ccd11bac239e70849cda4e035917790691055e2bcb677a4aab318ba50abba85c27b3058126208a4ce22ffd1f4ad2714caf2bd3229a8c8d4efe13cc8795e3b347beaa90bed7812241f5dfa9209f1faa7d8f8dbb89899ca53f0ec937da157646b8ede94a88d7e03a2aa96db78ab6788ad597aff1bad9574933e4c7bcad8667f507cb3cfc1841e033c71fb2f9326f5dffb5e941b86f65debaad7f5f0d7b428e40f2e65f70112d46eae0b5f71487e193c0ff27ac9620acfd91a2a57b9c12e59517de83633d02551c2b4b013a3bad5a1ce687e3016677560851673b179d60b0bea5f9c0cc0358f1544f9c9b157aadeef7719d2c1bbd80336febd69da785b383cb89aa0fd9122adb632244a8053ab265c8fb62ae4c9b31fc16e3453d4bf9b369b576db5ef49185ddc19200dab8006a827509566378f8b5f66ee9c16848;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha85ee0e8ef4c3080a53107fe909690d7061bc6ea565f008e49d8eebee8ddc8946805f8ecc4c18045e748be6629abb6599eff0ce18f4e04bb1cd5fd0f18ee43bf361eea74ab97c17ddce8fef5287b0b9bd964a9ee5cdd31dd2fe5297022c47503a8d803b41106725364ee7ea194de254809354b341c2022b6c04ff57ab72dadce0e81e5fa14f0830f41b54326e0ef0ff7427f68cf58775c69e0a788697fc23acfda7f888d5801802e79f9c1988360e1ed5260068dbf30e724de2c43e107a4a1e5b2ca80166ea9e5b34f04469760f36c2c0de1765c3cfcb173e65b2e72e37fac97aa4cd890521d873761edd8c193b9ffe7565e3806f69b68d17f254af1dce802a5de06536f8cbe0aee049659945dd296bdc1e54458d03f41a0322e80635fba58d3e84569fe10efcbe6aac3bf442064f8d9f0a1bb4c0ae1d91104effe1c9d7957e5d3c10ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfbf6f6ce13cbba0602d1c72156d5d84d1a5755524953bf755b16c6e66b60f0f63fa65a7b6c8fe15462392850e7e7c9d07446f2a143e8bc32157a690500ce8109bbc501371a29b63990618709d324a7b8370919a6e19cfeaa50dd85cccbade60ac1259ea63ace7e56c18715c9c4c85fde4ceac44ffa8c0125e3abda6552d1a4ee2db5dcffd855169a3e4092cba3d8a228d59efc0dcd5d0f9935e0b03d18111ae4241ff2fc44a8552286c3459a7a48b0e840e4dc519312d392b3b5c51013b3e92040763aac29798e38371fff4bea6cc07ff4526a5034a7b5017c51abb6587fca9f929cd7e9b7bc0b56a908dcf7dd150cceebe2122f33af6e4dfa1b3dee580f91143327ed5ffbdef56759eac9ab171de2a2fc9143aa13d5ce7de90e2b6b1d961e40ce7cbe76adb24052f219a7fb282a3f18ac86c2e6a35555eba8a3da1cf1afda7fa35db4e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h652d630d7c82530925f630252603e3f2128fd530e96b55175875e3b8319b4cc5c9a2991c4376ae8be1c923f5571c7d077cd0c49648c54e5ad6fa53f6845d69743e08407e2c558b4bddc23b35b7454a505b3b0729233e337d8d64a7df97a732916d05733715935c4487c271dce76fe9a8346968650065cf1b67ef978e54b0f8137bcb497e63ff20283d304b0f8ede4abdf45e36b82ee1107553ba7052f2a4d62ebeadc0e4129542abe06fe8308b3a1fe732eb0c88533c034c8160966f7b7743d19d2e088943d6c147d19d365e6e8c4c21477c87631e0344904715e2608ccebb7b382c6742403629338eaa4f97910b302e0f1103159dc5db4280860ddcf3405671e47fca29ebbdf1733aa94293385bdf6a908a74cbae9aa019e3c308acc1377a85536b43987f543cd8067d3f68ff59899543b19e003d3760d6a357a6704cd299592aed6ed8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha1e431fb330ca2682291cd9737f0a77761ed76960078e535fcf61cda09cb189ba635d5f273c217a833c35e3c3ff99bfa3ad4c697a273117854031abc3841e31b3e13942dadbe21ee23a9b92d1c4f7ef6df2cc2480240e2623dd7c1f9d15178ebd3a17b490bdede1be55aaade2c1514aa8680e832aa2f3055e398d34b0132235b3afaf97d436e252a9f3680ee797e8ea14be5ff60aabeb6e5aab9f67bcb0542bbc028a7a7595d9d085d0ca3ecbeca5a9920be25a59112f630d65ef55e34aeae3faea49133d9d98e1e8618e33194ffc9a11e08abe8246b4355786dcf369c72da89f887f230fd45f50910c8e5ff61e39bb98e730da1a05890ff62204438f4e6b1726cd6aa7d0f7b5b5ea710a190b4b7b52837d31b3070b98495b346a642c79a415bac71544db5aa698fc5b75dea8a4105869993dc313d6b8bd614ad87d358882ffd7b317429;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h93b562acb38851c25b1ac746aa3415abc03279f6e493594a76568369239ecc10661729ad6292765c20e83ae030ad62778cd1f7d27e9718a7c5b51e6d7f028f2d6f231d91d5a14f4da3ce60a7b91c95e02a12b4f67072de4dab4c357d8ca89424b62431951f6ee91473e62c01abda065b6e1d927347650f11684a1c2d7e091d6adca6bde3bcc1d81b5e54efd315977ed4d3a69ef1cd2562ad07bb3a3e3526ecc6d6e09f2bf56ef699accf107693e5a43157d27ee309ba215e2cbba00ac2e2df38fe6e7619974962d6c8f47b5ab84759333fcc8366c3a30a96bdbff12678640ebd012a3cc4a655b0ab39c530db076698cb2926f2b0a0bb0085005bcaf11bd0d731c421675efe068fe7eb8197f9c4ddfa694585942a11a3b652446b56b963e8e1d55091ec048179d28ebb51f6c3f3e77cef34e05c6c4f8c664386134db7a3881c0188863736;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdffd6e310642a5a56b73bc30c2ac84dbd4001860b16371c8e66cd876b77199ad6a348d1094be12c4275717b22f544828dfc64f93f9bc045a91662f5674614b0b75199f983d4bfbec143a91a26112032281979fb7c6a824edac1095f1a17460047cb841f3fafaeb7661fe88f59fe1476f830131020e394e6b9b413566ee2596ba96d7c8124de7534cdc917eeeef4c2d63ef6b481496832447b69944f2b41bb96a2fa4a000e590f2f00c0f1a20284453cad8d6702f91ba1442eca1e46d6f173920ba3ee2ae80c8ab2c96bf66947b6e5c7cbc2dd9d4330b7cfbd9793a2eabf251aa5230b083a2965b660a1c9d3bfb280ffd891e3cd939478991da8e3859ff121c7054ce72e379d526bb7e15edb97c59c9fe17e5f377c1bc6b4d210d46ed864835251fd3ae7d40917c9005a0ce57b95e7be62823e7836e7a2a68159a67587e1d20f90f12de7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4e8f04c6128ad7679b7ecfe69a30cddd86d5fa36ce6afd0bd070b5d92fa7fe138b4763140346be5c8b630f0d77d069ca8ecbb36b12e27d4cb6d3409fc621a2af4b0be59cf9fd33118a8b630a15b38c814b16d7c9b3879fbbad531c531e040ba10ac138cfe6862872aec65985addfb7744e87b91ae7012830946da46f6edf92a014c02b1c0ebf3348536d09f65d985e8db3c0637c4a4bdfb458ce8f3ded554767005237d60cfd60f282efedbcd3d1dd6f390349615f37cd1155246a40b2f359130e3d72d0f35d528e41d9f47264cfcdff17ffa900b697b60865bd2fcd697248a69e1780a48d2b994e40ee0fe418f07ce5280a18b5401c0692b54dd8e5fdfe4d82ac1dbb637ff8d58344d23cc2802fde3784f65a71ada44b64de82419a2efdc679a97981bb3bd04603f0cd9a55ccdee5de889aa5674684aa8512d4a51c9ca5515a49027e62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc7388707ad4cd7ac52dfd84cb12b9a40264eb6011ae9fc205a024d07b46f99691f613b32e89b652c593e1a5115fccc0edef0a561beacaab2df9a2f6e28807664742d3271ab32c28dddd27c319bedd0f77249c3e3a816698403f713e3f430864cba7290307eeec36db2b9423cd48a8ba9a4b7fad9c151a5c40bb1a57fcf98e5fc3487d3382213e55293c9e889cb4b4e714adb4fcf55921bab3cf62a9d4795e84973c387a30914989a612966713ce4867e90374f8458d46dd5730476bf27ab7478049842cc8568f2c6b8b23c2bf30e57ff5c7ad23b366a1d4a3e7cbaaae8d975a5aa8c2091763ee5b79c0793478c0e9f3a053e2dc234359bb80ad647c2e76aa52531d2b1e6be7f993573a47ef2d54578f250b8f2cfdb6e07dbdc7aac8130a1554365c447c152238640a39fd49f6c4cf46043d905972eba41052b34cc7300b53a7b7d31b279;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf229521d0f79cbffa3591fa8792467286b376c518702bfa3bc637c0cfe8a995ef64c2711e0bf5830ac23f4954e1b605be4a0d1248d0f5a809479dab98acbab459ced7b6b33ad98afccd7803a7aaa6ee391bf22373724daa83f3024830938f8949cda24cf362090cf6b169ffd87b5c8cbb53f145b51aca36734747b9295ca0fa90cd74b5f7ac4ca92787207e7d4b899606a4f4278ef46d44fb8e7bd81ac1373723dc8291c2926feb15d634ad488818039d3c43b6935de13d2a7ca854ad439756baddc798b0579d0f7503d4d51355daa58722bc9df11ab234688f4262f86377d0e36946b1cacb388fb0da6fd64d7672bdfd10344d362e9d5f41939573ada43986e8be45927061680e4c87fd44114c19a77c73f2a691f35514542ed4f9b77239f5405493e4276a0299c423c2753aed8df00798ef6322b4b63480ac40c52a32a9f1077ee1fe4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfd8d84d9a37473786fec8b47686b999bba3cfce691441d4a0a92fd103503c5f0b70f59177668f21221ab500cced12f79426ea13e8921ea8b60b1b1f930fda701403c777d04b9e6f33476944694598f28e374fc45ca2a92f6e5022afeca10fb96c259f1e48800e23b99a4cf03043d2f13b08e858d2cf1b98ef3a1ad702d85cd49e48dcb0c83a7a9270903371402597fa082d9bde73418d56e1e406a6d15ef46fc24f79a80be50ae5d2e589acdc3269036c585976a1a49c7985eeaeb194536de7bb8d63a1b5001e776506c7300436e692cf25b3f4c80e0841fa360ccf68694f8873462b60895ad5abf89ca6139b99be93f2c32d4564d00cf8ab656533cd871398c31e7987d23d150deb38821119f760ea3dc3e154a018c0da7336dbfb1fffe7825cbde607c25d8c8d75a7fa5ccfc64d84f369139eb770c911c005c8fc0c2cf1d73ad4c5ced;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6df7aacd3c51cedefecacba8d8a62bab1af146389160ee2070f8a1d7a66f18944ec96a3061c5e2187d70409b7ebf4fa18a43b35b1f6ff030621f3f4a6cc931124354f564da795af5bbb28b1652c703e62ae59c205dc014cc16c62a58d93ae008258367dd1324a60c188dbf7b3cb4cf937f85458acf1c74dac4048d4d56d7a2262bcf4473240b796be83c41504ae215160a5382b32f9f4f4acf8d0d06d97b4289bb4e09d1a2efc10890ffa793ca89f8281c8ac4f35e89d0d9c735a2b3211a390a220a1437b6eda86255cdd584d694e1ea50bb39568d4bde17512aa3aee74ca70f27f447610a14d7c25369c902327792779341f16cf1ebe731aab8a611604065d5e6ccc7f62d103811340386ed860dc43129fe0aeaf4e174f876337a454a9007fb8cfd5879426c0856c335e6524ab0685c4fc4d7a8876241a57097586bead33ddd345fbf87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h48bcb648232cb2a82161457215190a55581d6e60cc5515193f05dbae34f410dfef29c0aebd3fc515d60ee9d194c4bfb6007e96f55a59e95f1afc0702d678382d0a68fd26ab8a6ba7023e1b249865f1059338bb64db7991ff3fc9ce594f834d3b91db24d6dd02d70eb36b4217636d8aa687960fb63c569aaeed507529c3aa6a979fd648bc042fc220d688f28eb6921e9b3bf67a20f8ba2dc5aa1c72bf087b1c889aba9173c85bd7d1d2ba9c2c950326e9373ad806b84ce889408c8da846703e07268a68779f9b2a94a009c21023cad03c72da6619eefb7bb0b16b1ad2715ac1ef9231b0f63379f27ec0d38af84d9f3e95963d1f79df5ac8bf5e08c04d716a2c66969b64615dca31bf5725490ad13ce37dca99fbeac02e347363e5a6600d3c01d8dd3a2234fd728b5bc870ea19308b80a0a90e4d116a7c25438e3e2ca6449dc8fc2e852ce7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hcfd9fad62fd8656ad253334a77a9428cc595e265541bd054c19b1e19fb64f58f6dcba8c1679a8b0d7ae4fc4cda0669ab9a9ba7d4caeb5fb6dc77f374f239e0fae7dfb7d9ff1bc30bdb7d3e89d9d876429409c16c220da239438a2ef6e1b79b827d002e5652b17b64bfd565cc0748bade6ee3f4e6d906f5a2c81a52a5ab5c98f28114f03868685083d1895a6eb8d92b37feffa57f4550e4fff5c0e6e8a35d0e376e3daf5e8a9490b2b18348f78214f6e3474d3c2c2b81ed4ae298595ef8e93c2dc1925fb48a9772ac87993ffb262be7683b7fe2bb38158f98432942753057618e1f1fccc54529ea6d9754b5e18a8806b644437e1b11f3ed4d15bfa80e08ae40eaccf49a2a4b69441d74b6b1dd9b97488465c4a2929775c87a2b7f11ff031900b9a432fcd44be34850520044df3eeb081d6fe705739bedbcfaeb4887990477c61d67613cf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfebcdb190d1c454caa9ef0c5503c20707e98969426375425569502242b6a435c5e910f461d87f19a1bcc088c8d7c0ca0bcf774294db43183885c51b74355eb8a2f1916e090671f269db3d10a9c4c1eab48e0aa3c9761ebbf3103decf84c8fa5b325c0077f092441261555b256431ae076c13d87107fa29a5873d02004532d9afc313ab931696d89b64179dbee29177f41baeb5e0957c46620ad07530b83770d4293f3e025e018454ff0b6bdaece7bd96e7552c6ff89915c2a6688300b13d7a19f5296104d77f570abaa5a216d2fa8f6334c3eac696493868c50e6bdcc75299f6aaaa6f6c0b68a4367efb51d9bae135f4fc7ea5dd6d301d97d0b98cf2860cfdb2f5707406eff8ca7d6ca3ca173ca318d0c3c87773b54b5aa59ea02d1f3117b07e794b0e1f1782a41af537706068ef8628e8bd9e35c15506f15a0e84b84591ac5e98e7e1f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdc98e467029d6d3dd8494f3fcf3dd66772907f9296cdd976b9707b379cd4fb3fc9368c6fa52e002943bb5b6daa56c7431f7f49712ae094851ef2f14fbbb24df4164a6fc74398bccf743a9586fc3151292b88d84574a6d007cdabe7c9997f1baf31fb00d0c916a3ff8ec2bdfdd84a22a04c0dbe3b041a8341aca7929aa521058ae288917b1d956ccaa7c5bc2006b69c67226c54321e37f4615184c3f98c7ea88c0808c68d44b2ca74ecaab7e698923016fd3d6255249af796d3bbe3b6b46f16fab29fb6ff3ddec21486ecb4ba89ccc0d32fa9ded99c58e4c9882b9bd888a1eb40d374dbd97a253d8a6f632ad4a01ec835b3792ce66487b49cae93c862770f3444dff7f253e544b68a1432b5a955ba8de970fa4a51ba28bdfeb51f21291a96690fab1fbf360194f41d6e0a155adecc72c563733ed01a93b42276105b5fa32d6c2accb2f1d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he9985c71b34633c8d02093686f49a152f61c10253b7eb32085484a00442761efb5d50a1accc2cfad071e2caf4ac2d74e4a5c141401437ba80775dd9cbdbac63bdb5caede864df317c4baefc6e0605b71f8473b8af6f9b1c7a23d53b5172f278093da11589e759a0d222862d1ae0aac8654412cc990ddc1537e70344312d8d433e46148853e4d9e3d4b9ab809df3d44f7fb5c79b67f66a6858f068cb719ca2dd9bf64ba2cf3b90bab136c3c03932ad4c7cbb2b9b6fba2b6b7d0f07ecf9df65d50fa861a8c091d47c14e149700b7909d5c00e96fa5fd1b41ab315d8450f8dcdb484dc2ceec68dee77874f1ead62318ae733826b4a3a1679742e975e5e6765c35441c32beab2961492f95d341d6f546d0dd974f59e097474851147eeb94e440132af1449bdfbde6ac6ef31e584dc25060ef24153e832718d5636835121d7e57477606e4dcd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8e39a40ec018a1d26041efd6a059cd6e815bd300bd9548396aa19e7d92adbe0bd7b3b31c4904e06a329f4f9c1b4dda9787e55d6f982ce783bd969f8f5411ad8790bf0a4b0eab3c04bc087d04ca30e4fcf77cef56ff7c83627b7b93c0b79a85755d01bb9873aa812719d7c525c3a0f446867d30f4fcfa8f91334297cfe8587b61fc5c855ac5f6b03e63cf148d7382f7b805dbb7debb8dd20f67bb2d0062ad10bd5213d8ce6f6d39500d09459ea776f29ea0352412b32ab3cbd48015c67240bf5902e20fe2b8d983022534f3a7814def43dac6905e3168ca038685e7212afaba658aef9f5d989eb7d558e2fde5503bcadedad1a19cf362e947573d80dcc41893ea8ce13989df53d7b02035541844189e4c9fada918a124a99b623003ef35715aa1788ceac562e3093bbd4ec9b90a1591472864eed8b8d1a0e2ff3a9f5be4f0664a7d4e14c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5dd1ebcf24ef9689d197ef991c88d3207b3263a7059aababf2364c1a9f89024837b6a3b25918694a95684719821406a536c680c645ad6c88ac5c20ad585256c3efa7d223e5327b08e347d879c23555837909cd7e939f2a7eea0d7b2440bf77e12e12be91750209d0c5e6ceaeb4cd117ecb36631be6d92c940c8963e0b3722f8ffd5e4529f31206bc7a40709f259587f9d877fb05dab5b9fb3c891f86eb1e23cee7bd15588d491abdbb8d61cd352f4e251673d26e273b2214899c1b77bd7b6fe506a0ec217d1a9603652b7d2b62744063587932c89c94765909c6e2935a83488f695c2606c838edd9fbacd22ff532d9f7489a5ea1b93221230eca2d55d5caf94ae0f60ec41cfe9fb2b06b79852025c9ce4c1098d1fa84284725fe9ab16587e54c9a528ea8e81c82a88770f8a422f61b57d6bbbb8209340fcd994c1471fb240d65b4a1461c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hade21dd58d3af441dfe437e5cf3fa460a54180b732cc5077b76de08909dc00135731a4b0975e399497fa38691b9ddcb90e0d6bb3e247f7c7ab84bc123b68cc989a6d46db3ac2059ac5e986d20c5782f0a4adb60abbbc88d8d78599f24a1edcc5625388199545b052c12ccd24727d68dcc162b023877fb2c3450f5c1402c31e54b24e689b4bbe5cf08cc5599deb40cce71e8e97db37e9ab2e8dec3e38965f24e6dba6736a931824e408b1acf0fa93b3687569a0cc1949bd9656510aba32dbe06066c74cc53ca2d3f98cb82ff395fc503502306c119433067a87f9a1b8eac9c093302f340e095b1f1b60fc797b14ffaff230bf9a47cef7c9ab6c97c31824457255e9d4fc0618d145b20e5570c92a8328f1c2a8fb8704f29f4ccb19722c826e1a109f0b30c9de01b8ed052bbe57127fcc9427563e5639c6d91c1c706e65e4ae8bed8b890af8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hed660d5ded979ce84b56dceef1d3ebf0c8c963282f1bd321f442d89826da780f45a55abc986a49148ddf9ce4f9922bf11c5a45d7e06c3c7bca23bac6161cd7be02d4f1584f052e47e8cff3b58a72d1d2d7960550e5ca0109645f59ee30cffcca671ec5dd1ae3fb56705f6f0686588bb563f6627e7e8bc6ede4a146e953dd511436e660514b972c113c847690f47f99ba42ffeb225864680e24f7dc021e6bd393608700f26405eb17eff4aa5833b493b2cd1644ae2fad0d73f21a529bf84aace72691dee4ce907f25378eff04e1718eddd5b2c49f0a403dea6d22cfc9b3d2613870096e4ed97b355b544fe5ca2cd785de15c1df0187329ea6b13d41082a831bde1394a8870df0e207e7ea92889c06512b836a881c12043d141ca98b3925d1809b6c56352e94aaeffd01ca6917218b9752b41d7fdb7d4eb3e46bbc5ba63a74cac4fea761b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6288f22caf2dba25918b986e9527c77fe07dd9e22e59eaa1b3aed53e611b3a943917fa17b6f9e60b33bfe5b7a7168181ddd02892bfb688f5f7652a352b1d3e734ed3e327fc38517e359528e87f1ec2f125d3d90d3426a99042628fc6eaeff82e02e0eedf07d9f0b4a634de1d9304d9c6f223e52166e7be313c97d3a771aa8ff0136dd96373a63751db7eaf8f06c3cbde148ac0b048a4c47a761f4ae899471f55e9a7edf61166939967d89426c065c42a04be3babb67f4ab5759e1c93cec04e70bb2ad02af109718f48558a981fa288a541939e05a73e961961fa3431c1504687ec2d8e005839079ba724c848a0fc112ddde05c9aa2eea58971e2456722a94916d519528c7047c231542777bd67c02a2fa67d0e41364b35c01cdb3010bce15ae8953b32706001ed925c3949800d70d217cb5c5f4e83b7206a85e3177f033b4822f89e74b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha1ca16b370039426c3e01e398b2c0727e131d673d87581df43af1790a91c1f3ddde66bb0ebf3ccdb1352c9e2918b9a6bf26e7d5d47675be553dbf6dda73364cf25bbf7997352c2747d6d336bfaf956fd12ef07bfc0bebe83dcfddacd8f6b6bd0548847a7190a0fc0dde719c642c6898fb93cdc675f669ad656ab6f1a73d52c4f950c7700cf607ed57d5398430a02f224c9130a5394a7b4775ef6c6d44fbe3555dd653713595aa145dd18d27e1d0ae4d8e80e601606bc095e49d4a01e44ea2fb3dd2ee897a03fbe7c646da7f0449c558e2099a1a8243f40b2ef217ad6e8a4ef6f373a34b1f37dff5f882c115c991096f6f6958968a01f873728f4021dbefafe97b69452f667e6d8e785814f0fb2d13287aa36625580ef0918498ecca60a7ef391383860d85c6c02675f6df2cfef2e8da3f2bc29c860812f8905b759e8d58d0b0ad72b2b27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h406a63c55e048abb3d5ef5cbbdccca1a683e2229a699892846dec3179cb076049b48bf172bf7c930eb6d13230a0a25812f1f3cf11bac274890dc6bedd73ebc1035f3e25a32bcc6fc2af1b2adfcf598382a84df20757c97561bc9ee16aeb2922ec0e1f008888588d28d6432502788ec19d92a4d1fbc0b0235cd5708ed58497a1483d467b6d2aae41922f6e30789bb02baad66c73e847689a340cc072e161367d4135e6d354ed70955830d09fe2afaafd2ebffe65bc1bbaaaf88d06d18fcadb13b0fb4008d0c2eaae05a09c80d9a8948cea49b4e652b1234442eff6a43713e2b144dc667ca3a2045a820959b60be5aff7e29101765de95c688cfe89e0edefede50043a051f10bef296fad841b99ef498420ecc18a54fbedf5ec44b583545a83423938567cfe9d1743a08947c67be6278fd59ebb0090c508c97f7dc7d4e428bbd5754db8ea6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6376dc20dac644bd3ce0f1bd25ce905e4e6889fc41ca52cdcbc26fd2bf21ef59dabb5772b85363f2d48eb8af370a0d34619cf6d68cfd5e605e33e7286c2bf28e2703f6e90429ffa35639754a58ae1ce19e166a3f0252530f658cae1bf0e9c2139669d67be87f16c29861a42d731c7f761cc9aeed4e87fa115a11cb836c27dd6f5eac5d3e8ddb2d0d95b39a135fe6bc3e07ae6fd9b9ec1ef58e41e0bcff90ee69b5b2de49d04bc37ff01d85ed6e9ce894c0d400ae3ea77026618b19b69b282c722a90dcaedcfac528e53390b8caaf75a7f58c4d78d1149fdf664d14cfee4b08bd7b09f92ed6a40735fb2fcfc69156df5f26c63624bc1bc975e58953f3bf035f532f1bf4573725c7471c997c8e7a6d7d73f64df05a822b4cd2824f4489f3fd33dcfa92b58ba1264b0c5cbeedf32447422fdb102918274a120009f668df195b56c0308653e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf736f403f0fd63899c2e6518f8ddf66497dbc21dd2292d416386caf10e094f3539503ca17221f29b9c9930ac80e34bf9278712c6af913c4fc3955cf3f85874e7f145b61628b81443121968b77c8a9065de364220493d5282e28fa45a625e2e72b5d10abc75add4bc8e31c774a4d50e0d275b349b4fca761cb873e3047d4f57f5887fd204dd0d1ca90fdf696b3c01743b2f5d986b17b4d75549945dc340446079f329c0d802794e1883e06b7a4115606f331e55fbfa092c428b09ff409af32643682f40c0365149d2ae4d93411068fe8ac7d8e0cf591518d7daed295fde73283dd631105c7049b3efd2529790422ea1c8ff37f3d50ef2bd2d081fab30661a6da710f84583dd70d176b763c4ec55e20e1175a45635e8e610b71d598d30c9260f60d52c217f1d7a97d2ad33911763a2bfbf07fc6922f7be05cba71a509d5a8cc52e86db2a0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb249857d38d3ca6b10edb5cac6835c20b45e71bf579f15d062f7cec100cf87fde7688e20fb76d859e5830a51ad24b745c9b33dcde56cd834fdee099ef1e0a5db599031ee1b36d20517a991a9fb9107beb65f102f61c0b1325d832a59d2eea4cabcdc6d5e0eb82bbfb50f5d74aa2bd104393b3e4ed2b94e22c96eb1045f966e18246107260e9804bbcc5c5f326c8c58542dab15f257532bb0a78b94ae92eb0dde0044450d9c742102e4fd706416cfa5961a562befe7ec88b8ab0af9d4ffa30ef67eccec4248ec5fb67f83fdf932911fa38cf9f8fad8092d53f9823b5125e32c1a979a95a5374b38fbf41a32395a7794e8d4786a4041716f24a73467b88d0477bed14e03e44d8453c89d8c9167641b064f908a8e983814afe7f81b2d9aad5065c80e658cde273df017e727cf185b3abbbc32360bb09acac11919cd442c4de487a1eb085339;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha9e4a8144baa374dee4292c156f0b8339afc6bf1633228499a3ac680a6840b5764f3928ca2df27b2e112abfc4eae0581cb34dee8bd8c2a8c6bff6ec67ccffacc8e6e1c90ab5654529ce71e4975cdde0db2af7bb47309044470b084a2bf8b6d6176fa8e870a46904cf4b2f2d22cf4a0e9732a4b3f7299e7a103b6e296943707035a2de9ce6f1889f0cc0d653876d6fa47240f3dd004a2db8a37351cd558b5891a92c78d337419023aec7c268b533b97d36b8f6642dee7b40bee24b48f8be1c7ef26f93b9bbdeac9a8a86dc7bbd458f61daa5f3f71a4b08a3ec2bca6139f0a44b8387fb18a136fcf7c04cec42f9e9954e9b695e1df48cc63862a3201ac7562fd00b902f5815f7cae0cc622f3f2d514d58e361b39a330d0efe4eee59f604811019a23246ceaa71221b9e01e6dc73453ca497f4ee659dcaaa6f5c610757bca0347930e99b5ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'heb7d7345be045dba0cb258795c371cf3c2c8e134b832c987fc242c8e8cf7d85bc5e9cbe31c852f8d404b256adfda38bc8225fd64fa23a3438bd70fa3c4941b1b90d295e06eff78607a8ef482be89dd8f28f5140afb429329adfe862d7e490e9a1376d8a038374a1fcdae4e2edef8d347555194b2518eef95749f336f8d5a0bb084a5d9ac1fbbe8f227bd39fa5aaca080190fcc009731ee9c8ab0eefc3cc540bee2418c05b58363764cb519cf313b19c16fbddcaabbdbc30d77f035c336b5ea35083a42db009bdc6f3a51d5fa4ce4c4e8bddd89965ca791cc19905b0efc03ab50c0dc1ac9287d60d883ca83fc3e51af62b97d7fa9f88708c57618a2a6214607f4cb45068da3aea8563cd39e0a5ce9cb6602bfe0b242919e2ac1afce4cc1ea42b892b34947981d191fe7b89cd47d5700be87fe42849ed40cde2e32def8874890deda00d342;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h801c98e2f3d2d0df4f4fb43688b1184a758f3fd9b1a26dd7b2458dcf7dd87ea907e829c27dd208eb10ab8226525ad29949a9632ff097eb96e349bc4a8a52f65bdaeef4f661d4a1f22b146148d2be132588b5e60479856b831ff9dca5f56f770f2c1e52c448551bf64b3fc31b7632b712ad14e41bc459eac343f92e525078c4ae9618fd12bc4ef15d25a201d8cf0d72ca749d933fa4b044eff84204b8729c2da9aa85d62f42d7989ce6de710eaf2e9f3475a96705f0fd5d90f75288262e2d58652b0f6406ec9d4e88a6ae29f8cd8f980dd8bd91fc66e005deb89c7191f6ed0ed44c6bcba5308669c0ad2537504ac25768e2ab5a0e02579c2e18f61df8b5e4de9b370574c07bda64b3294581f2cadfa2ed76daff478bf3218c44dfebfb70d1740df869b48e5a5b45b1548ef4af3323172827da0241d657394d14a65d28447afdc7936e7c32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h320b64a115b731342228b53d7933c6d95bfb334aa47d7293983fb7f9740d5e8c21df88610e69042e2c9bc844a7d3f6e1bff9d3a94c6b6a1bd623295c15ef535da3b2b1f499e799b984bd441b85037d1e6f3c2931c02989b4fdbc9822042428faf5089d9250cf34a0d0c7fa358768269adccf91703570ea793cefa142b19d8062aba6e585cdb4149762c572d0f975ba9a79fa46fba950e87b39a86b3da0f05dda597746b8ab4a42f1b715c63a2026c1e9fee511c23056831332202ac7c89f167834f73e1753bea4dfaf06b14bf00484467d743cff2b17e397111e040f698b0100f4978a54415157b0bc8b7538ef7fa01cc39139a7a3ed41faa53f21c9cc439814973e065f5a1ba076896ecf45bb6185f9e46b3ab407121dba9ded943b1df4b606f482cea361546425f9485c1dc2aaed1d9b42ac900e75a1d575b17e12c7c51fed8796d6c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h78f019549543d65674cdb1bcea9836508ef5f191c14dfa8ed59c2d53c58b5c09483b3a496a470bfbf942ad8eab5973f23b14ada513f7137e01aed27d9a7d1b98e2d37077d138f3f78e079ee26dd56bfc5520fa1d56818af14163818c53fa6ea1415024edb0f7d3b1ffee124d59e3f7599e05ee6fe27bd9de32531ed66bbc66d2441e7d1cb6b88dcf5318e917433ff0eaa01c9d1889941b59ac04a1bea9ac172b55fc0ae1fb16b4ea1a7b45d471bce0839311fa9920426f8c0827ef87169053394c3cece81fb88faaf4d69afe7d9ec84a7caaed526fbb0c6e1b26b4c35d582fc9a3f297d498def313f68f42641b9cf2e0085dd0469ca8b5c814448cd833ffffd58d387a42358fafc36e7b4f81dc88bdec770f48b83a3a7eac72c64d52342cf105e45172438530cee1e4648b86217b2784bea3bc3d3f27e6faf8d7b6a25e0d6a7e6e9bf04d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h57e38fd0c6d7b00795a6ab48466fbce03d3fba9fb501477f36defba403bdab9e67496f7eb91a045b2ba659b32b5c5d8042a681bb7092ff38bcaf6b23b275539b6f51217d80ebdf0cc7b8114e967dc15296d3756d809fffd02d040522438be2560e4f33de573ca5f45d4b48b2be2cb0a4c6043817ca3c49dbd6ad8ed4416e8545ac417aeb63721e8e21c345b0c9adaf9a58320e74cfbb7dbcc25eb2f757a6318c3a6da6325561e84322bf0b4b6ab3ca405a422118649b6e0078b69162c9e7aec5edf3cf9a41a05c38365604b898cc68900654f61b66d1b706e93731590acc4ab16add3455ac0cb2016a8346f1b36f9e867adfd22fe28cc0dd3faed916b5d2e4601ad79787a00161c5736ace1c9fc2b7145a96539dbd78e063c3cc1b5b973b5176e17d4f85535fe66f26a6db2b67b2fd3063060f0ab12335320e02e5cfbacc39c7ce12e402;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3dc6bbb29b9334713cc3acd514a5a245a0b4b7ea38dbe85a02631d87c07efb76cd40634db814979505a2f3eb18c79b5a42bf9fa672af17e778bd4679f55b5d2893fd512b5476834b2c2f247fd908387a3bdb3f47edc995a012d9e525afbec1c33b636c2a7f07019e8581f4019d2d6e511ff11d67c6eecd668081f4350f5ad10d678e24488b499c02d74583de1206d7c7567ae4329c007c12040e597fb84c87d3dc7f45c552738c53999de8f708c1e2d7f6f759666d183a09260f555ec0557501c1f39ec093fd474c7dfe5cdaca3ed252d9e78ad12eae3053dfc324ac8b94d07bade05946cd68b171aadffbd8e33a1aad29ce3d7443d097ab68efa26269554e485a5a52222cde11580578557ff9a64cd590fc0571e482c60cef622e4ec589603c1db3040fd0e8571e096b05d8ba74610dcae1c3f981acd9730ec3505332cc1734a994593f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h75b297156b01ea434927e2c72009425a4c7cbb919ef1a58ed227158df6e4d59943cce50e5d20d1658b9dac38acb8f9d7ed1903ed24583a8e37acba6105fb08faf1966afc3a872dad06633c0b3086960e33c46b846b9a4214b27a88046c0b95aea89e4edd2a6ee29550f46879427a2b4fffbdadce46027560af46b049f1797a64261593f18b0734c88ad91e9a69fd99c37165cbca5bfb0772c42d1991b3e1573cdc0f3d4e2a7bcf56b72d8bf9a54ad07ab28e849b2d232050806c0c795d48d78319446a357a6feb4e0644861417d5ebaefc8376e6387ff62893b703c788bc32ff9ccdf8fa0e0ad65de774f9dc41da2d7c8851f922844486fbd10765245be60d3ce6b370bd3fff61364db9003b07b209687f19d2a1477866711a5b78b037302842510aec85ef984d09010d2c0a27966750bb214a726e44f64d3bc741a9042f00845e8e0261;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h561793f6a4894b1ab5bf61b09c13922d798a818b5bb956ee22f48f17ed57ac61a43f6d23bdd2b4f7ac360ffd027c2c92ede0fe0f6dda3554f5c028d79e266976f3d62d12dc7635c5f487564f959e5344480d80c1aea9435c0cde60968006fadd81d263d16165018462cf0cf33ac038abeda3555b2b23eeca453c8b474de010b3df62d06a538ba5c6a74f24912670b2eafe698ba21e90d5a1319f85a4c27dd3ee7bf4d50f99271fe507cbba7e24b22c28e851fa31eff309629ce0c3db1349e739681f16942ff5b599f3ab36fcbeea6d490b70432d33d96cfea5dac414fbec02c68afe1babddad11eefc709cc20d6acc6e86aba555e86ddac7d4f1bbd175600473bceaa339fa83751092666c02771c736aedcde53b6a324135331f0e00861240125bc531b7c3779f1ca13add670c17e838350b9e9662cccace5a7529f3d54bba8d3116d29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb0be3153fbd596eaca1ffcad971b4004e5221109d8cc49ed9e26f65e11f5f406f3ee60da791862a809b9eb6b53550008b7dca9bcf6641d33f14c52407314bd370648ddd98b7326fb938248369f68ea90b0a63ac8b9acac5517e8606f5852e00f1f43b27bc0b4f842b3192232ebb8d824a6cab1a17e90a457d88d5f1354e5b4daad597b9ab69340d499759ac64f49b9a1d492f58740d622cb6f2dadf9e7b5c7f9c029ad413e5ee24f0f90968084ec315759c9dd8cfadd4777c05b488e66c32b2672de2b1562c533550d50c8613513d287237efdd17af56dcdea779cf6f6b943a135d866602059064fcec58e19f792c2a888b8a3324294f95e36c3bb554845bf9f9416ef0701e8b17e35361a278468c8e796545bebb5330009da97ef0b4ac98e2ad30e08f00965bd5774e7e0a25fd858427884bb60fbed771b5b954e840f772e9b371a7ad6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb8d35337f117b1273672ef2f68bdce4382f1fdf2dca6c5cee2308ff586f7672d0895bd1f8be3e58af3f514b696105601ec0947a22b55cab28845479456e70922943829c73256bd9391bbbe59878ec6f70c122a79e9ad503511bf993304592402050e9bf421b3de72db3ebceff42886dc456fe244c8bebfcce0d10ff306feaac0059048d5b0aaff2f127696433c2893a73e7dd4d250700aca93351d3b15090ae19c6842eaf4a06b3f5f9e31445191d0f75b07bb4e13e715e33d189f90b20b9f528dcc0696f6cdcffddb4c63affab8f19a0ef3c97f18119b29ac963e6e5293f4bdbb9aa7a15a1344ff4f967b7e8091def0cddcd950e8ad9acbc1bd94b213841e91f4bf95d87a08a30104a47e27a7a79e635d74da8acd69b76d1ed332f02eb7dfb7641e15a7d9310b2be8186e2720cc22489e996791b5c29048315828d7ada7f3ad01445c4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3d9932971060071e4815fea14d1da4cbfe1ec58743467cce03fbb46c57d01f34bb68f2896c101cb25baaac89ae30bdcda22badbafe8cbc01b0e2555d3ec1e6d1bd5cc3aa97f6f81bae43407507e12b3d51eff0ae64e89031d7d6fb417ed76afb95381964c48b0b7ba2298cae085bee2921fe8d94e3de5f159a4ca8df1f22d4ebcb04c1167804ee635c2ec5a74a8ce40cc1bea929a543c92ceaddaad2fcd5bc9f358dfa7859713c0dd1244ff7e05818e046685513fc2e4a3f93afabd474c2c67d3c1c8697cba77ebd92c55651d4a863f45a6311a834413477a77233433a32f18892bca88be3312c4f01bcf11ea1bade6d81ebd7cac292c8f9ce237ae5177de8f200c13107adfaf632c07102f01cd0fabe93565c6b1ab4eccb70a16f6e0ae27d09d1b1663dace456c6c87e830837081506cd13d9ee890f4854a5e19beb29d163d62f49cbe0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hade11abd6f7b22a3edf4045a12f6b9269a97465ee712bb2960f51b42f25d70d2685b9f34b6c325eeffd92fcd486d4cd5263a29b4b636e82f9dd108e9be130f81dbcaa968e98d37b7a071b8bb93af5a1eb23712ad1e26dd8f3dd2284c4c236593df4db3b4ed37837e046819a79bc08cae6245f21cb468703c1f80b6b5bb681f291988416438585533947a6c1155514f5010bf0e891de3805f480e423192bab45fb126c8bb1a2545af4eaac8c48bf120c4d5672f6ea4a350216582bb5681fdc6f696191aec14ab65dc8eb57b576eff866a0f34038f5f815659fa021563e15643055e5ba2e874cc4fbc604b4c8270d6db1a9497d42842b17196b52723110e16a7fad9f78982d66437bf192cd76b904bcd507463932f3796f4b050cb6a4aa57ae1312da74f814ffe5042cab87c88d4f089c4f2d8a8db1a653c72ed9c40ce370fd16f2fa20fa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf8c40c9f48d1c91412905d8849dccb27831fe33e865c92a14250ecaccca6cee115491222a7165bcac0e1c84486d7baecf5f796b3ddfdf646efe12a6599871232fc0e2b7f26377481c99f9d3dc664eb0b356f1126c611df8e5d062f69ef8ab99950e43f275b9f2a77c7e4b1ae18e160f87d0a641a196d97065f8e75792114686240897ba24d77e76f87f2984d7a7386003b784558a9e29ebcb3e7eec463156aef012160476646bea4027f433275ee5115dee91365a34f12f27654bc345e5dbd06d4311ebbab1187d9b41ee54f59eabf6c5f0bd57d26a2017a926c974d3fa4f0c0cc5346e835225817abc1ccc042f8245ff983ea7c1543ffc9b13a8ee887f11c25f84359826adb42f8a9ea33ee3c19cc85b3a26c661e8fc6445164dcdb1adc72fcf60a044102403724fc43e58ecdbf69cb4f12564fd50ccd5af8ddb6b1c17a4a18105387f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he8119cd77d340a679709ac527f5f823fc7902488f32c88a8b8bb4777a1ee3790de5028f0923158f4e28c2d2195a05596daee561922db6479a0d897214d2456c276ccdda306539458cd686de269f9f2deca55d79907c19b71f462ff1141a38ab04dfcc6d159e1d8d3c5e76a42c3392c47117061d91138bc3a37d5b3ee5f712f99231be3d45d6ccd1b631286eba95f30cd6def59a77baea4041ab35eccb3104e6df68f1968c45b83a1245524780a39f178ee98fcabe5466925068b8c9b15c41676f8d78938364224f4911befb820862bbda11a195f739ee1108a49bd8fa38957210ef2d171e271942e57b65396eb92ab97e9a4d3a33a55f5b222b101b2d04ee591300401813c94414a492c937dde3f7c68dcbf5a39b057f3e29f8fe5028c7d72d07fd1c70fbe35825e043c2bf436ba72f54d20477a7549b9ace1348c639d8f6527b8b1c820;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdcdcc67caaef4d1cc8f4d1e6a2c008b62453ded425dabdec15366b3ecf237229c1ad785761d9d3264cded63f1cc8d1048cfe77a8a2372ab63e5fb7ac0cd629b4077208ef5ff696c2bb86b947be5d2127b28e82b368cd6ff9a681c9cdde12cdd4e3c5467837b7d606233a43cd91c3f4ba79cd9f2645d4acce8b2371d038ece2b093a46b05aa96895970916d18c6f252b6e6e6b678c4dfc33285f191ea467a08ed0e73db364a388fdfc40d3a74e74448a29a23a38ddd3e70e9c57df2ce71bfab64383fd270467151835788de4d0dfdfcb7ee9396970c1cdf718a2881daf01df40e104b0170e864998a0f7d91af749438f09fdcd5ef4864cb72375e99323ff23052e601f8843c16e03f147487812ab62daedff9b29889bf45429886afee14c110b0224fa15c29810ecd99cab1a26dcb28c1cc1ac7e1914d17ba07414c67d78880b35a2ccbe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he2618c59d7c1ee7599fd101c1c2f696ed57f784c05df878cb184d36b5045834a8ba20860a1f103f7ee660a41d373295d0c7a5412164f3a8911768b35acbd4331d031d980c019d72b4760f8e4485ede2c9374783163b99cd838263e83aedd84c8e84f1445a71f0c2621c558c6369e29f9c17dde34d7414e797746643e2925d42abaec8c5ae572d373ac7ebeaae9c20783c829efb701a1b094a551862ff4b9d364335ea1503aa4cbe613547300d1b80c782db6f91207aeabacbd1eb3506e734f2d8a1fcfed42a21a046aae06f691a62be69be967ec799242f32330d4d863977e87df526374c4c7c90a2c82de1a7cac2f7c67dc94e1fe2556c0a4e92fbe25d34dbc1c5f8f31fa52be69a482b371f76baeaecd9bd1ce8b1137a2c88f712e10c03adcdba4e97a80ce8e785d0f6d067d7084bd42fa13357fb53692a0f2a0236a19fc6148a3bc22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6cafd0cbbe6bb7b7d319fb33aa970b68616855611f3a2cf12d9d8a31bab883cc6ff452fb91351766e8380462724cc37fbaf8facb37061496e3b80876f5bb4d44815479703960a4defb7f317cf8c9d77d6df1de1dadd5c6eab2b27d4166fee2b13f0b116c5dfe279877130739c5dbe966dbfe1166698fd26693cd9f5eb5ac2d2a371bf562d3fd88a61ae63d067cdbf9714bd838856483d38c5823d9d95f34594bf9747710590f177743e0c3d1a5a9ee23a75d5363b9f6b8c10207074f25205f36942e6b318d6e849acf5f646ac8e9d91710a137ad10d2672e8026268da59475a88145ec99cb636d5aa660cc0d1383adf975753602c176f7b633ee53fccb4f6ed504cc085467afd8a0f3a46d0d6fae4df7d9523eba97321993506e4600b98ab15f3f61d4422c1fa54cf248f7d425efe036fd2030efe8cb571dcaec79de2fcf89c111d9df76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6faac4c3d18173ba8299e668216143311eb94b3566d7aa9fa7324b91fbec628ad9c4e3891d50d675e5479905855930b6baae95fc1a46275296d9521fa470a20ec6fed735eebfbbb794075983bfa9d7a9e56b98808f4002d62ac6e1909ec1952e0e019063ad1a79398134feaf2b8efe3255df954bd47411520c6c19b1390538b75c55e1b31d9ca5e9aaec6b558309ca76fc075d6aa30dede13298f86a593c0184316c43247436780b4866b408aa15f95be01ee998f80702d726af52ec95b41bfbff3ba1e2d38341cc3e1b96aa48c961c698f359ccaddf218bff18ea247c3543fe03bece508e052427f126297553cf72416b33410b43e967466a62d071e0acf605aeb85d0c7f90d3948bc2d1a44fe05a5b1d9ed8da37472cd6067f1d690d91819e65ef66eaeefed9e76794c921ae285f9531d3215295ccbcfa0ee69a7b7cbfedd6dad036de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5346f6a9d47078d03c3f50315cfcd4290841b57163a67917955cafe1fd7621fb5e8b90cc045a589aa96a30a0e41deac86030a8f7259e86039e852c4c142a515b7284662f452f6849f680fff23784710f78d15b5976b5ca572a3ffef883e18fb3525129431a1e1055e738ffcd860120c70fe19ce7124a17185cf3cf7b63248d8bc81c9119c2cf0181ed32408f75621357b256871d9a4e818c908ecbb6aebe40000da22972e137366eae6cd8b5a1675476b309c005dcf55d262bb0f884bf4a14cb7f634c9352ae23c7d3dc52f84085239373aaddd6fbd2b484fb4dde0133e618c48cacd3daac957a887ca43cd5892e7d738fa25f59773aa9f53c1b99c662e794b74696151aa370be292985fddf77f5edd3e5cece4f110473d0b566bd8f3c59d8ae430820f32cedab2ab3e81324eb67600b850ed82078ad94481e0d2666ccae87ad032151a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h744aa30ecd47d4c24686afa246a90c0f7a0b91e0240f8b0f9da2a512d398119cd58eae0d69d544de297116af95b75cf4d3156d5e8d1032e13c161f93480b633187d729c68c08c9cf9d975841a440d306ce1fec92281b46bd347e6dd14bd0d5f49ab077e76b7dfdcddfe715eebfd66399a0c8afb7cfa9eca5cc77ea95c4faa973830731d15f7e7f1ff88b19b21d58422d3423036220e963b8491de0f0bc4c64855f1689ae37add38ee6535e0f198ef96c2309943d980f472e9b67090522c69739a5e269f148779f719ab75fc417d2cacc80c21d2a80e2a3e934b028038073affbf9838474d27842f9fb13e3bf0c643cb46fb479445325a8643987282b2e46bf3934ffe618044ec62d1771b2d4f216707a808c1736c08fdfd8659b5aa5c4ba30eafb6e06cb8c7ce1fe6791833905be7433d709fea60f87876bd2e336e9f74b0dde18fb02d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h92609592102332ce8f1d1ff9a8ca5ea72f4a37e65236b5507e249fe864d3130d6a7b6bab11557bd6509e41ad0bac1b2ed4d5c2a334afee0ca73fd8bd8ff88885fba70180c096da69a247fe5a46ed527a3ed8d497e0e7b8375b4e76afd6f1b89e78ab44baf94f95a1879bc71e73b47fc2e08eb24873aa1dbe060d5825bfe3686dcb739e744058860b67337d824e8006dde4c581959aed7bfdd2ce3002c77ae198b41c21853d969e115dbc9c389ad9c81e62accdc632699de3315d747b5b9660ffb3478fce46cd596f485826de5141785fe65f588b35eaec495cdfaa3746becb9140ca8b2a99f86f3c393fb11a12136be9006ce630d5a84481830b99afd1ec4c2a33a483dbbbbe09d57b1d1afbd9f73529ae2ade059ff9bd41704fe3f78aba8573142b89b9946b456778e4c79e087cf33afffe28ff8db2458317483cb44ccf48ac3aff8c3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3697fdc8e46fd17df5c5c3c1cdb408f1e8a190c1301bf823b15f6bf8e38c581f9522a50244bb37cf5e2ebcda972a2297b8451b1fd58ed3c3d1ccd7b06ca43d104037e69ce7a0ef9df233f15fa0b3f1ed6f54d74a9d0c5bae0f5aa3b0488d2a2584f1fea12c0682457a681dc98f66ba65c3506042c4efcd2c0a7b909d4d253e5d4dd7eb1c1d635c1f2bd5e08818a3a868ecee9df1a5d31647ff844b828e0c342478cea2c3d5b45885dd7a339feeb2b41e3b7482bb6040f525d349fa8937a6bde18fe05585262d5f99d31ab895b231c572e716cdcd2b72f413ed636d4afe94b00aec4d328fc44befa87484bac8c50eccb3661f30e3f66225399e1e8d26e4ceee94d362c7f0d1a411ceb293fd529f3b064080d9e71c9c0de71d0ac80096ce8bafc0cc883fb1506870bd133481db3792d30edb3a1a8ada7eb91960e89c0e8abe64c44347780b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc5b4baaa749dc2ca6ffff83ffe5d2d1a7e3871ed057933e9950ad80d88d06206845eb9d08a3de9a22668f63e5c11e7c9d4a512d290554e215208c9b3b4e3d2c6d0a6c0c72134732a4fcf17f6ec8096104d69d57120efb1e37ef718352696a24703afb0b970360dd8a09f715af7b72f4e3f56d1a3d8accfde3e59e0520724789b36a2e651a195fc75794ac9221d55aa85222fdbb45f648080cdcdcc12081f05b40388ab9127366c722efda7e9c2800398456f2d852e43a707dc2faf1b3e1e5490d7d0ff4a7d1b911302148d591ced7a38f944882ba980122937f3cb6d56fecaa07e72eac279500f4f0c4e773e3ccb521acd2b4393846a08641ebdbba5a5d9066ee9698d2d7fc100748ad66d0421ea23584ce498cfc3f570c9cf42155519a53ca5ffd5d60a50240fd7db558ebaf46ff91a0a98ac969336b30e66ea034a6a2661983aa9a39c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h80ac42d7c8056e26f0d62bb7c22669cbe129e49c4490b0e35290a0eee1f309cd2e75a43efa948dffc9217699e2e9c150560418bd09c7c8240e36f56e05e1183c50c21dbfeba4d5b7a0df33de62566398065935cf5f701ca9490d9ee9ccfc79ae3016438285c2bb83bad8f87ce0efec6608efe5feae3d9ce9e2f2d4fc825a91091b8e7c482240fe36b2cb85ed8b351a0a00b3e2dd53fab5f1b7f92a6344531b122f804cdf8da055e8bc79a2eca732633f91db7f747c3bd19de1e8ce3d6e45b72716fc05e2ffba358d8818a19fcb9a008f8aee7847f052fc378bf6b3ca219b785bdcd096bd6d868ee172a50d593ccc5440abcdd5afdf61a4d8e4b2f463997703acc309d209023eaa70359edef3de58cdfe0c4e93951a0c6ef775b7db738485de12e51c835191b1165ac57c98627f45f3815e2817ee2fed99a1feeffb3debf800b6c70d7ae3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hae0f462d4aceb7039a60190c00be620045ad6371e00e771c8c93444e8c0861bfefd6e0af8b2d7283dbba9be5a9a57557f89159b1f292bcbdf7ae6daf5144013e0b0cfaa1fab9d08ec1a1b2e45252072e45d1869ae6a3baf36294a4e5fbae75137b591ebbb04bd49b304e204f25478d6a349fd63760097ae1d23b9d59ba421e232ebd510635dc8a817a5a5f2da19603aecdaac06928a8b9652d710add27e89d4bbf39ca71a2fe1073fd86d932325445cc4ea8a1fb925d793a1135b597817eeafb4a2a6b713cb1149f41d3ea48e4327bad8ad2dcd6c908817e58a5e7ad77bd670b31905813f6d347a90382ed4897dc7d64a3f3e0623af55e8370ae09646e50491656b84e4ebbab245e1053e3dd19dce80e5f2274bc7845afb4aefe9051292ec434b8182721f417049f89d2ddda1042a2fa0558d5ad035f0a38fd0654b23aec4c8fe13483a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1ab476fe95adb9b98a38ec1fbd0f55c3083d6c807f2bfc91840df984bbf46c3dc4ad14b353932f193ef1c31fe8e11123b00e5c36bd81d913b861b5fe6043dfecbad06044a04522f4e3255c45d0c36299057d6470aa5b46b9346e699ae6e95470e9bef80e44b2535523175baadb36735e0e05797ee755d1edfc35883c267f8e48952f1458f1f2d88bc341e60b65390350684caead668dfed3e5f6871ccca442f19e58e4b98ad0142ce5a8f22285313c0f28b8cbdb94cd2ff10e8adba4ba431f706c063d845beb7a3173a8b2301becf6dcda7ad9cbceec59b51de9264d9c6cd5819d9845b723c7aecbffab41a4f38f34d0cd8e8a2885454c91dbc2e1708f7692f1ba8ace784197a6a80b1c6888979625c26deec88e8ed497bf68e4fdf2822bc514dadd16717643623b4c0e2bd98894230a99a5c8a7dfecfd09de4619ad894f7b88f4723d18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h384c4d554097c311193cbb8a5b4dee68814c0c101e1ce6337cd37438ccbf2e828bdfab245273270c0eb49a92ed2fafbdfc6e770b250eec417106053f9a87aee6ef03599005af6af75480014310bd1e20071cc2c3ee0af55b0fed0bf1ea4f9eeec02a196d41da5f8f0c26b51e606521388645659f93bac2fa4c9f9ea910987a8a14a9485983733342d09b05f96f8a5cba136b6d6f011e0f6866840357f1216c8f595f3d16fbfa4bfa7a8aa9075eb51af557a4df3f59d8e83e1e367b51bab2b81bb5f95d5d6238d98bc089df93e9d7549befe8fefe42f408364e5197a5ec975a5a983d3f54409f01a20153a95b94901505e80583421ca9e7e5b9cffdcfc9f56c8a3eb9e2e30b988614666b0ff76239b3cffc3cbcb688754108c4e94e5a690a43d7130c6545e53fc96dc19d9d8576378d2239f1af9425df3e823c3e326846855eb321f00a41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1a544c3210ef1968ff31922ee2f04960eb90853bc5f0fe4ef580da0778fba3ec60730c8ebc47504338afd680f83c876bd38fd49a13e80b3cc0970e11bc484785c8efd573a2de5c67cd2f7f9465b3d8d073ad4c65f28b7e2c8b8c7f8756a734815555c3c65277c5b8386c6308ca26298ee48afb000f645b932d814c87eb0f6ce11e8d7593063438e63c023be23776f5747f4a9f05ac4cecf4cf6df6e30b838bf52251557d66790cee1aa1e6cca3a64e8362a8b8da19d7040a4ba2386055cbada2df9514b4171c1e55c5a37da5dea9839edcae93e606ab5df069d3300fc891335fb6a35b7ecd81a5c04a094f9baf8e1ef23b44b243e6a0c729e287bb5073f3021f3fc276610df55f8708b30867099dc0b931850ffde04c0dc09d384f5be7176baf2d5c221c03e64c99776aa181ec307dd8982276b6b6dec73f9fba4159b5ca773056d875bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h517061f4110291a5ed590ccf7459faa324b75535a9642a1d0341e746b109426675a5914aea20a5e7c37cbf75cded979bf1b163426497cba6c121aa252954f860f2f6f57ca8299af46db36e8b0f05ff58ce5b92c0d3d764e818a199fe23dcb05a705cb5d39a9021c1dadfe325b08528ab8dabcbffc7bf435032b7f46b5e500021613b04b7497c2a8ff9a37b4d2850833eb4ceb27e5d4577d265cb007eda4a81402d00ed6f963e03bb50bb5f17115eb172c5e5d2e53d8115b82b7e4ad4cfe4c37d68a329df7dc7d087219786862a60446001a449ce97612ff66134db3bce414ca4362cfe11e5ddd096d4032048cfa8ec64539ba6b4cc0be9e63fe86a52aceaae46390be27d02bc0aa1beea137a575fa947cbf4b1fcf4e78a44552ffd32790b730639f5031291136583cce4f9095e678d3c8d8ea0392e6c5b5d77fbde177d607c46d28a07cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd3c61061c4ac0e072bd745df2215ba8aa38f5a1e16e4ccb47f6126977d51a8e673198f99b7c5fb614d8b4932620ff65449058c79aa9a9bfb86cfecf4ffd775dc3df43432cb94185254075f0d99194b365380089b42ddee70802884faeb59a27e387e61348ec72a8072d50513a441ec84958d9471b42082b16a1978bf3feca9fe1bf03f31d08024a97efbf798ef97b4968a2b8a28d417c28d85521715fe4cb7def214a06ffaef2c2462fa5e00f57d032e9666b8064db1a292cb7575d7094ca36bcd386e009cab3ccceb8fda569e53865aa7a98a5bda8085cdabba2e3c5a163721d1684a752b52e7459a345818c533a33d9fd48c89f66c483f7e290672cd831bef9a491d422507cfaa234ae2461b75e342dd7290e3d90967559166e97e0cc80b02c999d85d602f17d5f3503d6832ee785682630f5284c5b7e94f6e7ed6cac4788a3f7bad8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd779c6f70c27351d2fdd3c0d3f91761eeebc41dbb9349faadeef05ea0b380756faf250cd15382c6a456faa69f1f6145a8a9a905dae3f16ca479fc1bea209b75464bf36eabc00df488646d0611c4d80f84da0a3fd9d1df9417cba0f8fb12bcb8b47c295fd7c205f22e5d5130d0ab2db7a4ce8cae3a34a09f4b61235edc743669e900fd507580bdd16441432fd6a8345fce7539895fd05c7ab5d74578df61c6d07e5ea22d626a8eda447a6d38114e69a78a082ec2b2dad6a2ec8c097dae4fb6a7ed662a98c15cb97117fb3f1e50270eb30a7c8a93be4b2a97ac859096c4e7954c03c29b2d8b91d9f1abeff33aab19fe95312b7a6c0416bbd154f84fa638810d8fb1b26afcd009e2c5084a10f719732e97d609a9b02bb4bf856604a5543cd915487a426a432b3ee1f5e74497b8f80a13c7258be9ffffb758d25b829662a6fe2e8f420d7adcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h78e2195f9a415e67bb00771d837ba15751f71add4016059be616abee000c337a365e0f3d30db0bb6e7397042043d0f41b016ff28ef10f4f7b74940e4fc486f0233d3c8aa738e2464b93b343cc427e9cb053e298863145d0b267cb8e31e20c13f20ae396fa76274c05cd881a1543e52767baa52f2f8f1d5520d453902059981e8d4a1bc3f8147e1ae9965f6f7451aa315ac8409bb261f5acc4274769d4510d1b4a80466d0f0c849ecb4a9c78c86493c4b6f504466263d4bada0a4b1ad4628559b9f898b08bbf1e419a9a57d9290de4772965ef1819fd30fef6d807652a6521a74275d66b0301a4602ec1c5114ab9cf97a75c4c7f0d3143595bb9faff7cbd9ace4fe04a80aefb952ccd44a798268616d07a7a8f07334130cba16fffab397bca12fd9692d7f5c6a424933f38499bc57449dc621f40ed7ddc0ecfc9667f4e8a8e9c8953b6fee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfb0c8e4c7a47f8eb018e5a5a81cbbf99538cba40de81e87f588eb09ff4d0bfec890c18e8289541f6a1432ba2a7f056cab646f553ec5166610089b0337f9ecefee61656007e49809cb9440179668f44a4c511a82e12b3e145ed53f56ccf957a77a83af9de1b4a64dbd594982817983ef28c8c3cb0d964182e1abd11cbcb8f39f3c62fc9225bfdb3a699c8e701fadf26c90a9b0e6abd4116da594bb7306181cde7fbde841871360adc37b10bbae4b6e3818a4de8daa084fd3ece6d96ff13ed05759ca937cb19a88cbc32444397e9f294c990c1e6b2b70e30fd26e75fb38cdd927aede38abb925a19f5c9c2ff4d1225e33711d32ea8b5e91a6dd79f0b8f9e82117b7bf9af6bc42ffeece84724afed838a828ea6be75d9a6f7753fe972659aa3e8ac098f4a3af2c1bf160c88a75b5ce8a204b4a97a5650527db93f9bf4055ef8dee26d3b10db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h67ec731bf65e135d5463d8e12e5a03252ccb59bbe3c43d19b67955df75a2a0a53eb8d436fe826ded87f273e7862fd387f69b6648200df280d906990d6107caf1f3c25c49054d7b8d7c9e110372828b251162c779cb89df34a664feee2892cfdefded1bd73a76823253ac61d50e75067ef437fd2a036899f287f33eabb991f910adf441ee20a80f5fa755cc2f469b21d9be5e309cbb847496910f42b17bdb87c0582ae4c20eea5b43e3bd30914208054663fd9de0bbc270f9cac7c907a4a931dd3366ca7e6256a7e66571c5c0f67f5306ffeb29dd459076e1b2ff3d5be996ca48473020f413b36b6dd53d778258f59a3812d556a8a95cf3bc1631628cd53e31f32a908999e4b6aa4b87a71f282e7fbd4ef463d20960d9085b03e2ea69e088dce90151d190bb584dd314e7be7f7ac5082c25dcd457cb059995fcf72c0e98969d14367fd375;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h619f0c8676a066fe48d90bd5d242b64ee0a80ce48dfd18bb6e4ca8578e661d053cd7c36fb464a5ee8ea81336dc5fb0d9a9bc9a7c5bd37888c6cf0884fb2b41c3394e90cafe586273773215642fc69abef6897d26f8bfac6af44a90128eb2a731baf100407acad1161f6041126327374f22ca5a825db17863c882ec507cc287c5606ef4b3784760f4d5b5a5fd092a3910e575947dc961b6de9cd25c3267a6d6df8402b613b8642e129bc3b0b008925af6387988632596d947a6609d702b2da31273c85f0db19c54f986331487ecf8ba1ef63d2a1f8a0ae365f17123e3dcac67221eac391820bc7070d18dd905f6d8ad02a223a970d380bc4a841e6ca85e16ee8d26684c492bfdcd3d954706ca462a34eaa555f55dfa3a92b54190cad3bed54ef04c850d53b98803c8714773d7bcdc902218f188da03c9fc02d86e1e629b8f2d69041b90d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha2e9955bc67c7bd7586afa1083e1f1ca053fac2d965f5f51cbe9bb5162c565cdafbaa591e1c3214d8d6f0f5c5c52cbd84509d0ee155e4e9a61645e369a8992529df32857240a6eaaceef8bedde54fcb48eac7802afcde2fdcc02a31241d8c374dce493db371b0a05320ce7da6df63b802c71480d6f6228946969980c07775151526b5af0c918a3aff22db2a20bedee989860283c010e7711b00ae6b327ea7482a504ae89fd0625c1363109276f743061b7bbee8f5986d7c36dec2cbd8cd73721bba06a23ab07a5ad79b3955603f6a536a3d4b68a41654afdcb965d79ac69879d814372abff8ac93e10bad57518a4eaec5003d0bedeb69e303ca4a6b8f04e0912691341075560294c27c824236672e76f2789fe3dbc29aefdb7d83a39a9a17ae1d2c38407384af4de8c62355fb8ec54aa69af3e3c8d4db0efcc6cf7ce81e029d87febb0c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h78c7bcb02db02eb23af090e4c25c4207c61665c5dfcf42994dea499388404961897eb98a6f76e77c6cd187b38b4a5a9638d84d382f36024ad4c8e3b8fafd3ebec4f684db666854d2ec0c008333e35a3ea36c9a2a5b9f12bf1352ff9e4f24f6eb58d955e7c723772f06d8ae5142596e692dadb7b3080f67d8f208e919d4874f353d1bce755ac60630c081e2668c560238ee7a9e10de24313d0a800fb4b7376252c22b0fbe0f9920b89b857a551350799e93584dcbbc55549449c1ffb395c3fbc0c39fc22045dfad7fb7a4a3f5e20d4dfd38dd587022b018bfef3a1ed696be99e368407043e64ab639a433c34754846848d056078728c39ec27c5ba869536e7d24f5494af8d408e91b7aee3a5ae716e489746d2add615db597a6b61b7d03776521d25248900d8a9909bbf685cf6338e50f69b5b2d5c62a95002514119142479159e9904f54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8d58206991d9f7bd83350b25a2e42a5c1ec64744c7589462c1420ab250ec997776c6c3c02e7e0bb3f4914e35babce404f52801f5244ed8ac6c7a4b0f2588994fee9ae502f205901e73ae5a3a18ee92c653e6a59231c6c32af24509b91e5155f9bb072a6d72c040248668f1b324ad1bb36c751aa4f11af311df467ef9ec62256ae9e052987ce51f355bbbe83680e100eb718a4cda2c825b995302078875d1fbacdd897954659af83a93af3b1c114fe796e37e8a211e4065a794d83d4a0d842dfa91cc139d49034dc4009b7480777cc6357642f9e3b55dd5704dcccd6590d9c978655e4bb4eb5f9304c8eeb21417dc646db32fcc63e1101ba72794accf3c475fa483c0b4554479db06ad94f4fc502d79e62b6f0846a7bda0cc44c7c5acdf321093713706abe712014d202b23f354804e0051977c179d2ba39e6dcb769dbbe23c00171eee3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb8f03576a568e1ab1bdd1b83dd9e4f481e233b7e650b4911bac270102505bd285dedab037c19ccc455cc9f9173782db13acb91558b5c8f649c94d931a280982ecc553ae721dca122155c67a6f824054879aeb5fc775a9acc494807a1e9318a02eb8c7970166f2a5c2635e297f4aa0f84ecfa4967891f77d0ff3d24e98703cb90e8c4bd49f2920bd76c532d9ce8df64d105e70bad29597c9879f2ea1c68cf265ce88be567732b33768481f88d704e0bf7f088104bf1308020f4db44a788362e61c1781d524ddf7ed673e9817df2703eb5617d6177ad8bb2e8c5502f384c78e582e3f05f714702053b5ecbc8d727b10cb2d5fe30f9a15ab312e7d1a19c84da89cd537efcd9b84990c84865466270b1e33b00ff0e136e6ae9b91014c34fbaffd267ee52676630c0b59f74ff2ea0127d87cf9290857c74ae8279af5afb7c761d31a856f3f193;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h938bba90f21f263533783bebcea4689c0e5dd5f0b69a460244fc73653880d94bb7c3190df190817164bf986fd9ac03fa2c8e8a3a66d09e5bbfb18e175b1eb06f0c7413b53c2579259203610723e2ff2edf5dc77c2422d8a03a520d29d66db9d14cd57ea95a623071ac46059068df766ddbb89aa6bc8258a7ff8160edcb758199cb06ff3b4e9d85c0af3f91a2e1196df91387e196853873e506dac6464d0d9a0726f920776794137ee1928c6523239e189f6fb1ead6014eaf689c0cf90465f1daf349133a38cc20213adaf662c1a6688ea11edb1d88ca1a31aadd0f33f7f809104edc1f57fe32a11ba0de8d10c47fc94593e1688d3e7bba2b013b1738626412a696e1068df33f2e151ae512154bbe8dee0b8ebb9540a98e548d51919b5e3cc2b05ded2d77c0dce453ff0fcfd49cd52d9277ac0c4c1e6a4988d020f88caad6bac404a5aee9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4f5a7ad754fe7e89ffe4defeea79b21bca71bca88988ce91cb8ab4d97cea65e988b636d2db8b948f60f09a9bc45ec4210819df686a003550c801124edc7b2f110cfe27336f87c9e616caf1e474e7420368bf7a7c61fd6610e118c0e2fd796331c5bcb8461a96b36d777794c5613aaa528b3063db4a7deb07ab8da7ef78fcd96f330b2d7ed79c60aef3a0b993c367c0ca42cf03c881adec516cfef0159ac0b7691959669d25411eed44e1823cd8c1f3a16e14588948d7d7dd6a63e21e947bf996e92bc9806bdd89acde447db4a59af3c052a70a5d65d8182acf7db42e1610e517c455852297780dd8795d2da71c2ae4a1853173965ff874ebf58e6862cc3b215daeccbcad7e4e4b009943b58a9a6cb854b7c93dab6e3f1e84faad70882ff35fdbdd6eec95b8bbcde365c327a052020ce0aa7a1a2b40dfa7f62c62ebefdc475e6673866d82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc31d3f03e21b4a8936297853f7be0ee6c462e7805e5622b0bc7ccce148f25bee8ae3f1126939c8eab4bc3e8e902b2096ec6317c147e95a267ce24ac3089184ea2841a1d286196253de7033a5874767ce700d67efae3f0029e50c9557043f13ff8d0e5f2dc81c00f2e819e4278e8e7137f14addf4861d08a830df79ede998e691c5d314a3ee3b46e595d14543f91fc9f11a8bc1720e24542422311e161ae3b4f249d05b261ac03c2855a2052f1d9f26f61473d1a305d11e5f0ed2abb167daf7a2bef37aaa1f46a7ed26ba3a5dd00eedcec9940acc4d275370f7b91fb930909c2f32540908fc44b132f31c6b3d0faa0765ba72dcbfb110b22c7fbb3574895e7001e277c91458ba245db57943e6d4ba7da03fc6df106c9f3421e05f6856d0799d9338f37dde429b09b5113a1e039c91e3cc40ee4acf85033cc49e0e565704e2ab6a6af7b3d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd0e0b620a3d7a8a48989c7af3f610ab4c80b4d36c946a4f473d5def9f095dba84bfe475ab9077a2e295435e638e91e58f459ab850d23e058f114978dc55cebd7b5ce2608fd18b731d5a5a488209b2efc6fcba8702b0d7433500fea87817d9f2789387cf47bfbd8176c2682f2c4965620a4c35e0a1671ef6ca7413971a9ff3498dbfeebe91ce64ab16f64f163fa95dcd16bd3b6de3addcb68d3c3cc9d3778f6f97bee840e085f012b3669778b61fd37889edfc13c0383320f867ef436daaeed81252602d05f37f26df36a0347e1e44fbc0c39e4bb28dff984e90c817087834f1811f70e6244336c549cc1d9d4af993b6a5c7624c0de839ea19105185345d1b279a9fba49e51e219dc40e00835fbc3a636f592b54822591697c495ca9d754b8e2a3610fe0f79ec076e4c2cd7137a522b57106c1fd7cc9d8058111da4b3ea686a9c80aa1c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9f5b1189a5450499d1f09aa4019512ca6c703639ef3af1e0e74ddc8ed9773a2bea0998e4bfb2f55d2aaa1dd7fb72e6dc05a808144321af1e9c2be3ba476e05814f65b46fb72ba845e2a9ae86c72c66244625edcad4da4502f15a973c54e6b24838229580865275c5684c956b11dd4fcf492c9b5f084b81ac55551f4e1d12c4875eff14f94b5858b37b603d8824f99b3b6e2b09dc9de8013052cb98bdb21e5b80ea82091b9b63a9c29850a0fc31b9c42ec2d1083ff41a497be8d850e6726cdd4ee56d725446757d888e36c96d521925f13468fe4c90c6d32df75613acc6ef937f30730787348e08a1016c8d4b2d7b162b3c2509e13d05720e195962beaf495239c706d03999a7226364c11b572f81539707fd9eed922609fe1dcb2e2587bcee021c4d199ffa277cba8f6782786fbc5aa5e1e874ee6ff440d3e07a9279ed91ff711aba7b77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'habd773d7ee55a8a975b772013f64bebd4342dce73ddd9e943b4e2a941c4c30dfb5b4baa65ebe30658e1fbe29353f3014760ba6f112b5627d57fa8ea7df20674d4149a38086388dade9168af9f60c89e6b3e29a2a788e093e639e60116960902d9f16d253d0c51f9761e44769d374313dda31e4c1e93c70a2222c5398a6c22123e6e894a43c15e19ff09615a46d3df6820d2105c3a178f754da8134c7e34317431895d7c9d90cbd9fd8f049c0337570aab7c518f2565d9ba536401edd3318b9f61d90fdb0b7680f9bb2e85175f74e042892b5e338c9328822c18c2623510a09b7d8550d27b0a4cebcdd2d48ae53e9f82855c2fc06cb79068cf97022cc45e6408c79f1fd5bdd1bdb1c1366b3d92f8c58b3ca8c4c83ca0f21406c0623665c9181220037346651c80197eb96926d0ad38ef6bdfebde59b357de93ca710902d14093f3f675cf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hbdab50117dfdfd317b9c4a2a1e7d6838cb4e53e34a64c82a03c9577a8b1eefcab3ca847ac68f2c3fee632d51cae157aa9c4880ce86f751f58a90f6e739fe241a899c26530b5921fdab505dc9fb86d5237414d798d87153b1149e1d4d24daf8e9365ce4e9433730c16b9a1a3cc929f18ce3c3119b332180af2cc191f95c2bdee7a8a2c3a7079633b7113d5d9b334545cb1ef32ebed514ec2591960058ae56dba9b1dad96281eb0a4558eca451155cdf4fe56d1f0d18db0b62f091723bf63e17efafcd8fe3deb84d9d32233be160db352c4e36df27e44ddeb58f1d4d91ea15ae90b8dc684c790860b3433d63f20da4f782e1166e5cd834a9b65be423eeec5acdf07316ce4a964b5d20b7b32a4c23c8de262da8246d91688c1bf13a6fafce9bba7470c8f7c2b8e8706afd267188aee4cc8883edf1f16217a743215e273e5c60b1fb0f571cb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdd5f48b183f706f8a8b1eef48a1ad044f3e4c25fb3c990c3c1b593fe267aad985d2c5cb8c5145c651401cb1a83fada0feb5b36731f270e11ba1ed0d57da9fffee5f3232a6f5fb7a46036cc92867a74f8234f0ffb84524069b0c33431a49894ce8418a81283708cca28dbd6a262326cd29a07500caa861ff8d579a337e5b62522cc8e986f9707dc913d46d9879d5f6053b2f3410b4ec2b020bca7a3e33c3c613a8b3c5621005cd2791e9cdd9fbca7a8d1fcdb1345e99f35d525a2ebe1b48f01337cd629a89805722c8f281055fee4a07057fe5a8638a85780a6c8d03f90a57e80c5dbc3c095a1f0a96d4b19f8fc704a2c23670517ac03fcb2f48cd84f546e8e9f68a65f2c52d7b34e04d8b547caa87f8429fff3e06d7bfd0da7d507458aacf85eed9c7849820fa88e7920c63cfa815965350e89b7892d0c552692b1fdb9199aea60e22bf7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hace7bcb9bdca56b13ed56b6fa9c03568baead7bd512bfa9fc56317f75d35c0203598e9cf4e3d94ced836f149d354a7b5bce33ed1a460c4fbb3f95f3fa4d61dc9f0ecbd46338f6d647a813ecad76cb74bb4efb01f1182a8c50787ff073f03b6864f6cb5d86f122078fd2d559b11207ff6fc3edeae62ede2da6ccc163eed2cf892136ef77d63328340f0ad1ed67a078ab6d4bec02027b38a02e888842066e4b5fede9a546ea20fc910e59ed4f68306154b72c7526a17d246342f73317020ce73088cf907c7895e2f92f8ef35cd616a50c07965833223f17a13dfc5f8a5f40567fae09a819fdf9d84793dbf74d0847c858ea645426133f986cafa4909412c5cd994f5160c473c1ac6b501fbad56a5257602179834e60fdffe1d64096df41b99436e0b67f454859567f63a3657fd55dd7eaeee76fa74ae916943818e760c000138d86b3d06b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1a85fd06d68355bcc40ff4b0d44e52b7883389c48d8bf44b893b18311a28ca5f761700dd09d8821bf3397b45b65b9020af6a883c01d1e85d3dd2ef4fe5e35bfbd33c8c24011cf85ebc9019d0cecb30b948bda1e6700bca8d75e476391a8170040b9ea2a1e8739a8e55bd958c1098df1643297f208af40170386e2f7d7aeec3e93d51dbe7c9a9aa34cb962c9c23b7bf5395ce6fce1ac6eb08894ea0917d16ab51e2443eeedfadbd7b7e5dc25e157e977a0a41f51593af5f789c27de7e715263361921e5440d771aefceeaf294fe4f4849aea58f32b35d6f1f9a5986df1f7a7f90d951d1fd2b697fe632e8c4533bc887371cf2054b72cb55d146ffcff8c6f04338209fb1719656d32184dfe649e2b7b1bd782e7cff1a87dd388df48107d78e6a50b3994087ff667eee2daa07c9e9fcf46779d270d41700724aa24784fc9e6be516b1089966;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h43b63b6bb39568b94df9feb5562fe95eb2bd02e4265d9bf24f97bebbd06bb591bf4176445ea4ebdb13eafc06d1c2378306691503f64bd02e3251a95d2e3115add1c4ce30deb363e21ac27e074671f35f1596c83e5df99f4f59bef24c0e996b9b9450d1096787e600a080820397a0aa24b827746f0b8ad87f5664bc2cf9b3b969b1b2b56d5526a6457dc9528847c811d4c227b910a58992bcccafc9d528bf93ec523888f57674c35a4be0f50d28b2f61e2bf6808fa7caa4c3f938fc1b173f31d7913358b919ea7d9a00528efbf49567de7050ccba216c39eac911296be302eab9d6c9a89cf59dac651f1cd21572b94244500c825bd9c38cf981dfb8bb6f0f5f41eca00ce6fd1f5ed1c15228805c59bd8c6fc80783b969f022b5670bb79ddcde9cfdaeff4c0d18e5ddf2b1cd1030248ba4a01bb310731027b56c0cf43940b12e0baff09852;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h646c3d801c66e240c62ed89bfa397745d881fb6517595aa4ad78809ab7dc5b563346e9c204c4c48595ddc791ab7d045267ae85e333a549ffe73bb7cf9d0a1da4a953b2ac2758da8af42ca7965bb2a9a7ee2637cf9edb11da7e23807f7b14c35dce05d1eac5cd30dd555c8e8f49ef132d3aa42a32c8f5d55af4186d2ba559ee197336195592b970362d92cb5269fc981a5a9c8f854fe9ff3b9a4832d295e14e5e3a21486728017e96504e7166ef771d9e18897789ee871c8312cff0ba6c942217f9a716c38a51a35381e3fc98ccf73abfb688f5edea5b88804d030ac7dc3e17e3561a6711b6c43fc0ca7eb9537350ca6e42a063d760772c361bd0fcb34d7b99c653389a9707fa30650c37f414c3b8d88118df556cf7c3a92f0d34d304941426a9a2dc64fceaafa40cbc4cbabff8fd06d50b9bf82c742dfcc6e47892c0095f7d9e1ebae685;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h7c2e6c1754143252f79437013eb814ba82fdcf64e12ddc9d0b413969724e7c846f95d589dd50b873181a8312d58fe57a9f2bf6b7b914689b873f9a9053d0cd6e26bdea46f51b46a3f08888ce5801478969efd3790d38d73d3fd66557dd3818d6419f93de1f93e57e8cdb721d4b826887d14fc363bb0ef5737d7ad23ecf4e5aff86367c6d03ba0ee7c12e424bdcc24b9c3a55115710cbb48f55e4c0d906598313b5dde2f9ca62acafbc20219c45f2d7c34d9a287eedc694af36c2ac4deb7c5c509b54db36d027a0424f8565e70bba135afb8ce8a7d515ff2d6e1591f881276f23a774ca69f061b527a189c17f68880731d483bbb8d867e97c6571f55790141cf8bd4097cd4f46c1d794353dd33b40fe1bdd8b7e102c734bfde2020f4577e1479e3cf28c277b63915adbd95086720f666cf0710212bd89491d01f00f767191eb239afd1822;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9d52f895762acc181a4a7eeb3e41dae44dad44e06db1634c2ef82d8e71c1cd3ecfbeeacaa1fbdb491d28b6e947daa56da2ec80eea26e8bc865ac976d261126defbbe826159f819628b0bfa46860ac802819843c98ab9f4c9477884084a4178c1f8036112dd1449b9ffc7a60a245cb0dfe7d5b647a7103c715f9d76f60a0be912fb705096370f3396c4e6aec317a5485e49379533a373a51519eeee171d5bda8611a3881dd5f4422cf07244c55ff63e3f3de361ae45366b3e8a14dc3070af3757731db5f79b89d5e63e5f967b156e04df0542da9506f002f833633cb192863819b5642d2aea5968eff05321c6bf5ae9852a817e1dc6c84ce4ffdba87b8d829c66451de11381ae3b8df73d70e4691ed9f4ee2cc62b4971bf26e32a65cc99a43970202b436cf023b0a088793f711dae1393d6b9250af4162f26238c023f08c51a1a1856b4a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd358bec03d06034b4c65c792ba23b52e8a9030f3743000c8c21fb05a8a05115a9b921b2aa54d1e0182ccb9b99edd0623b79e302707ba1ae08d472930abb37c52586b586b4a5bcb5292f81b14f903946f86567a071f9d95f70b16af81ca3353277b5bb75bb2e9ccdb878622fab64929e7032f01e0e41d862c493b0211ad8ee98c63aa5e9555f7bc002c307e81417ae2c9854933bc7584328a87df4fe1ff03a425e4efd83c0dcf906adc485c6488e086c403ced5f096e9a48887e3e7ac519bf1e4b7dc2de2948d442251a6a29d661777a4d51055e11a77492530576d24116e60ddf9c51018ad074376bf349cfd352c666a2f8bdd2e5ffa33ee6ddf24090b4fbeac68ec6a7f5fe519ebf45829c713a40ee2246952fde72f7b458fb13e29631ed7edf74e1f175ab41796e8cf5b33e4ddec81d8d6859956bbef240dc211f91172e22730718221;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h90523dfef7e6e51f1e41009513d37da8778ef4976cbae46c6daa0f188e421be8f51ce50ba3c034458d91511c9f9f15690f56ab94cc791ec9bacf358a7344501e86552c06ff7b02d2b9f57d524d3f2bbfa6a80b04c600e30e07f5f0bc980ced12a66926378232462b1bdadd2e46cb95d57b658c162ac755462ed109fcdc45af132dba4bcbfe2ad0d692c5bee5ba653c0ece7666533b8073800df0bc6185d2e224f4254d0d6b6280ebd39c27c0a2ef94ac11791cb048a3a3a0940995d730d8df59b7865c9c5bd6e61851aba7b6099a9f1f63bac7fe90b03272ee719cac17d7e72bdc8dfdf1dfc89e3de7b610f422355c4956199606f58c8acf803a9c23ae82d90cd6bf75f5bc7fe27a608b3fb89d48bd1e4a188294630fa931a19b137ece3d99abf1d6603b9a1c2811294ef7a3f7508303b35f1efcb1fd5e6626ece3a81675f05bdfb32d8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf42bab1d615852b1fcf53345765fa004614b8c4357d04ce47977d7f23172c4fd56646c8f9431031deeda0978a654645ccbebe0015b2f6c9ddce1aeda3fb1bbe77dc50319637d0b1a73291207bfd61b6fc1f885e11de94add6570d4b3da03fab94e4e9ed9f8cd50308e296a0cd367721210d643363d2b3a372ba9674ec907000e30690c515ac2cc190cacff9af7cb3ba16553e1ac8465c48497e80bee6772473406e69b238d0f567dc8bba28ea0c434b88d08522372562d5661d35461878ae9f84c94fb8f624a86a1a2c3bfe6653679a57cf34833d6d97e722a25b3de2ef71b6efc8201c3f851c410bd914273dc54f8a421666378a10847c3779119e02e37ed0e3cf0c6b3ce93fb4479e7819fa356a1885bed9f380da35be578a080665739dc53f1025c37a5d49727e2a275ee5f69cef6ccaf71252465fd1cd7d56fc0b1704f3252ccde53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd43bf8f90e19057b4b7584f5a07e3bc825e27eb4d3d281f6c63f5cdf827e6c36ead378ae5160c62d8ef2ef840947a2eb1126edd340e99f604c46067f04a833c37afa0f069a4834029484d3221d64657d6eb904c7ba9128374cb554e2dd5d83246441f914181fea617251536e129e4d67b7a6d63dd50cdbc0eb0138f47d7bf2b2aa7edf041a42f099f402d67bc4ffc415cd37e029e242e6ffeaf8b1e0ee7a9e76d5820e294ba495a01ba0d77e9f381e753084325b11f97fff31816530a5fc6d34e61a022fbc13889fa6d322d832bac0d2c31112bcdffc526a3135310a411b86931092e7ffd50cf0e5b9393730ece60d6dc16a282b0b24f3162c9e8c6a52868536036dd6dfff34f13dc2c6075e7cf7d27bc586d820cd2bff5ab92557865dc7c9c06797c5d3dfcc11de5c1a31c51a5946d7b7635f84949830613b83db66742e96fffbae5331;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3ccc36a023070b50d5ff57096e497790b4461928d2a62a37ed06e6cef1fa7b29e37c9843e8e87a946c30109d7755b203fcfe567b31a98126a4aba9d98169ef397e35b6bc91f704f304b336ac2c1c5a75fcb1528df892f340dec88058336f70fe81aa1ca64568b54ebf0c4af85f4aa180266015e10f00cd3919a361f5056aa5e7372fb80f376f439f9cab0a4da9571921f77cc9baa2f6d9b848eb004e25414fb284c426e258944ff8ad712661513a4b8c5bd582a25c0b5eb3d131843a49776efd40a101c76ced2282df8516f9c58a2f978f750eb56f25b7b2aef94feed22b0d880aa036cb925c0d6dcfc8947f6afe6deeff6b2a4c8b234431ee61bb5a36dcad2717931ac6b52e86d689f1c95ac4a034727aabf4bc6549a0a71beffc2bd284f96b2ced05da503d1fbdc6fdef8461be5681366b66a92200970cad4985531f14235e7ba8658;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8a0e62ff09cef2ea16781586c1c15a1e208c85b6a56d98e9b30d98593170f59b3cbd734eac1d90b67891189217e3b7d8d741c74e6c539b3a09758707ef48da2f01fa1876f4ee7f79320b1755626ca4f5a4489b3f9a25039e0372e2856c5e3bb7a2725028a661c6841ac3b9c705223a740a25572bf0acb9f130debc6927dccb949cac3795d91a5316a15f50f9289733782692e3263087918a21a9308be8875ed05e65ec297b004b08f169f79d672aa70b2e6da825f07abc62df79fe24b5ac59a789b7abd276a20acf936773b1c1b1c5c5bcba899e39d66fc27f90479cb2600824db1c7c32d77cee3332bf1574e79e682efa006fb80ab7144fd89d6f72500559adc17afa901c182c7e1a887a31df85f4ebf19f2bc641204eb9d3261bfc61552ab73c53c7b039f41b75769b6ef56f2a52b9d9a67fbd9c9befdfd4a7bcd0ecf3b4b6e77a39c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd4601524762cb0b49eed21d78946b6a60b0088e69badeff7a6661881f3fc7148ce4a97d21bf73a8331064fe2b6aef135d856a0c63a7c2aabd294899a6ec818f100ff7597bb47cfe4ee1f0fdacfd75b32cea93ac84ba0b5c9abbc9fde6edba826400ea942a96984415a2e7b626bb19dd431fe4391338514c181c073c7c12d8c38ffc16cf69d3deb6bcab291f2f7c5f7442724f24206c6f35f5a971c173927977166630b65f877107b30872127420cea746ddfd7c3dd15e6871b385b8d6be9d2e08d9e711fbb27a3eb905707a5739448c1f51f3353061b097ec9e081c667f3c47fba627dcab23830301481819d8a126fb457f7b2e91146a472afd640e5c840c2c1e0148744fe7c1df17099848d9cba550d14d8c789205a9da88a622861ed3d055f2d20454af87896a240ae331bcdb7a441336fc514c90ee1daa3226eb0ce753161a35d4ac1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2b57d8fa585c2a4bd971c23317f7351e5e97ab70a9705fd365c9715ff893ecd276555c638e65f1e17e57b1c719ffed30153a4849f10cc0d8736db76ae7ed8f23813926cc7acb80215bc274e670a520c03e2295ec5fcdd251266e7432773d8f4382e3b724829e018590e98fc8494f621b17f5ef0b4992e32a7ac10573fa5b1943b7d0b8a67a1b1af626341ef27a09c5e3a2d1a1d3c2b7498234060dccadf97ce4ef2cafdfd54731380b402a8c59d1858beffb1de83aa19f546259a4ab5953a44d1646a2f5df8e44e960f876876f4db30c256ff61483ebaf04b3f4f0e0871aa2f94d6e2d65e3056d864d1bc5f941c20a39a68470a343fffac02fefbf011dfae39f5d85637e252f4e787904fa52a81b00dd68bb9aa35053e7d987cc39f7be98f87e9dd314884ff569bbcf485d807e92f8c6f543000241800d03d620a35acfd1bcee277060f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h634bf579d9495a88c8f0250f62bdad7a764483936798cc48a21e61757d534c9a9abdaefb12302bd34a63f9fa9a14b6bebab315bd70e750cbb84a218d3ed6d2734d910a4cb94b2cc06a2eb865aacaa912222016f403ce3636f0b14c7a16635c098a45be2efabd6d2ca277f3c177325ee6971d5ecb51678a0a0ea619891dadd71e35bdda6697bc219f231c9a7a76937d94cba5a3a3e65d171e520ce1bd2a082cf47b5a52d4c15b6611f4b0308d900362867cebb3e425fac4f3f27822e27384d4dcb686d99d77440544326065eab04c8897e04d59e4ef3fc1963a7bac1ac0a9bcedbaa957005deaa18ae54f6326bde1c18a3b55f30aad7b9670db5e8cd4e72e071d3cc705ef15fdddc232b93b9f432481ec16cc5e0d8af7a59faf94a89e0d8bf9385a7369f3aba16e22c5dc95a8e5d7285977d258ab97bc1e3c558a1f791324951a581bbcc0;
        #1
        $finish();
    end
endmodule
