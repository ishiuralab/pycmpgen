module testbench();
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [26:0] srcsum;
    wire [26:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3f70db79c658bf39530d052ee760984539538ef17e5f4fd51d924aea1aaa884d0066c16aa1eaf72b75684e5f4c18709f5b17dd5750d61a2efd40f797;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae142f5a7e6de67b2bb8baefa631843d46466ac5dffaed63ce5bc05d044682cc52a5b8840498ba3aac1be259b5a550258fdc6ad17599062ea0a8392d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcac7310b3c104dfbeab38fd1241f1696c4671b92d9ccadb2008cab4973493dabd9d334c3c5fb43f9ce063ca8aaca7096752c1f0e7ca15b25e630c7953;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95f994f4534b0545ed9e6ab643835c7b7f2e32eec816db7604ed43d9b53caf88a8d37fae60c1fd3408c7175c329cf27ac441cd646f8c6bae15b5437a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e63c2ee6518d06d9239b34567c6aba216fb7490a20c130955cf535c61a31ee47f534206c33206354bd425903af208b8efd3e6e625ec00e9d1c09e8dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18cf7045ae74aa5ba0b1b6a60c087e6194a4053e86db195300fde6b888cb2b820ab297a79b49af0634723966789744ece0fd333e0bdd7a5b64167d25b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d30f967833a2dc23f7464db9416d5e857382924ef7a3f31ddffdcbc35360ea4637acebf054c0d99ca04ba84397e2112bd168ec637f3ff905b5bcef2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h433588cff376b54fdaeee5f5230c302e1ed600c039167b66c98d8275981c88c5610b1b13ef356d13a30bdc02f029e914d71e45aba60b30d738cea3b27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h621a76232baeb60bf71dd8eab2754d791a9ec85a17911d09e77bde17af18b94c7edcbac5f1cb55f3f4177283eb4b8edead7f332b8523a82881bcec2d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cf2480b47f5421b29c90d59ca765ccd34aebb226f5759e71508157c7e353fe30ca7618cd41189e7c34d631337c29c9530459e1cd15bb5eada1a77c2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b29f1d253c2d953f4654d337b50b49866d1b9825469ecb56e365f611407d62bbad299ea79c7cd3d09aa315790aca0613a5bb48084a96fae7f79984e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c4f12023d70fc2c03148ebfc62f4391a361d1facfa2e7445e0078a9a30310ddbe16541c14f8e59ad59497938007da7673c133cac3a98f776c8d60c9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb97d8ab2a060a615a860eeaa307821e006a13bbb13c4c33f73c44e058eb200ca8636598b03f58a22c037db4fc79a524d9dc1b0d1482b80c9150f47f13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1013cee8b43ab12b1469b440cab56c2077b76b91e5c7bbe1a8a67dbf56482b96deadc68fa20dc4fe8b873001b074c7fdd725fd308a0935ffc2c1c0e43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h715d65438661cf50c603a26f6b4693ec5078f05b30cdda84e991ef1a7067adb2878d16997384d04382ef982f2b34f20f5aee054f280e7e43d71835cf0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h446825092de25c9a0738d4fd6049728dfba6f42203c21e55ae70d2feb977d5a5b17b00a6eef704ed6a0f2de04b8fa6cda8dfb675ae5e515073db8f736;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eab817da3cd9c49dfed6907d2e12348337f7e6f5f2e77300a647e4ecf49368ad0134e545d38d16c423db548c054d50da7ed4433df3f4a07ec27dad36;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6176f7661f370a1d3b087e5309e871754628fbc4fc5354bb4df5fc8fe5279f241c7e92fc50dff3a4bf44d3ac5c122bdb3052772a1942cfc80094b65b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h453401bc5f600a1789100564fd60608e118cf1a3e95d1a9d2054bb2ef2955e284031f35e6ebaf019f8f5129a14fe1b40f02a4e77e4e4518b79b34889b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2eb3335a7507188816725bc817c4f3feb4ee6be24a4c69c6adb59de1088303115482245f269e9a6dfcea75668e6746381b9f6fc8acdff773bb0a25b79;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h184908bd55f52066f4a3d2c6ea815c66b98f52fdd1a211d5aa3363f240fc12bd8b748efeba8189e119f8b3074fb7d312792ac6bf923214be87bd82b8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdff445606d9edfed77eb74828301954de8cd4345fbc0f01b78d64854708392f5336317d3a46ef7f59f9e295060c8ceb598703b34b3d2d36c8b8355a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64485e9133a92804d60ac598e9b0726e499362ed72c06e07e7eb51a382eb980dafe09593e5cdb1afe2f4fc32621fdeab0f1978085839afe5993d5d7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habf780374a40bd91b9e2ccf032e15d134bc922e270bcb914406bc93a7bbb72485551131dd78e5516572f151d8517812f0f2c9291328c13965a6bdf037;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f6f88b9a60492711c17c2f0fa5b425a2ea95bac2f3b4c6130ebababcc14688df237ad004b365057581e811603050f2a5362f0f49225f56fc1174d958;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedc9da041306643c2dc053370004bf594d1720f933c345febb1c14befc8e78b31f962915441db5988be9dcd542bdf7ba26308b6b027eb76690759ca8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff748416bc3b276ce5f477d5bad9888afa482e874c7dbb0cecb97e12abb538aec3fb70a8385e897dba3070bd0c1bbee2cdfb544a8959d272ede615bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cc7120038196be96c53bbd66c8680575fe905fe85440cb372ac2c881f641a679d78e491d55ed930174cd2a89dd8f2cb8783fb5629258898b46b82720;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68cc6a46b2d0fe6195e42f6e1496e9fe7312e15a9fc8c236c9298ed16cf0ee672a73093e1cd4463b63df6e6f5489ed774337df25948283f8a138d56d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h619639626fd8e36d5fa98a0ace259986a91adab1385ce33812a009abd0c814c6ff19e11a1d2cb8b55349968a857d27a2ad9cee82ba4f6d00396d84bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d8a991b926105cfc2e99c7032ea73e1ec73ae677753a88db4269f0f2ee7051bbc60b80908abcad259c7e84363e1de9313f9346a5761b5eff342ee1e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e404616113eff4277ef9a686d325f862b9493a948efc7432f64cb43684aab32e98b84033f0867de8c5c30805942f60e2d061d48c6cad187cc2e06aaa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85dec5c54afa11a968a04102c50cc680936db794eee2dae9088a6d9290d186d23d508014b86fb6670d4319c696e9664a45e112ce0f0c3e13a541e14f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2053ec5dd96d438f343da30cfc0e46e2b95bab3647efb4fd320570a688f72bdcdee497fc7f499a0cbbd1de603ad0aec7e41583342bd6a0310017b9c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha00a94603de2a7e798abe2970c81a5446e07b233b0db0d512b799d63923a09060607e3069f37c7db33eba8716c4b18a4f3a4c1c5be9b7c22e4b3b6b5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2f9677665dea906bd2ba85f4b2fe17a2f7d49607d5713af50181bb1bf9ed994451673b8ecbdffef592206492cabed22202825801264296a312fc6043;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a469e68dc3754bc722891dfdb2d954150c95da9147ee6f87bf75a4ade55e52a2e268f94455cb65dcd17d79a914bccf29b562438d585b674a5d1e017d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h201105313f4693ffe40667f82ac844b817296f3b8594a997f5587ee9ee2ecd90f78ebcb6a32af327c0c6b91f923751254e4e6d11e3d323af6be032e57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80e596455991ce8e005974678e4b279ca80782142e0a6a95ec34591814331314e5e4291150ef69276027e761ddb50ca700b202c127c35bbdc5ccc247;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ccdb36fdc9c738e5c182521ed025bf2ed76154d0c990bd762fa6b3c648dad7e0a63f73a0313d47c1ecc27e91527c91e870caeb7e9d72a6a56b83377b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86022a9455358e66fa9835be7d1b0eb46b03ce7c85d39e01ad4ba7dc20d895147e90575f812d3275d5c734a90b134a51815937d6d43d27378698caf5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77241f2543f38eb9e658f0413e4234073db3b023a6c8220d8d1e35b79becab7a01f2a042c8b26b235d2481bc3cdd0a844aed256cab68c830484163ac3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2746219b4ca8229b9ef5742bb7461b6d6cee10ddafec87dc430f006ade513216bffa3e62ac2c4e24ced25f637ac7ba0dfac7acfbd332b66dcba58e912;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37cf7b5ee6079cb197d22e3fa1e9cdff11b9264d0a9ae8864afc5f6c207f9cebc291e02fb210b83f8733e17ac52d6081f24b0318b612b02b299bf6d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44b43b72c000c8d44290a03a0f3069fb35fbfb04e886e5912e0e9e02eb90f26ba815630961aeaf209937fafd2f991e4a2bfd86811a3b36e934e4a88cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91296b8661ef1aed7d2d4007f583026c689a5ed5d3da2f1360adcdfc0b7beddec2a9f48fce19b40cc412f5d1848dfec67e5642fbe6f22e52324de4aba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb131c018a747dfa3e8ea96202ac76d9355ab25d8b0b09a3d5e6975275959e71d05e5189a91847c61493cadb99743d5b634183053c65fe071ef1e01fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2abd84e43650d7b98b191267748883324dda992190480cf2ab40c7d3c9e4b83f708b51ec6d8d9c561cff11dbc1aa675561661e23e4de913af42088a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc929e7075a7e67fff294256a9aaba13ebbbe48a5dc306de76f9d4bc04b9d57714a057461f117d07695e0e96f8eee820fa5a6e9c2e53acbe9f25374;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b7deaa7adc291cfc6486def228a05c5a753d7c7ee24e74f4fb6ab79410123f7fb8238aa3ce8d5ad072a7b3131f53f31a67f3fc8bb3a70a6922ed2e74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bc249f7ac9ba217bbb9eb2d6e4f4fc826515cdd66f77181681e524c142bfc5995204d95eb3f6bab2860535a4e58a9cbef91c01252fb5fec2f525d555;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d95575c297a0a6195cf4f5bc81340c42eb2a0409b5b15ecdee1ebdb3e86a98a7f81d15c9fccaa40cea2904cb86fa19ae1bbcb0c49b06601fd4bb5601;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5e05de6ef69dd19102404908ea0fcb92ffcd9a7d254b564909a1562f615c040890f38c1486af3e1a65d7ff2b2391b4a3d54e4f77df142584d709ae87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1930fe1cb5e6463a418b8a328d4ab946c2d295899bacba365d4dfcf4f5ad6eb6c127d45748dd351ea5b866be072f7882e7893b7005ade55900391761;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18ea2744731a06fcb1a7385491a5efcda51afaa6e4f635e3f3ea21d72106b37ad396b36f95ad0b682eb76734230ffb993814872c3ef51501f88b34b45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70af83ca731c2c75e061bbb1c4309dc4ab4061e1636fa2ee6ffd7dee03c5d76726dfedc5e538cf19859efdecec861363e4f3fe0c1320fbee171297a27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f6f621cbdd4c3f0191645fda87aacc29ae2f4a1fb097e3cb8754251cf2bfd00380ea88c36724d38e399a4f9612cd48502964ef54a12c183c965cb10a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1346fbc32cd9e93478387d467fe4585f1cd5f0480819ac74a6bba5eb894c29feb9858df162d41a52c8df4317f5d45de873aabb7a13e54863a1c0ccd87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h598debdcccd2a82f378ab19f67c9f024f1e3c71fe23118db5c9c73e1202514ddbe3fa1ef13a2ce3b789d08287dd7b0f591bf7d42310393f1fed831608;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61d2e330a8e72e9cd37fc38adb983c664c6c18f81f89f5ff8c2f361da905708c1650f7381a4b460162ae4079bcfa377bcb91357f3545eeb267c02798;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h149d083d32f127b47e34e11cb50818c2baa2a825919e52fca606883b729976dfce79f14b3b543a04766c0cbc46b69788d0922e94e954b7139315fedfb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf865789e791108cbb716f463fd0cdffc3b9a2aaa1e7848113673d43524e711d1b74c1949ef82b8da0882004bf6978ae5a6ee6d8dc0bee92ee3c7cde40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36f9ee75fef113f86ca113a4819afd97e853af72506d68bdaf61245bd6dc83f9421401220a25e676d1eb54093fda1930a216f19b191a3e40003f5ac7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3df2b2273df7f0bf3c8afd96cbd4af211d5da5805b732d1c79652f9846a20e42d84d936dcdebcab0577f44787e7acd6533b01b62b692dd601a3e36da1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4601e9bb285b0efcc41f218aaeb760ddca2ab48a738bbd70e73085f2cf6717df36fe5de09399b3ea51e248186db5064cf5cc234be2d664ec91828c1a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2508abbe52f93a6584dc824efd06e38258b7a400b2c51c9ef71aaba9890087c349da19be22794de6ab77983c1dd74f4e28a23a4e74df7bac26e4633;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79f5a81f270eb4ebc615aff87a0c82456ae71fbee4206c8c435fcf74e7cd3b027c73da733649cad0337f7beb83779f9c9c04be5b725b032f15f2c2ed6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b352d4b4ef29c5e7f572dca626c1cd7d22fbe838a1dbc63c723d394ca263ce604b4cfd0b9325fb4a01c67e312fc3fbdb8f83d25d031090de09a3c5bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a8303a83aa824e935122dd2e6f16737c1d61871d8a78c93ad93ad0b21dbfa5722c6f42ae6b00e2d760591331702d6a63036a91135554726d2e95b70d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd60ed47c6f7e00ef77f3dd4ff5077e496580c0670402643aa0030cbe5f783e2c4183d87595b6b11b36c33215325d1bda6a8fe97960aae2a2d617a4696;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb81446c0116a771e34837dcad0ae36354bb4c01cacd7013aa2301ddc85a5460bd23725707192267374e9322ed1a0182e41856981a204128b803cceee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he98df9301fc4c79f66b8cafb5275995530ad6d8cfbc4d5b3d1c86b9797756428464be3e34f8b8b7e301735c98051d9b2bbe4f8dbeb6bb5569e6e6ade8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h673e83b3055ef671161c15ec0668b622585fef35cb438e8356d1d5c4c279b27fb008dea0699e839fee1cb0bdef6671774285147c5ad464b0e9b97ab77;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75ac1de42034ff3eed333ca2f00f558fff8f32bac0f69ec8160a559ddf4db841b5b1739b84d70aadd2ce9cfc301554e30f09507a515e053fa2f99c331;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbee88f7eb9a52f27df3770f23b47e69f1cd1dbedf8b06d4bd8405ac8e8956bc27625ab75c2dabfd85218d2d7db41f1e8e959def87906d221c980af9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfea43546933870f68d29518f33b729870ce6533033c0cc19bf176e8b3f62596880528434375a983228e085116759ed1c78ff8663b438cf3e13157b329;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4b76a70a309d6da2f172be067ccd6017703105728135347458f04ca1db56f7db7283fdc4b9d6e44a742032d9df39ec7151ee05689128a6b7136a8600;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ef9f538cf108db1594d43b2a51c5e4e3f0039450d51d3b2c1304a74ddee28cc4d7664178565e062324806fde063c907dcc8273070b03d26e8d0b8045;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e336c30039f830c33bf76aeed8b56b6a17e1e08492a4362495844f2451aff0419576f0f61e51c069d27d771ff37de3dc2d257e45adad390c85f8a01e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1900517b6e6da79bb7daee637857569c69ca368324045e3e3d2ccc3182d7f2ff6954e8c61a61e928086d7d71f057436d284de31cc5fb4871f8ae5df10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5eb53c2a73c2667f7eca5d2ebc5dc63eaa9d2b00f03c0b22adfc03f7dcb21e4eb63715fe6d4b8ced0fb83eae46d5a46cdcfd23d2517f1793f70478311;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd3fedc6422a5444df51fca57b7e967e80b61207fd8b73738835ddd97b51d1808cd02905f3467267ebca302a8eed5a7a3edfd0fccc21856739d1f6e9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85d903bf427d447884b1f0ba70671fb673236dacb324c2add9ce35704f3408cc3ba2fa834e7cf14f9f680ebf54bdf733fed6a373435d79fa878c29bbd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56f12008e978447861e3034c339b2cc7dbc174c1916fb03d10288165a27eaa32cb9bdb4439469f9a8cec4ab765c245d0f50ad4febe4514594f2eca1fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde81e1f1dee08e460b101af6f4e4ccd6d52861e87c1374e193cad9bd1febf7a76ddad4f8ffcf2dd5aad2ccf63e3ce8b94677dde1add1e484222f428d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bc05d6a09cdc26e6a540b62d39b62ea58687066482ff95ec5608a5ff0327fa319dd9851ce5b36b7ef6589ff524b08a1ad15950a0e0a6b3a358e76e4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff1857a83d36fd85f9dc6cdfc041ae13fa5be56207953467712d8d6b03399be3675a5fc83c18fdbc62c58780f056f04e5b79a88f63e738cff5014127b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h401a4c6c84277752c0e60d957d5bcb979316c48b945b5fc4612649948adfbb9bc869cdfd0c52992c4e9b3706824556ef5524146423affbc748bef7149;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43f5348ded9b07ee40f1b29184373bd183196fa459aa69606ad8128e0189588f61541dab73170816ba122d855b481569330d28d99a06f24703e5366e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e6eaffebe0d15eec854910124bdce539f1dcb65bd5a256c227250d16430228917e1eb89fd661f1cf67e3d1104e53a64d71d6043a751e6335967b040b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcedbc81cfcbbc6bd4679af75f8457dd26835cef787c9baf8e8412d1a15b1dc5cd0331a2ecec305a26d495f8d996d478102239455cd93b622e0b64c415;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5a795e5b01d4d44856ebed8fb6a5cfe6aad60bfbcbc39903d8ef9d7c2a0788299b627cc621840813801daa3c61bca2be4a7ee74c8375d51f2386c98f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd48b1ebb4fa69764881e82fb842e9eba9c8a42fba41b0d62f3154a3880fff38b72776dbf494b6f56bab1fdfa05628c46ab1c140110fdba35fe4f2797e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9380341e18b423c40ebbcdced74a4e3131652a39d36a5b00b9a87929330a71827212f0e2f39227c2d0ebd52c2cf353ccb4850f34e8fcbf73e55f5a22c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bea1f8945923279741275a9b6f1c98453f3bf8f733223b56efc25f4f352c5428c29ffb6855ebf230dbcbe0294e8e6291e98b1316de9b826cd109f987;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f5fb6b5904d0c012a9808fb3f9425852b9dd30dc9f55a09a30cdeac7442ccd15f3b4c6a3c02551deb721db1ce65f9b8503436d6389eada90d34c1cc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c403483dd4b4491857150e8b112be52551bf2742e44d67ec91afe17b922e2c27a7c51d3f12ad35939b41be8486df24e49ae8753f066fc1b3cbd6eb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32e09ff9485601eea7c4e195a9964583fb68e95846dd71a797143e965fe7608d4848d73c4095e622baa8e771168af16840f251cff7491d0c9850e3733;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h393bf1f2d15d9d14835be460f6f34cdcbb343c929c2038e13d2a9bc436a4a34a17628f0aeb627c10faf7537fa99e620a09bfaf75f5789f215bfce15c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6aa51e79fc8d523ddac96f83746f0d4ed55daf969238bb7d61e7f8bcce8368679660ca5646229cefd9acaff8c31986447947abb2e09934ca193f782b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4cfbb3d429f5d8090786d62d981a124f426667e8543ad52c9aafc7c34bec931badf9027c0a64743fffe484c0dcfc39be8e5cf1a6634f999953e6121e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b3dbb2043c607ddffd07cccf37022a7290514df4cc072548a8d96fbade848758651cf9b37f3f66a467136e1eb1e0256ba5ba80d59e82128e7f9c716e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99ce27690493fea3d51da028f4a68084206a3ad113992204bf66ecf5041087aa6e7af6f31fc79a832114882534daf136c6288d699a31da0e0ec497a70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5368a0e124cbb03f96c2e2b0d0d77fa779ab23db5aa27d307fcf396535e50fb1203fc4f8704d9da31e93803a1e3ecc1db88e6526b4055556d382e6d6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacd944770264b29c67589c14c7c59bb59712724c1ba6bbb33bb8517d6055812d1d9995331c6b6d904bb3d376dd70b3709a56fce800831b23bc04a05ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31450291b7e09c67cb002aceda3433a52c88af046b667bddcbbdde0e27e28f20f2eb2c67fee3e3845929444c12a5a7517b3e627fe5689b5ca1cca51b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f1e71004666ebd08caf278d35a9c552cc2e794fb4542749bb93d5debe28b6176b8609bf513db1c792f6b1955b8858b66bfb8989cdd68d5c4e0a1beeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaa4956b8291b7e6fc351d9a79717a45fbedac4bd55c16cb83b2717e2196850e024152e239ceb53cf30733ab82951302b863b11bac2b69ab8982c016b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf080e599bdf6a62e1e4f5a2ce05c916c90516b37f34060fa59845e62e18ee30af6cfd1203c45688fd8d005a3b9ddb15dd3053ea110404038fd144fd49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2eda1f088bfa653255e379495b9c380acb29a99afe8ec4b41f4b539269490069c66d388939bc1ff0971288ea573be8b4f14248107da1f745260f815b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2e72189a369bbf4cba03bd585a2237914018d3fc4a9d1e266b305843252ed989ca598a936e4de4485de0b100a478927ef54eb0a7bf3763445d8d30b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4db31110f6b8024686f438af564e2415d4f2ba954c8d19ed64099e551aaeccace91ff05047611a3b33fd7ed30e8705da8c8404b596803e912aa72769e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94fada4442a6fd372ed025532f5aa61f4f75250a053526c19a7339bfd5fd8e0e5d0519d16ed382c65ea5dcaa5af0cf15fc4b04dcfcfa97f710a65c26e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfbf8e53b07288c60f8acecdca7c014d4f4fc3b16c2acc192c69950365b267e412a0f34556809d55655b7b9e3833afcedb567c5611efeff6f7e498524;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb89b948bc8ab91e201b8f2688e824eb85920e3157d6cb1f1f11fc9a5810c614108af84a5de8a3cc0e8cc2b80d7858ceef2382d5af752d6a7dcef3e71f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe230592550ef4fd7e25cfff3a7e0f88663746eaf2ffcee7f7066d9d3c3d30181fa3d8eb8c53306594fcb0da73d0b81d91040222b2e6c02628b230823;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7132d95f8ebeefe3ffdf5f8d644c38a1e91eb8efdf8f23618867f16a27a101e978a2e9535f4a925942e6b57978c20057033cc8c04fba206c5575948fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88a4b88aa395468803647f3b0258090a31e0b623e4c94729172d1aed1c238338d1534e5cb125d32366dd98a933b57d35d2eafac92c307388caff0131c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fdc3aa365d2846c4eb0a081134215091bd779ba2734a3c9d232616b4ffc297ea67860901c30bb63f2a8505b72472beac770714cdcc2248d83c495056;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c740a2a40f8d46ff8b161cdd27b6a7eaff5cfba6d44e2dcad4d085bc7486065ea920e0d1655374033df815c35c11a8b88ed2f309ccd2f182c7b7b9f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9829de6839903c52a59f7cace0c1fede0f99cfc2c6b82cba81aee1e787fd5973c520287e0bb6be3b71f882a73c3be0fe5130ba567e87d35b67cd26ce3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4392927e9078c64823b056ed316570dec3be29e70b9f1780e07717f1998f9bd9e7886c5d39cca193020672ce15cf04a3569cc23049db4feee4af8497;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4291d41e59265cd0eec13ab8ef8041eacb688815c8186be039c60ae1842fca012f02b1d7b5e6d18746978fa05858936e2404488f98d5873840b7682f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3844fad927e238d770403dfdd8384a1b41339d56e41e5cca855c51695785979fe26a7b8d14d8fdf333704b92dffccbd5d3b9ff5d1c473018dc14c6424;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac705fccefd95837fdaabb71f3d715031a214f6d9fb9843890fef798b915e5fd33dc38a3f44e158432a43263db8082dd8f29296f7982d2af40f3b67c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haabdbb401cdd9d83e33a2cf07de43fef9fbc53cfa38a54b0a6e51da005e76b26e935e1664c9d730964d263c5a4337f8e17bdcd5a3b6160a85856b3623;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habc347fe373ac78998ae689b2cca769dc0f37cc909380834b6d20ba5cad7f31c8c1717090f619b74d2f2ef7f432004462eb4fd3fcca68d7da6f173790;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6dbcf4be74ba1970f2f8df1b5d03f703bb02739cccb336e0f1dc64756c96e540fe4f1fd3ee1f7465d1d49d109587ae78d5635b6083274c95cba69bc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a95552c713040a3d481e05f30f1c2b13677fc0f9f86324cabc16b21381cf45dfd77326ede0507873f3436da30c64601a7614a33f1eff2b252c6e490;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h423a56d26769ec9869a4a6f244c9386f009a3f45023bd0fb82323a4fd46cf5e7fb4b755d7d5ce08c6376672ef06d8f8de8eb2cd9774db132df3c745a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd79c794c7d1f8d6bfa690cc973a05f3072964bb3628b5d90db35f2fad1ab5dfd6e157c3d581ce68fd808f26e0eb45a8ed842c63e9ef4763c37ba81c73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e0704b380645830e2574ede58130fafa2a486e7e734a80e76d71e8e68af0b3c126113afc10a7ef285ff74f8be6462906fb58404de46ae1b35a70be53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62a60793637d86b0bfcb9f12f0a48b94c6ba149a2530289f55e474fa35eed06bbdddbbdbce252b25e1b06ff4ea09a4c5a342e8aabdb66c627e082fae4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h675582496f1ef9c10bbfcd0501ecab47c5e600d1937c79f56ed27c55e236b21ec62eac28a353c71e3152b843267f8203ad9b507f9bbf7a5458dd2e544;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h780e90a7ce4b38db2cd373173500888a69db6f39a5c46e5ae2b8211ae316fc71d9eefc84a029711e2924971e151ebb1516ef5fe8808955a305671d9cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16823b02e23fc826b9608c2a7fb8641a6154d717a3a58bbe4a3c63edb006d2737b4995051a00fa38747b33e2de44e318832dea552389aa1a1975f9cf3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haced6c11a2d18679e298c2b7275cb340680067bde4ca8d62d17fe66b00fd51a65110ec3db21e9439ab5974881178d6fb744ac3e05071b00a4100c7310;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4e017021f2f0d312059de55013c1fc73046236dbab7167aa998108650efb9a9c4ace2b5d359a0e4372d1db2451b862d3390d51511769fb31050522e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d049baced6e77926910160a5952378793ba5260f853fbdfed73eb8de986618b14fed303ae2f4f63694d0f0634b9d2252d3c48939a03702df79a4d4db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2d0388f74946f6b074fedb7704fbebb9fd83eb61815054a9c6b542c2a395e7ff91ee1013e07a11e5b30bc050b4d3521697c941b9b18daa4be6b46b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ebc37695f3d7ca0e19ef2efab0b9216432c296027c2f47c9ebb5fccaf84d4674e3c6372fee12d11e8f394d7b5cb59e323b7455f3607261524cc58634;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf0a94d8e2b46653924c4ba51af440758f40e7b9137bdac7185b76a322ef1f3b284a3511037de20bc6cca8c2f578a20e1741f62a8dd6768e7f7b60155;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb89c9fe2bc70788b30dc3b8238687bae6be85695d687a127c5f1bd9d17b48afa78699b6c5435eaa8fc27370821af8f51468d3c8232a94db133cf987a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cb947e025fda8c9eaae007d85ea794020fe7f640eecf4b2092f2c406b5311faeba0b371609b31f4957576cfe4393234373bcb0e63bd5213cf816fb30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fd45e536a7b28c18141a11d8dce4ab5f98fc5bbd14146f8de37d44b31ad0e8def70f90ecdb16dcfd02ef16039f425054baf2cb92adc7bdd1f04d7f6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39ff794b72fb5a9f7e110ab91eca62a9aafa780b52f97473275e42cb9cfc09b7e8c9d4b417dca88a254f8fe54f902229c9f02b182126d2e5e24e7a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53756c933af34ffdc2b78b89a832d6e7188126fe37405a9b888b90e492422a7419aad95060962b5ad194d24068fb30e2900c2598e03ee2f1a8e2773ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11e83a504d4d5fdc6245c480dc561b4273497d0b1bb5b5949f2e88b1ec8343b46dc3c5c8982f7590842b1668ea663c24ba46a567917409d11e31bf81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7b6bc1abac24bf20736b18e077bf6e8795ed94c82d19dabb26533bc76def09ac27e2e78bcac38dcf88fb3178fff3700db77cb8de49e47c64d934c407;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9d503ac095a184c7649a1ac6ea364482b5eeb7c28d50c9ec644edb5e6f32ba05b47049d988d436356ae3df4870e59927a2880ee547cd292cca755e41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf106598e0462eb0f2e64a2706f8ed8b0669209517239b2e415b274b0797017468f132753c97b06089eafc3d6be27bcfef0f8e5b01c46469c0807872cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b232f8b99bc65794164a5ddfa3efef7cc12c48f819b1329ce83ad35a9cceb98eef439062d1ab270f738400b75bf641c6db45e8a6037e045af0df1c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9038cdd10200acf3df0988afe305cde0a3b9a9ee7e5294717607f0726b764eb80e42a052151499a77b3cb19dd7faedd9f0b23c7aea03fc181c9d030f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3890b77454061202690fb6c7f55d588ab09bb7cc675db038ea21c2399514044cf33dad5093912bde8b23dc35192014bfd1d674c4e9f05c84c7b3cfd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69697e6cb1346beab4adc697e947938c98bd9bba08600ee7f481bbf619cb7e7d5a36286bc5be2a643ffc1d9c652f9425c5e5373555313d20ffef00c8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d5dc86a9e44324a046435e5e61cff354b9c67d1e142d4f83035c94f834b08fe0ef520bd85a6a6f888482ae6d96e89d8285db23fbd28f3d490c51de89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfba9d95d2ca3223b49f14d65184259f56539c3a9941328bb295061e36f5293e28cbadd6ad67499f997e40e722a9af6b775a8291768a26740fae3bffd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1a3dc7d9240fce0f7ba66625983cf8d023f507c81d1f3ccbc9269656a57f73c041cdea18e85c94fc0c90ae8ff081b7369fa38d18b3f1c10f49d1d00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h722dba7e646d224a4380af5790005becd56f06039e2e4a17100a21e818d66b97189bfd9bd0a9d3c1e59e1544ff85c1a2457fc6804cbbf931fdd08f287;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fed38205911dc02c7b80930ec54d9414f1bb8e6a4b2d803fec2f271c92bbc04c90d8cda61391e0bc1c5ec413cd54825b3b63d6de1a9928d6f0018df3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h667aaf286a0378be3d4e6cc859bbb54c667de36cd32b8d5768fc95170e0a6dfdb7a3fcdf74eff121ab2719e0693ff317533cce04cf7e31ba6e2ef5e6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d6f7b109746eccca36fd96a4287466ac999d0402131d21c8216c9b80d70fd4a45dda553b7555fac294371238f58fac085b25d0a82de4c69dc0b40fcb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d61144efd12c63bf08b3d219de8977746e308f446a26f805c37629c9fd9e60458fe366475c1ea196c0258acf8d89d0314c3c147fbdf4cf4d708db14f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9c468d065164c19b2fe9533564d00ea382ea14efe5428c233f8bbf37ed86d221670bc029a6037bc55eab23eea290d927bf2854cae55846432cd3c696;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfed0d5f5a4de9125565d1ee4d2514ae6c0176ed6f0a0320cae1446828f42f6a76a5dc6b4f7d07d692ddea3d99307d40d8b3eefaf2eb012cf55adc3dc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8c76a9029e5d6c19b4db188105cf902ee070cfcda854b4994ee11e98d9d22e244837792f8193147d63a267b9cc7ed09576c4f5a55d4dd0938a67882a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59963c32ff9e58dc792fe4cf88340d661e4a28a799a5b440e14b9f432aef34f8e8646ff2a69177d149033a62975c20bdfcc4f76a6ac1ca49f05861799;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19bc35b886d6a6650dd52ef7479f05bdeb164bec3e9079425a75c213d37554757640516b66a055a034902ccb53fa539ca6beafe3cd479257711412394;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0a513a1b45cbace1362c2d5a17ba967dbc3922196a85855a7f4ee081f3f08216c561cb2caf674de4292bde32108d8d14b92e3da5ebb345960162ec06;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69595d09f89a44b6b025b72090f31be20967c351193db9bd9beef8186d8b825c2cc03d8885a856975896364f5a5b9105f6b9394fb5464f927bfa14b22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44e11ed545cb3669d166f199ca2c46ee84ae0038a828e3a5e64f5538fd586f898baf3545ad689346bb5fa6114f3ce2523ddb644abdd9c5ee1af705882;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91fbe9af504bcd35646934435d7987726f4d183a256ce115ce7873acec3d027db4e0ca93264b480ed50fd8339b2a68caf68fea812f3f180c4ee4d1210;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48713efab8726c69f888593bac50053714c524999e1670a310b70931f50f5019ffa5a80df217a268e637d3a32829684638699c70e8154d94a0a7cf07f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf22a8891b0d90413858211bc00c9c519f75ea1af55b8b2e401236b169677ab8aedad1caceb8357e24ee5c137a9d9954c7b3ffa719f4a6220314d73d77;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7baf61b713fc16f67dd04e1efdefc9e7c84559193f6ce644c1f146714e4af55d4ffee630af10fbd310a91760dad7f11a3db516d7d9c1fdbbd2e6a392f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7478ac9873770c7cf52b78d01b26b1cc43d944e8efd5eddea1089635989c6fe3d9e0829e4a0bcc439a45da4ae85363f0795f8be60728ec68d15ecfc2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93220237241fdbeea2a5c45f1c48681996d227e16cf5bf9a41ef4663f60b4269b03ff705502e235ccad7d88535d392681ffb20a188f07e979bf9f2189;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac3ec18b7799ede1f44987be3fb8338946b43b7d6f618f3d9e56dbd4e49ac9828397fa91bf9fb4bebd99d931637f50207167e7dda52162ca1654b2fb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha94f87bfa9b4553beba2c5ba6690feb67f0e9137316a93b6090eb9e2f7385ede33b2f6b5b1d6405b508b4e00ecbed5091cf24af7bc2867379a2f5a3f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcf893cfb5c732dc91c922bc95388018cd6205e914d9735af28af7462eb13c687cb7372dec85b4f09dc4cdeeb611b44455281c5dd2059ad6e8d6a4801;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde3941438d77fe44c8b79576cb0cea23c50e2fd00b6ec44965415235e37cf7a7308ba092eee94b81280e86878ce39725325d6450db481d46de0b028ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacbeb3b80aa4d7ebb38000348b69271410428a28575a6b901046534cf99919022bff05211419fa7f0f585ba4714b4565de37ecc0d7c56b7b1c6cfbf00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habbf47f705229725f2d964bbbbbd61de1dd9f7d62dffeb2fb01bf975bd3e65de8c81d7c904ca9b4c1b759552ad2cb9cbe93d3d190bba19bb2365e6c6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e8fa2be631bceea34e673a290a38f1e4234affdffbc4bdc4e894608b786c50e25d1a7fa617e923b75593625bcf9e5e7b655a32d8d308b3ade98fb99f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1901e3e7c3a55d46f491ce7009be998df65ffc254b692c053f811229e2ba999f4b6ffbae38755cda95d3b355c66b57d378bf74a9be5a516a74aebf435;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h187ef3842687ddde5da1304f49f63c3e0eba465e682f75c37aa874e427cd41dc7306eac07abd1015b9bc13717a364ceaf990e5055ac357ebfa2cb6a95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fe474f0449ed36b2053969c1cf554d0083cc4f9b555b1a4e58ec761400aa24f4d12f5dcf1279d90efc3ca09eb05dc8237da4ba80e036d32b0a0bc71d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50ada832e5ba96255fbcfcdd79a2714fa4ed6693c73f9f4b51e0fc2405db174074d0ce022c4519d56abb74dfead99cd9a41427e6f9f18a8aece73f59a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e667eb38c6f1772a722a31066448c5cceb2ec5a6abfe3ba6e04870900731daa264dd1e60a47d4b01821099c266bafd967b2f77982493813faeb088ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5be0c338b8aa2430f34188c0a25f5d6ea2c626e34a10823753bae43b39cde271aa0afe311ca44d2ba57b9e253fff7b4181d51ee64d2c8587390f11f02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96277f31c00dc05659d58cb4cc06619f7cef0f7feebd10c624169273d1f1bd1cfbf4bb046e3a053fb2faa456c4aee72cb976f3516d877a65b3111f222;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f427ff311ebb5bb47cca3497f7b2cb577ed3e41f9ad08f24caff787e9da47903de5e9bcb73ece34d56eb819c59d6328c1d2b221f8474da81feb7560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a08286a29d89e4e85e9704abf3d77f76ce7f74668cac4a3bd730535bdb56d6f72f4eb6a4e2154767ed426d45f774a89590de36b45223c06f2ad6c290;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha72a90a80f2c9d387ae348f7a833cfcf0fa906bb8753d69d6dd91bbaeb93ac4a1a03d09ad296df668575de866068fb8dced566807dfbfb8fef0b2213e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haec30cab477c6b12dc4eb133356ba7e00d9a0a42b80abfe205ae99c4032132c7c57df2680929011159c94a93e232d74ff4a3d611b9211d631da4ba8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37b72899e852fcd89eee3fa8c88de11da1e778d5ca9f67c1bb37b40f5deec0d42d090ebb68b21706422c2e5c90edff3081c19403c0ac13a8875499e40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bf3cfb72c386d4a0b197dd568c4b4a826edc4c37812054856b07b88eb42e6c04b21805413d0828790792fbaf476030e82a7acb6de15301e70c595182;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd808191e4e154cd112d71051a6485ad8db493a90cdd66573ddb8e16d0ac5f9736f280d0764ba94b0ec192e92b90c3b50daa361a061d288622a4f9754;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3a9c3afc6789f84bbc4ab199fb583681ab1b4cad5de8106d80b23dc86be73305806a43d194803bd556745bc137bde58acd921575724151e31c622134;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h967fd5fea9e4b637b4a4b15f42d2f99f51ac8be90083816a90cff43e9752e4fefd6502b387088a8c5d7c94d1eca1f72d05231ce6dfdc54536b643dbfd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0e4e9e4556ed65a9c2ebb38b8cc2f166328a770e34f3270f3277fd9f054f932f2eceb4a6575b6dbf1d0bdff393d6185e713c158339391884dfcc2e29;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h366f308beef0d5dbebddb5f0fc47f4d7a9c7e450bdd9a4ebdf901e709ebec6a7d75d9b049b13fa65b27c6db7cae00ec9d5130317d31a22954454fc372;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55e7e1afb9a6f2b5c606b1ee57fc77d37f4487544275512ddc024de6af1bbc76746cdf17e6a3fbebdab6b0266d532ee499f38349f0bfcecd421e22b6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21e4034816333d89f96b255ac11a56b2c95319c2e52b0e22376c614df82aa512efd17c9e21b7e6c9e613435ae962bef774890f65da9ce20a32c68f9a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h597857169d60663a8b2b7f2030dab38f89a5b4bab93e02a7c1fdcdd0b1990b4d177128c7e67d9afd41e053109d0848d5c84c459e471166342eeab78b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe91aca34000f13a32f4ac19bca2223e1b732d270ac96580e12fc20acff706a32f6a02efc63a59cbb316281fb840c11b0af9e92857b7a355c84569e0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644de85478aec08ea561ba40a0dc23bfe8271133b3791226fffba161db6e5dca57ca91c7d7be2360337126fb866b8708275f7eaf576f1e71faef909a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a23e2272021e6161fd3d4461883e133430ca1cf9290a7586b0eed6c4f82f429d6df3a98ff247f5b7866ccac796f3d3f9ed31e42ac5a01e4dfbe7996c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c31e2320af5a81cd29df1a4907d9b65ca63acba1000d4c379995c97e3b16c3b6ce3fa8ad2dbae0dca12ea7a2f6cea532391c5c4c5041c0d2afc1083;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12918991957ead159d3ef2414b8d982a89877419d1ef744c1208ac532700311192fcf2193dac38274a4a24c9e89f83b4cb5388376102e468b94e5326d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5be696e6640bc89e135b74b8c6f9e8059fdd62509974f3843c8cd090dbb2a0869a8a363172e442fab72b7dfbb71b7295899c1a2ab4c1884b18f89faf6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0376b3c60be3063b33dff7ef1fcc4b788a66acc57b9f2b6e5b70fe6138d2efcd1aee35f175002a5c57439bc310ca38be35ac9cb807c033a9c9a041c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd81ae4b4284222f071c3a099d139ad2b90faf5c4c3406d28e6793cabb4f542455ae5a114b21fe24d88bfe4c1cea6ccf28c6674330f9d3a3719cf99847;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59567f5262be66f7f8ad44ae2277e04ab79ddae021231bb828c7adfee73f0b3f045bfcc502ecb72fe2afce080ced91ba45ba57ebd34f4e5c1e8ef54ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19f9407ba4116bef0143f8f84a507a8941ae0e89214f22f17930d239286687189c686dbb596d69143757f0381e51803ee0ce20019778daec515d4987c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90a799838004bfb2aa4119b3afd57f7c75aab617a4ef1a5b76c7b64486f4eb4770c3661022ee38a648d734dec53504fd806b3db0e0f152742fbf2bcb1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c8a8a03a920555cd42212771c234416b5a7ba3cbe07d3f1f856f6ce1f0649ed326b6a128177b2b5e1772d6e3151c6745ad4ccc6579cc2a697fcfe891;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf724d6dd9f4ac1b3db496251da88f5fc577f08d21dc1cc06962843e46e80ac4256383015f1600b0fb05a2d4206145d5caa779ae1f02d678ca3625b149;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc5cc4846388e726276e8ecc8312e90aab9cc9ba9311caec9438ab2e46868e7af3b83453ac97b4deec3c7e017a9e1d538a5185de66b9ea12b341e9bac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed7a686ede07d55f78066263f69afea01b57581c4920b817da23bcba2c649636f4fbb6bfed9847df2fd4e5f560aa258f814aea7b36ea4e7a19d7415ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d392f3f56a61f55f75e57554c935854b99f20993b2c4c025ca6b8652d88c93ed0aa6b77fd44d69288a0f14e68d72219d8b289a79cb4b6ef27c550285;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82e276e43cdc6bc07ddbacd35c251e6a0f3a3f8f76b182d155598dd1c4f7d1b3db6234b7d2c724d05bbd972810b1dfcadbca915ac8a4dafe4213692de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf3e6e1bdad0ec11be169e947ddffbc120d4f58d0bb8388f22527d4c2bb0c78cb83d116ec1b8e10c1eed70977d462ac77c0cdfa0898249585c60394fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5252c0016e6cdd60d887806baa43c263c3e07d5a1596baa76f71a137d25709ef98444dc1f04e4ee947025e657fb492bcc00cf67207f8d16665058f5b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5d637afa9781d184953ce6b8851c878d5a144d1f16950ec4461c20e05188f7e3a39cb60bb024f7627860b0ce4d5ea186f800619e230857caa3ffd1cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h936f2c6655269af37d8c3f7c8c330cfce315bfd9f9dda695f869bb8bd2252c7ae811517f8e57faabe23f3a2fbd1fdef6ce6616f8fa0abd6811cec416e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb8b610c8ac19651340b6bd44ec02d16294286f9d312a99216883fd4762568efb2ccedd86948b61c3c731a4860a3435a8f607cddd40e771f607fe2614;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d49951089a3c26a18cf93d9f7e92db8d622dc291a7670234c3909c0f713472aaa38ea1654b4edde8d62f83b5e393cd8c0a9907adad12ec3c3096fc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h956d0dcf36c100282597b6eb1428aa4863f11de04bf68905b9fdc14c58bbeffd2f30fd938de13094547072c5476ba7ee336443c56f285aa444574a165;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1850d44ab9e3dc692fc1da039f0028381e9c82362fc2ae18c3cb53485326f2b30c0f1a53ebbe4b033eb29858b6fb9425f1b2cf1bf25b3a4c5121234e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd57d543026ae2709b3376a2d1ff7ea0b26f57c13ec4ff3c0daebc64ddaf501ddfd68857534c69c18686e067aef276ba7b29a46a125e7f058666776292;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc10c82c2d835aa722dba9ac011676fde68dc73f725bf7d8a903a3140b4096a35df7db5328d1455b6ce7912ff28555ef43acd5abac36f2b4a5dcc3a7e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5d7fb6b576b03b94e4cb5e4694218d4d1b3cf6eb2eb0deafb036d45b5c52ed0b078fb25f0f7cafdc0f68ec352cd04f6a648bd8d8aaa7274ab8ea9722;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2c39bc3bf8b690a97638ca906a7cffdd6a1ff898812be617e7a61c43a26f79c0cb3e790c0af2b44c62f1b5cf6c5a94c30574c3eb7da9bb78e6a4b3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3be284b13b470aee977ac91c2266ef09e686bf265adc1636c7ff4470ee2b912ef3614913a5749bc501737b1fa1f215d2d26615ceec13d125b8415225;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce771a31ccf7b398d4cd4e91ddc8a2b62d048093b0db983d9795243f4053156a55faacc2be525e9a5b189251d8a4cca8a5dbe30eda599677699952534;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbafba9175f6612c1b429ad37c351bd27f166216284cab67a8362bd6918a4ff60816c634c03d7223bf4be7d13c021b9cf6f5be3f8513113956bb70c34f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92754f7c6e2648c92c75125a01eaeb08e05d4f28f39690dab97beafc6eb50470b175857d651f722844ebfa09bb4a1543f9a8f6b5d63eda12994bb0bd9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc905d6a1a3e43b75169d97697e43b3df76e45a2632a4c628bf9172c810a49faf21c6318b641d926aed956bc822253902a57a63c2b9013af553a2de7b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d59df5e6bdb9b7fe5332d4f8623cfd1cb8141e040d6943e9a90de0f008b544b88876df919ffa760ad1768bd524e9481a167e0d97373744fb1f4c7762;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3a432c0bcc2c922c45a10fe55a6bef7a7ed0785f983c879718c1223204ca2d4b0fa398f3e54ae00987e0173102d1793b76261fd5d4cb3809bbabb69d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90ba42f5a9f4ecf751533cbf29d5b00dafe7d2535d233553c35bc2e53e7c46e88e85e1f3ea65f852c5e8cae008dc48b2b607e15decaa370416b4dd0d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h512116c9023d0a77504485c4aab4e2e698d3bbc73ee765c2c2566ac2d0701b2f4193c56d63a041e3f0f3c2fd41679911b8ad999602cb8dc2fad439e58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7a291d9bc77465dbdeb7910f8c911eb4e1d808d15d7b2ca29c8613bae1d6a952417adbde187fdd6ab9ec93ce00400b1e76461bb0848e078019b4e695;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e726f528a2629fda5b4563c234506ea3f61a3f166e7efd4b9892be241d6753c2c446cbaba4f5e27ded3e5ac85ff69b66faeed7e8fb5b618951c8b021;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d82e5105b06125dd2a75a108a18b070d7cdd23b866d026c7e9a7c6c85c24f415348e11aae1a875606ac3b75d1449f70cb9f0d4264563f168abd46ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h138c6a66143c1420ada99e3db38734f74e17547577e6804dedbfdf7bb091db6d648036e1463328858559908ceab6a8111ac171f04b93dbe47fe5db8bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h101474de0ddf336d10a56d6b038e85875acc087ed9bdca6962f0a802bb4c53af4d53e5f7228d9d4a0549f18e82dd15a4f0692e91b1ecd6a96a7be8ec0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2220209b908b7b6bd9b3f051d5f201d3e1ba692687e5f714e2cb83549ffd75606918cda124b43a3dfd23e8384f75b3f847f3c3bc87a2b332553a4b817;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2705fcee9f3d435a4b5a3760e62b2baf5eb4d4ab191828034720f0b3cd18b4f20221e3b56e2111c1359c5aea22e7d726c4303b191e33e13f448cd4b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bda88a0d42e1ca38534018234ffa9575c8283661a7494152d0e1870316b13c5fbdbc84ebbf258c35c8972aa58afee67bbd3beecc4f0a5c71796b30bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b7bd483fb7e80bf3cfce138387ab96086a2be6cfbeb559be8f679ad7234c6b6a473b1a9c18854302ecdf54863175a1ffd8507ccb7ffcdca258bf106;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec176e24365af189256758e1234dfd16ed84f221760a6b7dd4fd9df0f74e8b3b6ca156516e705d22fe750f3a1657fd9e3a5d37f361c9c4c3718f28ca0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9197abbf22ca03aa5d768a9e474b74b3edaba8cbeae7b34d1877ce7f97cabdb5160a4f6f0f3b465c7d87ac5eabbabbee1d0cca57e954d950a0204110f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h754359fdb3ae128d9643fba9bee5a7492858edd5fe9617b5ec7ac97f1741183916c0a135cd130241e1739ab154fe548649d29649df9a2c9cb2dfdafe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34ba13a06054ab0b2effcca7f553654d3772eacedacc16d5e717aa8397a823daea6ad1fa329dacbd03a996531d96590b8dc76388339b13bca1a5b2733;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ebd35ef0b8c553c6ee6aa82f7d28d40b43f05317f35b90f7bc7dafa6494d80604dbfcd8b031a0923fafa3fd9841af1eb85899b7f262929284787bf6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcb710bc72a22f10fc3094c2304cc380fe56fcdbd02513afff598f3e5734c38db4ab2c4ecb32f386a021f10242f43c1799e767bc259a1bae47a44c4b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae54ebf68db91285ec54a269fa5e071559678e9982062f454f9f9f527470b3db0259d1efb1b85dd3d63e4cd0e0667abc6168122027c5b820e008e75cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc67c37a04ab0769adc94b2714526f66cbdbf912884668bf149ed6fb1eebae4bca3eaf9a476c0b356587a00d15a8b976e7da7689d0a96d57666a145b14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56aeaa7cfe6ff3757b4b7b7132da392184e2f1b5f88fef27ca76926d582c442027853fb43d05c06b27e70ce3dfbda2be3f87cbbbdbe196defa37a781e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d80ad3cbe4ff6ab773c74350d3576df0bf7d96775ed0fb33442249b2fe915a8cedceae03557740447305a041b3ec4cadf32b082f7782b74c0c7cac02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc24f70a964b8457480e3969890558976c42feb6d1b6516fca3ba9bd94063e89a740f8a39a05c901dd63f25618128d4e375c8c838687faf74b6de8d001;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2091867bd625aefae2e6afafe3a2ac5b675994b73fc8e2928664dfe5756faa71d736341aa5ad450bc82bba06c24ac42081cd4f10cb53a87d2b924f7b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8ea7992683c29d21bbb69ac5d8bbac2e53e710065a6c27c3750355acedf68f4782b3e5316544978ef33165d9f17e3e910452417d0d637ebe3bae015b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76affe7da43fb0b87b3663b9828c12be6c3affe08907f14a0ec978f6d127697ae8ca94d5ef669c5891db7cf5749fd01679c999252c4385499d8aea77c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fd0a5af14f9b64980b391416c6190990cf185ed6569e5f4132cf67e0da2da2c8742733247240fab36645c26068f03dd434c8875fd3670fc9c739cc62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb1befbf3c564f504f267bc0bcea860608104c6b5df4a3bf03f1b5f3c56060f0ee439612ba6b6917a2c51177b3c139fc47e39eddb1e254dd85a05e854;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56021e41bc57b90171d44023f952315bc55714e023c32824ae32120dea42d2227b8f92577093257f33762fdc42fd023329212e00b817c85c934a583fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf69757cba1256cced07519d2005b71fdc297cc61918084b92e9f9074809b450f26a01e7b377d83da5c7dccea310d1b0e77d686ebff3fb4f01637c35c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd266ac47a99b3c0746a60bd2ae06233d268963a969762db98d030af9087619b9ecf9bce862382a40b820dcedb81192b49b40cd8971a1d9396de95ccf6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8987fd1d81b6b6d09e4b253380a710c6d0531bb2cb35a2ec27727d5182b20d100d782e24dbb583ff581a52859460d96e247c0033ab941939a3f041f2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5728a575116fc6dbe98f2882f25ef34cf3a6c0cbe9429d907f3d89a7f8ed34b6e23f7adad87125905627fb79507446c8aa4b8a64c0f98cfa73670b5e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2aac7322812bfea6baecc5198e7b0d0d72a674b6b3a202d9b8bb58a4e2f10e51bb460433e69b1506089233ee5c264945abad6869a4b6e0fbc30255c0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf03638dd26cf6c413444672abf09eb11ce1fef9e0f71e20ac0423ebbba127f261b088d5639398c7302a07ea657c8d051038c3cc9ca38cc7b1618afbbb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc855f69f4da1813f506986e3705a6a37118f597540f72599b52b27f8236cc7dfbc18a9ae0539c561fc186d3ccbc727e06098ac2f12b0bc50d0aa935e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf8cdc566b93f24e8996ef5ca79c77eeccdf9ff5198b4dbd14bebbb51832a1fa71865f7829d4c617e0e1a36995c94f1c3fec61123835090b2fad26079;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0fb799f736007bda3c6f6b173b0865ad5b444c63598fded966df3cb4306b4ecef6e1d2332dfbb4d14f4b3454624a16d1cd15b18b8150469491e63e89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f0c5af6685872137c5f03be76c444b2569c063f88b147b9ebc80d6983917391d2feb14169eca6acb02bd46e1f13c202ad37140ca116c4af6ef6e5c9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cc7750c54cc55c5fa8d477a8e5a32d1beb0d509a47d48b16b108ef8f6c48b1ef9fcd730c2a60c48b7ed81249aea5328855660970e2da70495edd5543;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2366aa04d4cfe45ee8dc7dbfd370bbfb8cfd6128b6763eacf53905330cbd5d0d47b169164ff989478b87ff2490faab3f1ecdebda489c282195d0031b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h333926870201fe4444c6ceccc472ab732fff784fe51c33b131eab4255f87ed454ecafa790bf5c605eacfcd68c802a4643b11509213eeadde2c5db4a0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb6daef097a2a4ad37f28d98ddcd47281d1266c321188d38c53961a797420cbeb6e7d351dc030d0d72e852f06032d3dbdcdc824bd3d35a6a7ac9866ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce59d9cf3aff6ee1c78dbe962de90cc1b9042033483e49b94fce1e0f03e30a7e58e1c46b5d802bf1cbebdcd66f645aa96f4e74c07ad9d5459e7169d67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcef2bbc139b909ff990499255cbf84b2abcb51688be69ad479664fd3818b720c6bcd293e62f1d2fc222c1df76652cf68eec96245337f3ffa6335b71f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c54b559c0e4089d9fdbb8e32926b2e017db5507c44f49b218e9b7aedc6960c12a9e46d6a467361296e40a67b3c9c1f4bf04e5584925e6e9dd4cb6ca2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d581895186e7a572ac591ea40ca95f1841bd12cc2a52f1d91f2df765b14cd37a2129ce9ab57ab46f0c93355a1e70cb5ad492747206fe921c804a2769;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6db8c02ae0a615295b8beb752bbf83875222054c07b010f7a4728de8de1590969fdaa086a4dc43e8d9bfa7fb3d1babe2c05e88e9ccb0c1d5d2565fd8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha93031ddb4f85ee7673f122809ca53b826af9f12a642fdf002d3f247751d51a761a969a2a845d3ea3ab63f67cf4cfc1468cca2e1882f0b570d3b08848;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd76135d1645057498b141088df64e5cff49c2275cb327738b52435a935664ff540307d3afc8afce09126f221c379c3c19adb4cf501d6c0ec9270385ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67791711a0917e4c1d63644052d3a2e76ad4f91d370784fc3469c50231c86bbabc049519df975913b01c620f80a8a36e0bfab83a57a8ddc6340894031;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d83a12ff732faa98ef25fd24b13596c7294ea609c4712abe501fe6d1f01ad9eeec6dfa2fd19f60a8636c26cf3ef009fdec3292c54972c11e861aac6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f33d0a0387ca220db38f9c7a9afaff95e0f39ac8c585b82216d37dc2e2d842e53a87ba2f8aab0a1a527ef418c8c5bb721a60a8ffa68756d233f94407;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c53e2c9598a2d1017c0593a358a0fc9aa7158cddc04c7ca845f8f4a2e63c894a3ae7e5d9c10e6302f83d3debb692615f950d890de55c2e133a235faf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5dfa0f218062cc8594816941a58dc9f218640e5c23b371471401e33c66b2d3aba2967301da0734469009c0c009b990a964841edbe5adf5e5dc1935b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59a08295890d2825ebb434916b0e37756cf69471e6c97bcdbaca7c0daeae788a09b24319341881226d8b56ebaf988668abf1d61922b7987d7adb97ea8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca899b66cb33aaef4a6a0e37af5a0b3a9370f6342f0200478825b10ee7d8e540b5a86d6b9993e95fa56a9c600cf0b8d3906713c1ff5b7ab7ddc5d39aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h396e3aa65e978400886bcadda76b19f1ffd04d3c2fb5cbc96345a4256fc6fd90ab535f506c5fda6ee7c279ea3936fe61b836796f0ca495927594e4c30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb3e5d0bdba0693353c5bdf04496a102edecab632d3f59bdfb6e3982155cc02aad60bc4829c9ecc38721417155883ea68f35d2aabd0204241da09e429;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75138cef1f8918d0d24a7707ccc8c207d49ddd2e7b9b20d441cf28d6b6337129a4c2a12a980d2c8e98e72fb2c0f1693952c5d403d9cebd677d0aa3fdd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c1bfc4422a2178615ee9b564fac4b9cf463543d6e075a58d1a53597ef53b4b1b8dd6a85d46164f131b44f4400c8a5e49bc52dae275f8f2e15e4a1335;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d96bc9bbea4fe269a5b9fd52c9b5c4e25160708d8ccaa7ec9414c39a426131f21ae9b4446df64718255c0ac9f9ac531ceae6dfd7fa8a801df99b62a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h316fdb01c1c51b9248fd985187cea0103cf1f05e33bdc6ee965a2f9059ac93474cc5d2e3e194a1f301eb1eec87aada411164ce8b27dcf949263badceb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h123f502e3220a11f1c94aeb422566ed08e99c7af1ceb2514139ca055ecc7b20268e9da0f016d48a44fe20a779a12ccbcb7d50efcba847761fda4f1b7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h893ef68235e1ff07ae16692ccd3385bf42053bd2f8cf59d36a8a1762087d39c3467864bc4754cc8a4aaff77d27a54cab3fe602bf2ed293828d2f011eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76e1c64319ad3ee96608875519ab584508940addd95f7d5879b45e50dbca32b307dbe4f1abc8b92aa70e9f89bdb8cb32796444f6d463f30998a99a9b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab5b3b32adef49b3fb2c5d220d23a2edd7710ec99e51891567c9a96ab76093117ce491dc5db771c8a992bd7de367d313bc2c69d26e58bfd0a3e8c01ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf26a409e8cb23679de35a71b26b30d226a32881014260d82e18e756960253a3702127b93844bcc58eed053459d56df4ab7afb2850598b05469ef209f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcbc2b54f6e764f6bcc5e040d73dd92a975e279f9977f3695c6f649f896be5b1eaf796fd7c152b74f2f81f7909a63fc160bf69e9201cd051d82a70717;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdf594bd6527b7847dfe2c646589e2712e7983543d2c7aebe3708e9ca4f8a7b09ad612a7d820b0a19e6193be866ba271d2fba9b3e77e0937f6c4f04a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3582007990e91ae27650b4cbdd4c07515b97243d0e15f7efb6bb9a6bc6e0593bc7a42de0db4557c84e4650ae153f35f34600f8dcd8496210fbba3ae84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h253ef96b2556c3f0b679b63032cd7d1ed2e475e7871460560f8dd1b3572e39ad3ea29e5503a81b0c9479b9f72205ac0b5d80937ec632d63de68f726cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2f42f83a52471d81d01af254936d2f6817a67aa03cad64ff411f2c9c5aa5e9e8345a433a22d93fef390dfdb884213d1c3d2f9f835cbb268d74b2eee8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8bb542d2583f9155e55aa452c82c5b8e32933ad389c30b5cbb9dad9b58e180dd33234cbe4a70a60239390efa5e9bcd5e4d6054ac840ea8a5e688cb33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb7a40233ee422933b7c0e22a28f26a62ff0566e04ea63f4ebee5ca492cdb99755b4e81bb99029d00da758eeff7d219526b5b5deb181504e726b7febc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h340f9fcc3dafa8ae771b290d1a285f2371590c03b3e73e5bb20c5f346ee76a8b163e2855d118699f5c6e8b337e8bbe8e071b0a0ccef5a38a9bfa10d80;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bbef7238a5d3c5affe172e2a594bfbdf00d924b509a5da3cea09acc4181fd3590e9b84bd104c0a32f62b6930acc51911faf32f4fb0d3ad0ac6429473;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3cabb5f50cfe5d3a6f3f4f6324c37ddb2bae0ee9818b9df1bb0845daadadf48a1d986738a7fe4c1d56377a021e7c6f75e3c2ea95c40d4aed93b20745;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c58bcff88fb87b50e5dbca69f1304b6ebaabbac07f08aab13af169978902a31364ef6d9be42c01d21ee792ee64877dcc034c29528aec53a64b7fc015;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7190b7419a24ff1e4350ce6124b729673916cc5c8b8312bc62390a2468559e077b7b9d30d888186a86b4bfeedd7b0b4a9b1080897bbd33ffd8c9c5d65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae77a97e53126a684e93f697c3bb639ce77721c63dea6563730d0d37972a089f699f7ff13155771e5172d70b4a08ba4b1659145285c3e09f03d9b8f90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a36092e36dc690bc3542ec3236b1f6e6155891152c3d0c2991e4e2feb7e025ff6698beb48780c701b6dad7b9a7fa832da14ce3f0aa1ef04022f9c2fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9f8c880990fb50606f0eead3716c481f80a92a7fc09500a6a398b63accd12fd6f1be6a56f06914289d1c99dc051c80d9fbcaca1ff5e511ef6d5253cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3b2efc50c7b70a5092cf7d446e4e9fae81c7956f1ea7bb06875520ae2c39c3fe59b7a847c13cfabf36214b0e1e4e332597fa3cfc28e6c133ed7f7a9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heabf061a161178f8be7026740949dbe3e37251cc3a5b01b30935792aec15c38fc1f14d4bae8a89571bd32b6ee277020e76e2a3eb724061b69d602bf2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h749ad2d0c61ac0612dba8c91578581111f8af5a7d334809a8362e560d05922529b2c7b0f444f0659cab727c0fa043a7fa67509efce7d68c32c8a7013a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc34206a71dfb04134473625096d03c77f414809322a388b138873e8c0c18cf037b1109868673ec80f960c1a799cb9ad94ed2b17915a454325e96d404e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7e47458e9a7657ded88389f0e2c7222836d0d0127daebaa76eccbff8bcfaceb7c73ffdd00efc5b8f2fa218e52464cd162ad32c11022718a142b28e3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e037785315ccbacc2725ca7ba0ece229c9ed07b6818f23565150596a1399039d7d236a27853094d2fb4264eb43d608b4691b97b6aeddf0cd1cf498c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c7351923d89570f8440862c97ce876d960b00d9cab3bfe781467a77d1539a4357729750aabe96e5024641c4e3d54a236e6c6e0ac9129f05fad45a809;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h827766c242498aba19130eb34abd1d8c3c7774d8b0ccb53027a40f970e012d561b4da76438d628ccf35f7834b32f362d0bb2b08498fb9c85f95445f1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93545b8a69710aefec4ae821cd0f6aa6dc52b86fade9e57e7c5ee5f9000c0f6808f9c41a4028b14dc08637af5224cfde9903bf8c202f1565d7b7706e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1422a99a8ad0fcc3ef60745f0563a82840fb675b4fa995feb55577078080853aa1445e1dbba674def923384a8f27c8f4d9f824ecb08b8487a4b0db40a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdf6a436199b52d5c53fa289ef2658b5f8c3873e39ecb55a9e6e113df738d60cad669ee149a20274678e7d13d01cceed3ca7bb557e33819be1c7eb69f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6239fd2bd7ab5d70a81d5fce206225b07676c15c581509765e7725b2de292b4d310bb3d8268efc9cfa05ce93056846abc42431ac1d897318929ffe717;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c37556bf7226803bb9304c657f1274f3b82eeefa9a90eb364f60ef84c2c2a86c15b48746bf2f7859e530d1b3bb51f813d40c37d7924db8c33795d702;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93f2fcc3db114bb2d0997ed702c817297b11709eb7be087abe72f9fc63965d55d0bf6b94eef591ac777eddd800ba6edeaf02b424e22f7560354e52f9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8871b559858c5050d209382e5d22c014a831e09619ba8018db0e9e6223d95f30f8749b77f61de3d499bac21cc39d9e82eb1a80e59cc992d78e239bc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5d372816290b3438d18a3f5f7e1776611906801246040342aae9a60134b7735194ef2b8cd8e5b0dd7b460cefb1adece57128493689df4fd6c072d1b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h940a0bffb2e682567f9ce1b0c3bf76a38d0effb4ddb383344a1986c3c58a9cbdf90f81f3c3d9354b72b776784754d644518070bc54282bbacccbc8eef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e63c9360dfecc9822d4ce827992d1c3c7d19c577f6a27e70e501b888f03338a7d1f9c5f1eb730822f63f8aa75d32b4faf783d87a9466c654e4681991;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h720ca00777060c625bacb2db84aca8b81ad3382979fa1729404583383fd46679935d832e95be1ec93ad99aee87fc083da4d9f8b22fd42153383af995c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34a6066ef0e822213df2d61dc2790709651a4a90c59d4ab72339583782edaf9546c8394cfedb051b171d1d26a614536b5868daec9bd26fda4b4664176;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h156267db7fa8f894d05619e3413da6dd0fbfa165b1a4bf5bb1729915e3b614e672fdebe392f652275a73a3840832dba7c1e2c2224b0bd656b018f0e28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e24abb9edd41884ae7c1a302748736ca6ec021c202e0d5e0e56e82500286f28ba90f868d7e127144d6376572f48acf6a99eb3e00dd78bcb9b74588cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b2ab149c188d272ebc09cce4f6dc6fadce0f44804f3c64daf4928a4b2a6577f4538200690b16b7b03270a4ae31b42024aad4a50276d6c8e3790151e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h465c8ecdb5c049871070abeb843484d0aa5fb3515dfafe5d8c0717fb7a753a89f826f5b7bbc92401b480d2f08d2fb0a8f44630ddb78f4c47341e77fd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e93979a47130ced7ec9aba957aec41558a498bc39f69e1c3d6a938a39a323c00af0b0c66169014d35b04e1d34d5b642cb815f7f0d9c2bb3093a8d1aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4013454a57913c504fe80bbcfc37996e865e5e7d9922f2265ad07e91212321d3ecbbd1ff8c254e7edf7e0db08dbc0e6beb7c42bd18b76a40db61b9f0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb14cf4a43f4a32f0653ac11140e61dff8e6c3b5a352b48099238f83d9e6b1b7d2fc6aacc2c0ea2dcc103c3c6749bb6142ebcc270e99f462af90efa76e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha375c4f9297493f3c6f45062ba7c2d86f6d8dff6d4839739332df844d480c3d86d98cab7f6b0eb612c3d24f77bbab5e5652bb1430d849c7d5579baef7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9deb4b87d1f29da2daf9e72f2a4d9c541b8626eef020687695b5d1f0dc149c685ff77c14c5f44a0252a636e0e58755faedd5608c12c8cf0dbe2511b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h207592d81ea52192ce850873907ce61d0809e917793158d2f18b1f6e372dab85d07328b3fa90b339a94b6ae026b72ef5dd31007f48a429c36f0f74305;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35c837c21c30d5b8887f401d3f5530a053e51276496f41c9f08d46072c27694974315ffe19ef8fb944bfcbf1d640536f26ae5ad8fad539aa9547f0698;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75a526a1eaed1a5381a52746ea64ebbd6ba3888e6eb9e5136d5e80b910a793fee12bec8592ee20ba206196620598ec4cd7971a36feb868afca4a917ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h151262e9779867cf2306abcf0397e8de92515d05555e412a1969448d3ab8a7cc78192b272f2569cca3a10ceca49b7c132a225380fc3e51108b3ce58b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43b4ac85b9c782a7b941c0dc758ef98960892ecfff2017c19ebbdead6992d9b93d49d3437fa48b27398f40254cf6e3a2cc919288450c917db5470b3e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea32c8fe32dc92e1837105a0a14e1deb734862e85d5828dba15d060de40efd68d2873a552399c14f9526d67e7c02d2b73c2d88694983a6f5b83bec55a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd35eeaaf38d77c36da91084d3109092f25327417d7cd70277309d12f09e74184ffda17fe39695040e23a858d6f370527e54f7c69ba120d70203ff74e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h142cbb88ae75662f4c530484ef7b55e53ab3d7f8a13329ac4d4a8ca778f6dcf26d0b3c332798f10851cfaa4dcb4f458df557994156affd785369511dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h278cb70007114dfd87c2070de46861b385bd67f0dfaf573392292cd2f18ce614c135e5c53a27d1532ce307803018ec232340ca35f02d85b5fd60fe8ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb7ada7788ea6b0997d320e56e6ead27652a297e7e70148044bbd1bd0a870691bc6d9faa8013637b4a402a598b5f9cb1a9d4f728d1d4887d575375e2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fab8f2ee10d08d10356df4a565a1f608f404c8fa256f8e8e7bc8570c276f0b0c360d8334fc633e9108b71c35a2c0fa91303afba1fadb74e4f16c5cbb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9df34d57a04c1033d43002767d12672c63913ce8f20c31432d8c52b04ffe22192393c7f6ebe2f1e2ed2df1fc14c8309da7e6a0610b7c14a00424696a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1e329833d90249a372413a5bf8daea50e4bb3e355714cbd2562af28b279651f378c6300c18736de8ac8603c260fe21568de2aeabeb796cea5b8f07b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee26186d2d15046fa2b73151559377e0dfa579660d20764a8f07fa6e9d0dfd68f0ad96ec6bbdca7c519afeea1c9b7267066207d73ac7bb4cc1abd0464;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2400edeb89fc60625fb4201b71df62f09c1e13defae5fef2c955f33638552392f34f8120efc61180cc1faa623a23e25a27c3a3e4365243c0f2a62f967;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h248f95845d3c8522bc933820f40ffcdf6afc4e07c37b2eca694a1c7f86d5a9a00f78ad26ffb64f2fa89d58c3bfb80dfd377704cd811c301085ad2a048;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e8b9d0fcd9da6a120e7793640f675338a154dbc7c63f4188893a7cf396ecbcc3a3c97ff8b0c7b804611591d6f3d5546eb0556283610eabeedc7c1134;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41da8cb45c2be8dbedb30347c20423ee85e9557bc8e8dedab0e3605e647c40482854c04e46b88229fbc03944890e86a8bf4d51c173a8c4982464aa6f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fadeea0ccfcf9f35ec85831dd76554bb6e9cc50910ead3db8ce3d39a74646e718652b8b40119d57e0ebdc5133d245b881fcc6f2c1118f4d5c61d8ebd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74406d4ec82d6c45d6ee20520921784cc53bce795da0a3740307169ef4e5402214f2bff07c6391df20ae32de4c587cb6e68af279bf388673aeb2b7dde;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1659c3ecb24874d53dead2e864113b7c5e936729896b6ecaaea4762d6d7f2b9c48f1ea5fa50ceb2a6a8c948401acb0aac613ba436f9c8211c1e203c88;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h119a2195c8afe1158628ddb4ddc5db028d5d4b7c86abf24d887e3015ba283607a28612f6bf6b4f47e4847739fdfe97cac68a11e062b64d3f45d309295;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6908687da0931b22640cfc2eb00efa5e711d7d6a8a27110a7a9e46728d7b848de48274345ebfb59d7f566c0dd46f728aa803262221efe0b895b1f9654;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc613783f469bccac69f8b5a5e7e8625a0ef41cdfc518b96c4730ed8e87af1187ee831a33d8b14e588ec5fcb869c5dde202539adbcbc8793e73632f8c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb50eb67e6f913eb8e04d074da376df1337a209fb3a01b4bc46d8a8ad2d51698efa22bd8d9daa697891ddf5e3ad7d202556b82275e2abc7f42cb1068d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b265413426150a4e26b6ada29588c655b22fc1d9755c95a99c9999ab1f60101c448e29c83e6186d7d7593f32cde1c59ee40ae9bb57ee7bf8a2397f72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h147ae5076ad855054b2c295d763dbec5d8b7d2275d313275c06b98acf4af36d46a00cbad298fa8b838b17ff6f07cade5a411d56c761edf3a9273dd8fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fae708fc7c07014ca1760c72378523ef676f7765930bb67e485c8a250cf6ad90bcc449ce125e3e4858cd75dea1e965be699627ac348680c8147d743c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e86c7ef8f870abac35dc3238270fbdf28d2f38732ac41f1bca27b788a37a55892ad688f87e667c55bcecd30157e87042079bde42de92824f88d5510;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf56d78a513f8f2bfe7d5db9d170695964f0e4cf01a79e27f81df82a30b377a0380f7a3e75fe033acfaceabcf8264ee04c1c0e914e15c88f2b8f78add;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f816fd06a95605f140482c3b104108c116a9d40ac22a8c331c196b7a1b11bbdd0155153db950bdaaf4ee9cbc074bbce8617392be6ea23c481713a79b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he465b33ece2c1ce9ef383dd0edde3e152db5b5bbd0e5d2fbb142863bac3fb9c9b7878a33b35fb0f079cb4943b54e5192417ffb2928af9e7dbef607de2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1d44339b66c881109a5b4dd099c5a3702a5043ee142de1fd5f170485652aa5ccfa1b6e8a8cdddc3c506e5b2ada853357699e0236f1cf260cd813c5ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7992b17203c537260f919089b788133bc3dbf98e4a8383369d0bb771296b942c38a6bb732d109c1a178922a96c7833a1b92f2b367a85054b31c926b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he63fae8a662881f92dace394fbad95fe61e4eef3a3c882b42d858b720aa17c515d26a19eb0e094ad797bdccd9061f0bffe4fa725519c3bf837e73587e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc14db7a0650342911cffa9c1307c3f64016ade1c3c26db23f3ec1a0bb97fcb107351e3042e1b104d526e80d01cc858e815dcbe5a3de7ea35aab4b3767;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h770f85a353e0144733e86eed81e82e9793056a574fac85846b4d615caf84742323215825bc6d348dfd363c3c1fc68f9b61d8ac5c0aa38895e0d230e73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52e9a7bc35674ae737af32aa4789bc858e97f0e258bbde6683341979bf1aff1ec88867154ff54b945d4546d692eefd76adcd5b58ec015776d3bd0f66b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf59918fb181abc3bf9b1a038d6ff05e38bf82861916eab7a8a1e6a35b796587a696eea844c9c4b5d0df8dba8d556aa979e04fcfa38f2542f96aaa861;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce1717b8c1b9412f49b0a7782c7e62d6343abb3146c70effbbe8736a0168bc2f8e76618d42deb0c21ebbf1c0fc3ebaf145e099516fe57bff0311bd7c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7dae38e4c137e811388c441c285fd8ce470863cf31e5796494339a7b5e1420f3adca7dff452eef209fbcabe806040f472abc20112e7ae754d1d05e10c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52cca55076d83fe7e5c5fce28485fff89e90b3d191c8380e63e9f920f742337d5b2f3e9a6435bb5da38302e056ea87bca65e95f8db1338cf8c9ce50b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf72fda0f6b4c06a65d9890d79d564b166fd05259a91ecdcfb54a8acd140e5925bdc1d8a86f7c1645faf3b3c35c50bf5811ffae7f8183a8be6c7de5507;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83760ce012ba20431085e14594fc48170cc2b361597df0434b7a0835aa31230721c98df18f8e2a8d5b22efa81a8a25fea4a274bf0159d0f570c63d412;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82d7372bcbe8c8693b4751094d9f343a9f449a5d8fefc1d8ed407de23d21d503548416e7cb973ecef8e99eb271a201e7a2abc5503e9cd66b40fb66f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58a51e866243062520fef29de555d17bceabff28150f1794e26ff4d4ddcaf5811abd26abec3fe274617a72d29e74a6d5408e51a62395256a60bc4b284;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2114fd8c35d3216bf950c2aaa6ae18b9886dc1dae919c1c6e668cf2273233242ff99369e41d23a7e4cb3184e0ac2f9cc75aacd0a5202505f89f8c9c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd81c9a47e55a4fa98cc713832286ee9c80b05ce4fb7174d8c8fbfb062ebcdd9c12f78ff8d7c73f983ad9e593a951410d6b4688b9afb3c9efd9038724;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf81542cd68bfa65c0376e3c2a24dafc895875eb348eed879ccf0c465a7b07ee175588f593b72bce791aa6fc260b958765c45cc82fd35d27d54c8c041e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h592db6345278a32ce9e78ca62ee4b43c7b24c0feb02b857aee294cb71d5215d51edcb289183b260a882885042173082ab6ce89ae8c5ac53bc6d638654;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aef65a3e626dfa505e58cb7c880982d32575c4a712ac3cdc7032110717a4f489480c3946a07199412cc919ccbfea011e2818d0a5b674648c6311dedb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5938b758f10cc86850fa4698cd975bb7780d16a43a18a3bea82fecc93586f6463073717638108778038e6b8c8637c60901d3d61eaae48a5fe7bd81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56e2b6e25dbf668765e3cdf8ccbb079bb493bb00acaaf3907ddfc6f3769bae66d8f4691eeca90c5c2048f5e0115c5155e70a400f0119a00b3dc6b9b87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf566d2aa9af9e3bbe569b60e1e116c04bca468bc3a4ffca7325f5cb25d53e5c2149209f4887be8e4d466b1210637f28b230cf0bff546967b9824d2448;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80c82a3cdaff61d60da0c78081b76f00679599a1b7b82526d73508106e50e811aedd0fb880953600ea8a5c8c8ebcf03cbacbc73a4fe895ac24c2bfad3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha567a6114bcb0eb5d3b2017eeaeafbe14e807a5323e59226d9f4023a8b28afd19486cc0ebb4e877f34cef6a119bc2fecbe6cc42330ca5b7bd3f488299;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he549fbc0cc891d2061d469bf9c2e86e6a1db0cae442ac5f4be9d4880383bfd0fa81d63df71bb2a155d7705347ee2034b3734fdfd2b432f0effbe19ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaa8850dfb17bd3e8ebae0cd605616c07d9f59b2723c3b8f18b740acc68e3a7cf7d2ef06d455bae07eee87eef66aace7393e87a69611a0f7942a40830;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb96a411299547a119afe84522efec64a02ba5a4fb2812cb3f9bdac3f9164ac7e7e50b776e7172576335be250a096881bf1d23ad872a65956679e567bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b91a7833de05c05a2d0e8de14bf746adaa42d82de1fe78a67e3f75ac90de12885ea756290913a096ba398b61b4706269273eb201407285bc03ce905a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde98367ca96d47c5b7ffeae9107ef5c17f3bf0fa7e983fc015c22f40816ce21d3a581a0bd9b5e523293e9f01bbe3def9200fb67c4c5b364f2feaad77a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61d14b3838006cb57308b9934421bb8bf51518815b60a388ef6e10d75da6346c3fef86f45783c4d2b022520a55576cb5b300fc841ddad8fdcae66ccfa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h845cfc564af8a94824fef099c71c278efdfc1e07674a39130e738d29d4828259f6a4a2f52842f3249f512bd33a25a1672566ea1b26dfe8087df111969;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2a973482a129004c0484986bf11130786db277224dde04a7c568bc8a22a44d82d4c1ddc8342c86f79bf8645c7cc9fb584ac950cce9557eef0c42c404;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h563e3f14f268a8724dc8e034cbca75eefb0cb2bf32eba9cb25c6520411ddd54a8aa92914dbe777f03f59b0f130227dcc6aa430341a2accb0a70e035b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f93dff1c832a08a25ef27624db6638e5a46a96e7f22e4d8db895f26791eca8eb95f417dad19221b81487b22aa0dfaa4733756f0af1c1255ec168319b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2fd0a7c12660ca97e7f4e626f9463da190d2c2d4847f6a3ff811741a6ae6f3f63ffce745ff1017dde94c652b3271aaabd7fcba70fd595130ca1ac9c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb763ec98d2634ded5e5e1d973a8c5eedffef35f719466d39c55fac4dbc6fb1c348aaf58737e1c2df315f5cac38c0a677072ee23caedff273850f140f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef6750e962728a62a7b39d4f8e94ee8410a45772cc8ca2bc7b663ffb8a522b8175b9badc157bee6fc7e753b5551adf043f903b3aa8a80121b71a0f3b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f279c2f2748c1ff4eca67060aec492fd2a7a27eb014912c7f263d03ec1f844487f11f8b2158447285144c07ae341b4f88b2a86e11da7a339f94bdeda;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he961ffdb4b6bc28662d40b5c7f26fe121a7529baac93d751a30f1c8b0f54dabb4c5743032ae1fb2180049e33a5dfba6b44bdcc2490a7ce552bee88393;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he634ed0ede1d1e70692cc7591f30f2cc9e99fda141277774881cca513e69ac7dc444f101f8b1b7c99f3420775ae7c8a30249832965fc3b69a7477572b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62eaf0fc67a3ebbb8466f38af054087cee0724cc641d5093afce7691a9a8613f9ead7b925738774bfce65937100ee8c502190e67ea5fdad019586229c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77c6cc9699c511ab4bb5419a9039387f47e802b23859ae989b62d00202e800345aec0040a01354bb1452ce6388bbb8568af019bc2e839db6857842748;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf9d99bea461da8677c4b0157e77c588d222ba81858a7ab69bb0b0072abe5e24c270d1b634439a0dd2779414140fc324f4d4e303297692eca32b7f968;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79dd9921032c8abb1f4abd15d6df68845482a3802a58c57866940cc56f92722eba7e3c419082e6b36ccfef1872b3ddcc76b6fbb80f68922d049b3d4c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a303227f72b088a5582727a7cbfb4fcf73ee84b6b749b127bf67878f71e4539db93297ea3ef776717e211115daf444086140efcbc7d440dd8f9d3a57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h370c9e132f7e7f0bbae29048df5815df0dbe4fdd1d7b38d1921fba3a3f1f635e6fb6fd6b40c33d856a2d675ccdb084915e1179fc85ee7e59af5ea2f8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h248b6dd0364e53a1a8e6d6a85d7a96cb62266ab6e6ed17facc0dda7730a9e04f86a53c838e7722df674ac12ed4d10feae71a5fb4a395d36bf412573fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haac56d84299cd573ec663d9e08d315958e3bdc569f5579d6db8c356ca6794671c27ee7be7fbb8fbd966b6cec016bd22b1884487db1435d706742d3d0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4de4933f2b9bc08499ee1d453f2456d8f2051f4d15d18dfee1be5569f21e3025dca0c4c5532c873e5ff4a68c39d044a0e875553d2a18e3f2d8f1f3c08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83326b7300336cabdc9b6de40024fd9bbf535f049a3d2804d0903219808abfead2c130b82790711af2ef2ef50da9da84cdd6d267e20b932b1a9d7f1d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7763ab9a0f6e6d2de942049eafbae1192b74c5a11ace940d8ee849c2931df7bd77c94419e52535283c72a56f879d82c2064b2499165cff842175fce93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d94c6da99f82dca88f6a39ccf19e7076330be6e17769b823c35d6c6ec3d6c6efd18acd6e3e94d54703ee38bc9f6fbdc04b4ab2535deecfb7dac36baa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ff80f16763bc8c2cc12e3ed461308d1942b30b69f05fbf7dfedb918bac9ba0565b659f7055d6073954fc9def73db9ae27eb7f94a0b0e3b47304578b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fb5e66ed2319b0019b45086930301a61c2400643b6f2b8ee13bdd8fb6be52978b8b0a7185c0ee23a4c7025510637f55dfa88c85fe1edb65693c7af92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2731fb2b7d946d7e3e32f5cf6efde418b97d9e75dd5bf2571c0fff8ef1fd66482368b98d3344aeba9bc8a8e95a893b1edcdc653b9b3815fdf953159f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb93e6e6e924baaaa47cb643487e399f9d519262e034234374f2f6ac9c792fd46e4e6b69c7ec719507a5552881f47b93208b41af619d475a634c8463b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83e44f22778ac4b1078a3cdfe7b5e7f828288ff9753822c08c3451871e2ddea612e1d63f0f4376422ff82e28fe34f6d8a2b9ae9231d288e789c36e54;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h720aa50a02c38273b1b026a9de40dd917abdf213e1c36335900e8adb007db19095650d36157636f127ef6cb4803e568dd800a0896fd46e7c7dcf49532;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90cfd8bafc05f905942365f47d573a7a0505e8aa1e5e81ff9a9100bf33bbd35e464cab8c0b49e5d1b09ab52d387fe16545152d5bbbfffe8f80cd9ec52;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6da30467e637fe768f17466041b030f1897082891204f566466e8fad25d0a18195f5b50e1c7168ffe7f355b07bfcfc7d4fcd29be29904bbfec060809b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5959c902654c937467c70eb38168bdd33d9cf8c6354142f6e657dd6439a49421378171be24fb8fdf1c539ee87f14af373088e75f1bc4e483a74a209f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h861670df6e20291b901b317a155d82b0be4b6a65a7378c0aaa7eafbcea215f72cf1199c19458397e010fb0456b5995d59c07ce0ff1e0cb0d9b3e75c99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5592e5254c5399e1b2dab53e69449348e4a01a934773494a3355f97484e3413f3f98762974c1e95c321fa1c2c3b89948e317a392b6c1b767146d176dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7328ac6f5221de1e5be9c9672e7c7344c9c8cdb8ca3011f9502fbc5bb081fe9c09242235dec112b6bd9ec083f2ddf0c4f88732b3ac041f6db0f591916;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba39065fa1d3f9859d44ce2ef92826da4a70d4a2641b490ff197400bc3b87545473f1cd620009910247518181c506028dc42155892960f341185fc1b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9028ce3b425ea344f34ed485deaf228093716a86959b4fc585d78b3d4f47d7b564d2b11eba1992ee9d74d686801a1730ce49222933dabb35cf592510;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45b4a57aa547ce076018b209a21c2b31039a152af7f2cf50e2536ab063b0db5f008bfb415abef57c2f8f2c637ad8b707bc5384475205d66f2184f37a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a074ed1a52e56a216689349be49148bd6773728442be922b4724f4c640fd27afe2f3b10bd11bd4ca6777997398175ef4a005c1970833569f206d67a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d0e916dfb89af000200dc489c459e330a6b2a62519d2c4608ad525266af58aba18321d170c813d082a3bd822138d98feae2e101df1fe56d7e90bdbcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h771edbf0b0fe918b9f49c19be7398c6598e54fe74b57650d3a3a4f59c606bba6ee219e27d6a9d2288cd04d1ea9c5cafdd52b6040076428391057a2887;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd9ebfd014e0d1bfd1faad4257eb05275a80ec0deddea6267324ec62bbab715e83cf5d9a0fbca8713a2e688a1de26f5c0d2f413b05dede8671f3ed334;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h626f28f97ca503c7400af95f2af40dfdba19469ab961a564d81e97cfdffe128c94c98765b605ba9939fc0be509c582e043d8c3688e6dcfd9103008c9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcefd3bd5e2f98d4478c9636e0a4d3ea0f4f75f438933823c132c114009c6aedc365f5666f7eebbcf74085243ac537569a1ac21259b12e99cf26ecc401;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heeaf18983aec92ca60be75deb2ab68f0f1f32e3e8077f8189eb6fc07da2486aa40e7b28a29dfd73e928a60e1c1f60cdeb7b8776dfd05eb061a8448b5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h704e04249831770c4d2fbae4596331e06d08df1961119a761d0bc36e35ab8b3ad9ce725b1179ad0dea19e70a47a0e80b3363bb4504b8e6fee6fab4e6e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9caf134f7b77128108e95727bf2a548fa8defead1a3125926f987f236b6de3d8d644c0132b31e3320ba62da8e09bfce7112139243e25fe0056a6a87c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61bc347e7465588f66bdf27b84482238e3562571460231dc274c2b0ed2ea89a2a8ac0c35aa7f272631377729928581417c03ccfa884a8dfab536dc4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa2e5479755be7f21b4ef6a9a6cc7cd14ac35d353dd3bb534f604cc3a91711f281bf36654d1ac308869be080b1e4f90e2be5c52757f79b70938dc90cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc41b1d8cff9d59eac791e926bda42e8252d2c04ca9148bea615fbfc43bdcb8cedf095a12afa8b96e553a5bb8d8f33ddeccfe51a906e0d884d07c98fb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72a1594585d22add87362d0301255b16272fc48ef28ff08f353d5843ebbe063685b43f1e312886b5439468b9602e3fa50c02029bf7d72e1c82ad25731;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5e75d11c977ab2df19ce44f8d06d4232167509c792b1a69526813f734193f76f8b116f537eb15931c18c02973ba30644f0aca46a83b3932a95bea386;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e57b1d669fd6a1c669b4c9311abb417f375899ffaa6d07efb515c565e994e9639efffb39f8fcb69742547d92a0dddf73613b0b94955e07f88f9255e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0b84378c1fe9732d2a91d6a187672d5a6374ca3cf47f8b10460598bffab5eb76fc57b9918db16a66a863ba7aa1fcc1ffeeb93d7ddef6cf8fefc52840;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ee1c80b6882a58d6555069aefec73d61903c594223a39f58a2e37f75de64bd31a21ea09911b6c4f4ef6ed3ae6f64bb87a42f49dcc3d3ef7ae1612d41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24d110baf1afa4a46f4496fd22e5e06bb9d50528007baa09f303eb1cb9601e4dbfe6249ef512cd0845ad7f3df59a24779cf4013b1b84b82003b1a0f6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d330a45b0d3b384cb503975e37f7dc40d63461249cc72c504acdaa66b67224e8712e336aaefbf34e6283f0e2669092d32da91199eb40cab2199aa38a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb810a71e3d2608d618ec19dfb7f60c8091d3cec6055016b595f2066718fa1c8f82e10dc88ba59ebc76bc5d5e01b26f11d3a4b8d5b4dbeb7aa4e1b49e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2c3b08edaca2fdaa702ceccbdf4b3f849e6484921bd7c1657b771cbb471173d12da571912a8dd14298e71b07e91c9cc275bcf2c6ce0be6faddef4198;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39457bd01cb2536305426ebad1ff8229fbda8edcafa5e087f096f67b0b8b1681f24c57bb7b5d781b322fea8ba9d9c3d5b15ec6e340c0b5b46ff3add27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda97b95ae89494f5ae7225f9187b6cde837bde4c12730673ab2fbff7d85ee666a29c401d9d491e4e9925758772476285be9d13250edbb2aed4401b37c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc747afcd7eb1a9b70da4398596c9fa9a8a19dde7b518a6a1534c26ec1c197f4c94de8b78c167a12a21ad66cc2fa17efc27419c5a567e6271df47b280;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haad3ba7cac2fdfe6c45535609ca05dea6f213837fc5469ed04c6656d98920ce3b074d5ce0c895c27ebdeb140f1712b73c2d6bf55bdb890b959f3514c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb855698673da4bb63892a9a368ea83504d4060cef47488268023902cc2d6fc600f3e74610c07856c73a4d6e0281456e9567054f885f98bf2b4e6a47d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6aa1cff9cf7666e4713ae1e3d98f07ae484c36f48f7c64444602fe2f43afa3f216adb76cc496083fafc86a3f48bec465e351ae67b1beb4edab20bc99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h243dfcc39b1822ce43ed61f57e327c9af11f0190e57ed070e3a18c269d002a8a935b1d2e084ec1bd4ea18d5345f4d1a120f62ef91421d5d85bbba1d01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27d912b04532ff958638e598c297f2c6a82d9f61d0ba4bcdadb2ef5c8156408cedbd6c7fb33b4cee151fa33773db0e10e9ccaa68af756a3aa241256cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35525f58cf883ce26061ff3280ae8bbb80ce92902582353269fa906ff3c906c6fffe0dd6de60c3350bc5d1282d4b2761745c3a75c1cf4a5204c16057d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h525a3893017f66bfb1a1d379957e967752887a685e24f884d81213f554d9e330278f8c4b403255c4ea71fbfdd262f0014e59de667577d2315df922613;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba206e77fc8142e982f7f25ede69fa38c30b61a6e456fa74e6ab66308d4c377df795f53be9f80b2e997b0fdfaaa50be9adbd7b4df97fcf9ac5b26cb71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21c4a1072944b90ab1f8541ef52f7b272837701ad1b3e93af1e6f861129e2676292d36e7270e212f9aeb4bc2fac1ec25eceb2d48810357d6858374d87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h242d4ab7148dd227e2c14225d120a36f56f48d27a23a78131595ff27a1330c9b0a55d9a61400c4781d8efe4354be90451ee238a8f52207a060242eeae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h316faa794ffcb30e9f2dbbac1e0ab8c76bb1da00fef441570a74d227c580a1c324fc0594d29f27f711cdc449c8dba229dee951d894edf5d935324b5f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd108fc2ebe81abc7af70ebc0349b00b045f0ca825070b5de25e9be452436bd891815e600abb9568ad75ea16171ea7afc0a976deac720f00f37b39c358;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fb274f58dba0df2fb5a41e45063d22befb31cbb6a1bbd6c4c5e06e85643a6c6da4f255503b7ac7c6429ebc6ef77e85822a356cfb3c07709737410a4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64764543ade62b85af5a363e6111335a851741bd2d1f0c73d83f5d125fa8dc5d7f97649a86caf04d317ad309e20a550b3a9b4573018579168bc41d939;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4892fedd81e9444c14ed2a8cd7325febb0408c4a3becfc173df1f06f8181efbc29c78af952d2574a6cb6cc0e6ef25d2cdc0f61d88d962037d329f11d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8bfe67a4a77ede0cbbf8a703e114709a28f5f5e7477612cafe9108fa01bd29cd2846e81f2ff27e0f70055b827949562f1c1dd9f432891dd4b2ff2ad2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c736455d1fec2342a000f033bb88a85993e98cab9b1d8b39ce9629c903e21a14c713c3f169cefb01418f6dccbdbf809023df45186cde0203ac777e5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h623e9b5b27daac243708d9727d611442df9a653b393bbdf6d668714ff84de8f2b83e1f70a937e3d01af1e21db819af44a70dcac51bcbc8f36767a9bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacc3dd5dc6850df140bdc0b65a897b36606bc71f2ef820a29f4c7f934b72988c93d14be2c6217800a79812246a0f694356e33450b9ad9609fb742d767;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h245874953aaf8ed848e5173d7216045a6aead4afd7b3f3eecbb34d1884a2e6f50c88af955fdd4de1d0a225221dbb97434311b63b5ab3140ff9e6a80e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbca520ca6a2976c8b10cfb1aeab6439dee6e30b6a66aeb0a4e5f294c0e0e8e611d151044bf7a38816294d106a6a0b4844203a4e8d36546ed413ad81ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e92f1b0d36fba74a890324a76f6ad43805eb6f959a71f42d8e9e212a07767c00ace6fef4e0dce02a0c8304c5c96becd4756f3fd97ae0c87633a9b060;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12f2f5f057ad4a2c8ccba8553a271d6076255688d70b3bdf2503921ebb0a83a704a23eb1620927a283db5998aacff8fe7a934a002b2a2249672e2dd37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85049d2f92a0910ae72ad4d3e6dd8045cbd6098d1f9530401001b57fa05c25941291a57f2bd119e7b7ce2ce45544d8150e239a163bd4c441faec38aeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha23b9c81ab3316f86bc8f3d42e8c76d3177515d80d360f02c2e99a730fccc334d0983188c12abf1d7fa95bdb9879d43e7d79bf31066ff848689e621e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63ee4179114d5acdf2b9ff8696ceab47198febf992d1e4efebc4557062589370d359f419197d32e2e97a52f875a504f50f70bb388064914506151ba3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c28b67fb0d01c8114bf067141bb5661a471491eb5c57da869b677836a227579428feedfb5d3af000e4927d05a6550fd023020fe1029402b51ec1860;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d4375650c9d1a97f6a7541363af7b3b0a324e990c91d2dc72afc0a3f384ff7241f3bcf94e6f098d832701b8674c81f4bb7dce099f0cf27e78ee24cbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3191429fec378e98c99a12f8f62ddd65c0acac44387975702840b303507baa8582d4c82027d15fd48e7f3b653f17beed728f23436f7ff79a0e9b418c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfddbbaf4be8edf9e6ede38ff26fb3e9c1009ec0e3414d12e964f1403bf826dd975f7bc94575a61e7540c7a6cb99dfb00f72b886d60bf25676326e2de2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7451484e6776a50125743dc39842da10aa510e7b0367bc0848b43085a25ad9343ddffa4f4571f09c1ffcba4ac1bca099e5e2bd7c512f7974d16c01a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2cb9e52e87e9567b35cbfd2047e85cf8e1c91f22530cab097b5e6fb746030947b12490a4dfe2ec6524dac953fab286517b2545281988b4856ee6a0fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc02af01fdb0bc97d8882d1830983f5030233a67cec8faacd5891372b2377fab564d09f68fe9352767dff635d19b6fdffcab6d91c16db5e43aad7f4df7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc91332b72ab7ad93f8008c2d764914e324ff8810074186de0b136fa297871516f5231537bf78ef0be8172c760f7ff19cb77c4edb0a3293c3126f0b967;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he576c8efad7b32c5284814a693a83173e69211b69f4a76be125d4d79fed4162f60e5ad98ea2142e1e047755ab1d0fe6456b91106cdae3973343ba1d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d9e70ee0f1206e5acc190ad7ac322f3ba1ea03f3f4d379f597a04f8dd1c1e4d574940455b8df7f075d9c707c52cb62d97d2421c0126a481f502e8513;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a2a20d0c21bd12c1ab9ce95eafb5ccd00be955ba8d1f7afadb67f82cf5d0bf4889577a65256482886f368a4deaebb844bcc2e0a99be2b95ee6641961;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d1392f18dac285a4009032cd1693e5eacd0dcd38bb7ab9b306ba8a2fb8e793212c8ee58a01d50b68cfdf2ab48eab6d31ca56dcd48da032de8abc6475;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53017c94e728b3dc5b674094ec5e6fb6ff4d01fa7ff0bdd776a307905495946cfc47e811ef4ed1775c26910d79b9128c4b0faed054e0635ae1022b5ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he60cb11fc06d1ae2debbcc251379c631a262a8b0d2884ae4ae8a74a6f163e8865a87d20309276a3fec017c564392f9fb9fac77d6c09e2de6154b525e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habb30871ce6d7df1a487e1b52f96fdf89ba2256b3f9dcd1a4c539f81f0a18408873a3e723f38dee505cfae75046ac2c297eb677e9a820947c7f4cae1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h309e883ac77bce3563e3b7636b626bdffe7ff0830ac9456b73fb6c9f4efcdd2bfc4d4736d0170f4754a9728f06b43597bba8e1cbb2410bc92058d87be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ea26778d51963ec51fc31460457016eca435435d0b54d2b7455064600c7ad098feb82a31a8885f6fc86146804f4d26f8c3ea91214aa6024de29cfc26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28b1ddeec7944b9c575ec71502de517739ba004a54fa2c0bd4805ad6b84d37b997097859f926ff9d1f9ff3f6d1dcd0d199e11abe69ec269108e0788b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h570c6dd20781fd249a4bb964fe2d9eeb5bb1ce7c46265a3dd87bfd22948014d6ea43dec02feb01b05cdc903755da172cc6366bf2b36d7b75f3ac236a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6916298ecdc0c0754ff8c1f7d8c309d3fcbfa8c26849ac89d119e82dc36e514cf83ee1091deb920150e5e4800e2c42d6ccefc7e8be51c747920d686a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8917e149d97df6b095ca276b5e839ebfaa82dfca24cbfd921e82bf24de8afa0379eae114058f8c4bdbfc68fc7bd665baa135ed18be108055afd57e6d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9508db6f5551bbec328911050507c70511434e38a9395b1f9b712a487583b103af14568057b4b8cc5e065c0e6bac2b49e6c196c9fc4dcf03af39db194;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96e177ccd5c9c2715d40ef11cdb1f7e5a69f14394a44102703e80b77b925a676812ae31ea180110c8ee8ab7133a0d3e460fbd55832acac82bad5103ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fec083b0da98872e996e510e7368cdc339821c54ad8f34b946c246122688d3a741efbbf30af47db1294e14e69676431c1eb3dde89642403e94825d25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13d8d5040c9de7343c3ef5ebe5f975d1e4fe9be7c926e6ffa29b5b508089c9aa224a02c524b26d0c7181696010565d6425b0c14dc552f02d6a0e40ddf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79ab31651a8512a108ef1de202e8b8d28807d1cb34ee898e18ab3d0835957a2be5bb8546e2d1f155a05ac6745d4c3c776a267ddf3eb2cb3fad39e3555;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7391ffc92ee76b326f1f37e1e1100bc01c173bfc092978f5c1f194607d1c7b6fa65cd561e0d8a098af839c533819e8759dec48329afc61b804f7979a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4a992d6d972dae7f155e7575c1c895eefc2b008fa0c9a880224d43695614cf9fa54c8b40a483769f1257cd9153454e7171c2295a04391a78de3a6487;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59d017971e926f38d46bc36052c0ac410aa2f5a239b39d513b9707e1245771fcad928f8cd959c8903ecc99cd0aefc6f38ad9c9c83ca51c81bc9515ba8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24815d01de3f66de5ce841041e003bc420284ba2f8f7c4897bfe4acefb16643689f793a1aa5348b493b77efd4e2a7e1cafb8b390795864e748fd9fc5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fd3eb581f8e041a2c799efe0d7d1338b5195b227cac2822e9ce87ed2af4d58d35a3ec680451222c5e3920f846aae1e2b05f9e2b6d269477504af85d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7abe990335af5e729203e8c97e973d9fc25af4d89750c6098de3406bcfc0d6643a6c43d48671974d29687b59e1926e70edf564dba6c76850299a78803;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha23b6110f94cb7c38df7430f772775fa243358051f9483ceeed87fa996d27ec604ecfee2f70a324ae1236034851e69334e797a7ce4e04e98a2186faea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h971c581950cf8168a2e9820c52e5d11a6cb098931918b2dcfbc8e7bd5f0462b4d4de75211a995e9b4e59ac22dc1348e9a9a38656889649036dbce5a84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab4420cfe33204c678754dd6231f555792ca47fae1eb3bea75e2a38bada3c52245a2c68ad28f32de0dd7955cf13c7bcae0286d1dafcef93de31768e1e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bfb1134bb5ee24d58b4a5966979a6f12b99bded68d74ce15a0b01fa2c898a3ac234d531a594262f38d036d8fa07ffe9f783f78877e5941fddd2f65f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h261b6708f1eda1f112de6ae288ef88c19fb59a8e1e68193cc3287026ed9159a2f9cdc6e5639f9c58eb7061d36a606821582f37b52a3ccfbb1364ca2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd27bc959cd429b38a9c8de59802aaa445582773b0bcce112c165a650442d321ab06e91e9a452d9b37c100e5e4356c721a012b0a2c7e46c9b83e9eb0b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb8e89a1f884bf7ce907f06c78dc18c4db646eabe3d55c3487be48b75fc805aa6eb769207f95523566bab23ef6850ac4cba5223ec2495f8347bcc4990;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fea8e0ec04b9a01016d946c1885fa69cbddf2eb04d8c9c7cdd44805924453ab5bb7e27882cbfff67e1542e95c2e3238cb5e15c9676d958f39eb2d7fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ac2199bfe2b04073911a44ce3be2e265a4c366650084b1c9fc55983e05b8d68f9b9f1cbb9669b823e308364d0d3611d573f05be354d78d551bc27d81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5b603d9a6aa83b13bef0ad6c8fd37a330c7488a3f0005c5f2917a4b2cad91cc13b23c835a02a97c31da16a08b2596448d970160acbf72bca73cdfbcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h619abe556342cc29fb0225da538c3e86b4d840ff1b9ada16cac8f2c1e72567fd06e28ca6cc7e88ac9842fa98fdc44f4d78c22a97b121c544987ee26f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb77e19918e99388c529f1ea81ca278f39f48f0e9b437f8a0a9a86b9f78fe57d85f47ac280f2d12fcd8b97994170f56171c11db5cc27c77e0e54c6e3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5de8d59f4e281243afb819b35e80e6175c72acc201ff42bb3db101e922cb7b542b2c3eefc9d454a66e0265b165914d428244d8303e724ce805a0ebf17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68b41b5c2bbeb557f7dae07664ca9f2a2e3521354bf43e3275e7f6b60d51753fd57365a6b9136a25bb06f7f371983bd4e9fbb01df5249332226126600;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1855d0fadbed3984dc93bf8b24f9c992baa1dd458c240516f8b5918eb71294a732167421af78e86fc170bb73b67f2f015a197dcbca20c8c51d100ca8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd082727f2c88178a5f6cde98752d8f7fcaceaf4ba91070a8df35ef389ee9a1fb9a85a416b25eb10dab48906e2d8c4eed99fbe4ebc99b2bdb3aa0fca6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed53cb75aa6e7e0022f2696b855e2264183efa89a2aa840dc1a86b055df876efaeb2cce7ca6b3a2d8ad8f355a246abe69b3e1bb5bd29fd869378589c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7816c021f8542d7731e4ec91b3ca19b467f49e0020d3c1619289e05038f95144f55d9e116e7d49e5f708f1b13de2d50e68f6a576ba937e196011cc59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc81a39de212d4347b0f8bb266650c8210a6860e1e5363992cba2afcd99abfe421a59fc2e3879c6882d728e4402d27924bfcf3f89ba389cd1297c2815c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h327c246d1cd49122b6e5b04ced6cac388265992f2e59bcf1ca864523044cdaae44a583f7ed74d7e0723ad0ed3d0906a5aff0aea1d68b493af1ee946e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3664640b818df8ca9f7cc0ccc51834d01796fc802d36cc96bb61c2f1a216d60606f7329220e986cf348b2d01322dceb2e70df2e00345f7b3e35645e65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3f284402b4ebb45e8189349788525f77d6b86bd12b96393a9c21caed1a61b028076c80d6300acdcfb5f93b4a9a60bb8c7751121623bf874aa2b1e6ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h521ad88205c31016eeed23fd3278adedf3b0445b0bb8bd5f15250e0e0227369cdf3e76579952894adde10fea6e0b4b8cb1b9969846dfca7d94c717488;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ab02529426654b751d379eae192f9015dbffac13b1dd5528eb610ac4cd4a6137a3c98c6c2c896ab154187c0347256d805c039581eac3de5ca185166;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fda3221f93cdb35b98a96e4256ac5c0dcbc0894b38447fd1922d23d12d0f376b429cc3dbec4d2c1055c8574e591788cbf21b064bde978500f37d784c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36316104865eb3671c8b3765fe5e13dfa00b7f6f5c64d29f7e51b79c5199dff8661e8adc5aff675ea8065677628784e346a6ce5809b5ffe3b1967e981;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7668864d7a1a0fbc47e0a3a161f60bac41cf73bd9af5238a5ca5b6c9652a190631dc83ab70c8affbdd99a844cd757e0e6681a9ae3941a45344ccf712;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed2580b4e2ff397dbd9420199788dc54f862a357727b476a0caa3da7acc874870f5fc8d6b92dab4126ddedba17e20aab852124801cfdfa42907df51c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha30fe4515a4cb7ddfacc3392a36a17a971affaba6dc55d6c6208e574148cbe87e81913f6c74016f0397eefb030f845a8ff8aab4bcde02ef083e1305b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c2375e785ae166b64ca2784d8d4d8701bcb5833681c109f290fc4da409b0ca992b83a44ca4f558c06a5b7930e573436348f9dfbd6e3a6773c3b9d3c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d9a09415e79451d962cb95b5ad8e65dc195a942ff07d8c4b7dff08cb91c59e94be32aff10c2356a3eef87441739c3c95ce15b3bb4a1a273934f1f4ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5007a50bffaade0beb2962acf58855524fae5ec85fb928ca516bf7c53510989fffaec85e6e0777ece305957ee84dc68a82773fc59faef6c126601495;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf52eda1da830a5916f622b4e243178de03ef9f305e1c0fba35d0b1de779866f16f3022af5b9a4977a852fa3ef96cdc67b8c6d3adf51db62d95f627eae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6acf56b7b15e0461dddc3f4f0f87e7a58dad64ee4f20a12a1574f8dc3e8c357628f4332466496735470bf93c935d005264d87754950a175018becff8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2497259ea0ecebb1a4cc76588af608c78a7636d80eb64fa785c44cd1c809edf690c8250b452ccad418756bf9b331a5f35192e8f6651ed0c29eced615;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13dedbcda4cb07ed98c111c6ab9347bf8d8889d10685db8e3d029c5693b3153bfcc287a812d32c0d8cbfb2da67d23beb49430f4447fc6baf9108668b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fe221edb0b31a847c5b18cb6093605623d391918f2cd19626a9a4b975275dad8e8a4158d7823127a1cc52aa7c4228954e80f66da74c154b5da126ae1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he36ce7b82c010861ff3cf1831008bd7784264b69c8dccef17787fcc441ddc5ed49206c90a7b8191b2f663450ed278b304aaa465e8cffff28362513907;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91347729a221de44af60fdf2253eddb31a910e4c796f49a26a2e1c56509dc289f64936b43acfbeba8de2a3a7a6af82650906608cf89fac87cb08784df;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fc4fa9cd6efb9ddc021e66901d88b8e38caa1e04d3f0884a90944d0f1a4c6600b7398cc29f2f47e640e059c5e73534b44173d38dd320d39a952e034d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fd3e487c6cde54d75a35512657f9572fea35d590d26ae95838f5f38d3cb8863a22ef184ebf356363542603527b802d6fecf7f9adccc35007ad16a68b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he50dd3e8cd70c65c52dd7d79879307ac73104494df0f6f7c86c5a96db5c59ebf3a393a75f80a4e1ed57687a45e1432983cf1d153730c71fa5a4e4cef2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70e979f1ed760477ec78a5b742789e7da1f64ddea9da7b0fbc885d7bac57ec9843e8a102832ae80ffd456ae94a8b51330777789251684393537225009;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c5afe12b01926f37579559dc8c52b8e6b3e7f747ec13f0c8832835ea29cbcefe9a58977f83d5a0ac3faddf4a8383c8b754d9e7d9fb533af4dd493623;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6d5e3fc53280216e54b9279454eec166ed23ae5051126698be87dd306437cd1277ec5c3b6715f0a9b3af9adb6ae5de62d6ab0405e4c00c77fbbb4d8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he877cd8fc7c1e22fff902220f483896ae46e97601eb3559b7c7f9b988ff78e503c96a4de9c9152a2d0e8c02e0a3e17951cafa08d461ff372172d27abd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h571c5bc2b5b24a731d0763b2d353d8cf401dd3d26d20230ba73670b04240349329b5dafc33bdc9f784b122f5247666ef4666177fdb38894ad0aaeee59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c50c1701be4ed8a5ceabaa75ce31a3501b70072930e1dcaa071aa233b3fb471c0294220c63993dd12f30b416de27e81f2740b5c7c06e7f4295b68387;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6993c5b7f83e31badc6142da074070dab370e03fac1f3a9abcb0886eee65a9dc784e9a78065bcf99f1f5ab57fc64a333d0bf9e4192913873c21e4f9f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5fb71110695c90df8c251a50c6afdc43bf91c9b68c66d82dce3f2abf8ed915b9ca5bf21a0b9034d8822f5f5d54efe08959aac57aebf12acabcd1e8ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5461c405ae3f11f02c40ac2b3d80ce5f710cf34632bf71d957a9f5266260070ad2138924c447e9b72e1f28e46d2024d00414ce978c3800143d485325;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aede4d0b9baa78f1f438fb6c98593289ace09927c496d965c0f2244419fe3a211df18450af9d4a7e49dde7d016576ae1d605d3ce2600ba9f3ac09fd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h945b6ab834a72fa0c5fead197f4fde7688ab8850690f7847eb6b27a7358df8e00275c3687919301aaaaeb2986fd8c2c0bcd59b714a2c8356d5d7a2f12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc22b4eb4f1cafc260491f38d72c9d4a2dfe48429dca48bfbc7d36e745cb3d6ad71678c4050f71caa5555302439f4b7cc0d8f4e0db3dcc034a7b0354d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h436147aa2722186dbd46228b94a8f0d623671ae8cfab2553a328b2995ffba3cf8b4988f68f19aff865bdf182befe41ef40fbdf1a03442db82fc571f64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11756fcd91f2663b4e4ac17761cafaccba5d64b55bc3f6d29e23aa1f1ba86272811b1095f9ee89087e64ddff2b1643d0696a2aa6e59b9abf609fcf388;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb3507b5c1d660accfcfd42bbd1f95a5a625639bda17347bfdfc0bff0dd5e7f588471f07d5e6f8a4b686665f01950b52ee7cb5c914186b2caded35592;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b1df3df3f403c101351c75e41ead8445f4544e6795b75f1cfec46bf53287e6e40c586c17d8a6bba1f551bbb1f0f823483db5e4586df645d95f7e671a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c5899ad8849fe8956bdd3e65fb57a81a963471127aeae2a8b9c977928aa1a8542e75c547dee8d9a84b934c366e3ece44035cb8861c1a165d8cd95d43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0859110139149c1974b9bf84c6d036681fb7db4f7c7210cef831faf028610791bd90bbf37912101cbaab2bd7ac9d634e0a1f6244eb60cff16160a206;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb0c2c82e5e890970cb7cc8bbc9470a246ba0051185eace0c6a23cf860c275f3aa592b6a003e8c6cf080d15636335da9d2f7c49dfc78600bdec770df1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf508dca61c0083c86ae91876c1f7c1ffd2792cfe156721ea9454b8d681ac0398eb1efea47a82fde0eed0b0cd64242d953f08bdba5675a9ce8578db71d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f2004376786acd7dd4d45eacd51ab624d471ffb0623f8439ac26a73f366cf5a4c26686be8e9e0edc0b7bcce06415a728aeca75ffc4beea549e20d7fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h133f539bd72ba0d02f171bf55b8a2b835525d04caeeb46c1d41228a967bcb78fbc09a1313b802a374e6b3e317823f964768e0ba8e7bdce3e8778b1ed7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23247a24f86deda0a82e04b1d6d4a751b0b6e39d7392260fd9a04a9067ae3ef7f8c5bd57b8932f3de4a756bae9e3fa477a7857e442e2f58a744ebe78d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2b351def3512d0e2c073bb28df49f928b1dd84f8b26bf84df6dcb8afd91c1cb723bc7ae71c1b26fc07f0bd489e8349637ae92e2e4e41b72718614940;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc83b326d9c75653e00f62490435a63358215ac812fb7610f33f3c575888b01a79a016915abf5f017533742d9273071d071461c8d3bae8228ffe77994b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a874646f295ba6e94de5ac02830df37fd9c158bc7ade857b846a5bee6c070743ed522dd917ef6857c3ccd5c410179a609bbfdcbdb67509e7a5b58a35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89610ca8fb2a099cdbf69e48997d7a04a5ca2c5427169e9de6e1fd90b917d95055d523bcbce0d541fbf5c90207f0ed6e23dd1d915ffc05bbf832124e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cd52602010fb2d0e28d98227e3948d7facf52860f2a72de1d45b2a041adaecde3f5cd701efaa290a3da046cb780cfff70452e5d298026bc30b8b6abe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf70d669f8a3b733ee47a0fe8c41fd115b03171f4ea050e915948819e798eb2795ac7a1184d2e7a4072edcbf2b26f2893c263e464ec375d1769bb1fa11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c014920d7a3d7ff8a2c61f30cdea6d15ce6e1863d55011fcddfad7cc795fcdfc5a879ae1383bf2b5781bb082143cc09dce3aada7cb797fec07d18151;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f8979f8d67ac22331400b50742145eb28d225be905a5064bb28576fd143d8a5b31dbb4fa071c1b55b397e63755420a7a3542378160cd68f3332686e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb84f37015252b8729279fee5a62266abbb91ec6ba8d2ee7d7d48688cf5fb5d8875c0a1b0dda445761b119c747107bcd4035a47e9268694864a148abe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29fcd420f661ca6991842c6fc15cca6b5a883581caa40e85e708974d0dc51b626d96587b50ddf5f0365c99e77716dbc0615e35dc582aec9901c41e56e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h661c3d36fc383dc8b5bec004881e0c36522adbc3b1d18a13829676474bf416742aed28ffcc4ffa65925dcdddcac41f3baeb188c1c02353341ca010c9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69c944d1c2fc2c114a768b2426f43255cce6a2c5cd30e9342689732b003ec58cf7099b260926c5d53bfa9538ed496a312b72754711367b959e2543220;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf18ff450a9ecab403678c4db7a167ddd5f604cd935355f415725807a3baef07cbe5ab6f9433b9cb0aaa80067a9cac7a05604b881317e0ab6be4ee614f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc44a3646ead288fbc298d70b9f0db908d3246a8d10afeef20da56aca344dff560c47112c68086a35901ce493ac2a31625f40f9610d9f65e1eed5a6f9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd87bc44ce6d325e6ba02cf51ec1cc4841eaf8181a163751580cd2b1352a75f1308734af2a9cc4f7b9928462bf0528401bace24423f296a8ceacfff084;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7eaf44f60176929b6995546aacf5285b1e288d7ee8f199504252c617399a27ce61e6233062b5a3147cd89ea1c376a742b73e8f3b1bcc079b9cb4d78c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc55dec463d39697dc613a9f582c44bc747a526feced3eba9db90fa0820fdbacf7c38029305bbcf5e4535f2908a0c1cc310e24da00ad0b84a9646d2df3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf12188475287d4b2ef5d0538f0463a2915a7054b9707a849af434bdda8b487f041431ebd945f5287ce78235397d46e2f593e01cf6606d0723dec5203;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cf76833494d47dee8dbfd93ff4fc7f8e771c23bb61c37ae96baf2badea56e4091853183aa595d034cea5c6004656053d584abb7bd93af3133a8ca369;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc43ddb82dd9ee206fd16c8476270a9be06436cb3b5e8e7694cc630c1dedcd33fa1a43bae80cc8e2dc38045367215796cfe71607c2b41f7f2db9289357;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he68c4fc8897b19b7c3f2ba5116a44c333385d7f08e1d93086e1ea5a153273c0a379e3f04418a440e11538cac311c8bf69436111d2b18714382a296e3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b687ce02ec29dd311c22fae4cb02d97ac2b2cdca82d51a70a54e49f02daddcf02e65a982c8c5ebf13d6f0d45ee1085d1972e9081ca252dd4d42be7c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a1952ae1b91eca2411d365ff0b03d4fbae3cc819601786195c14e94fdc816ddb7ff1331229a5148d2cd9bcd6339035020e829323f88636bc81364abd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he74a3eb54e9306a6eccf5f787299d235e4c510b13b08dca3b77512069152b1007417203e2d66a634e85c777c9d14f9ee26e6a6ffa1012a9f137abe7e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h352624f1a9e2bd46c8b2d8567d55f1d47d9e4c5dd6741a7adae95b6168920987f506d38a10df8b7951d76a42556298306bba0693d1841f55aac2a4097;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea6388c40cdc08615886867e6944f75da2784decaea763191c96b85ec4da95ceb72382ef1592855f9312ba1f451b614d0d2ae5ba0549f9dc8e366a33e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6f514c2c447e3826223d9cad27e27c9e7fe79b33effa5465e1205adb81b4c0cb82136d48f80480e7e886fcfb816d8faaf3b8b87d0ccb04c80ab0ca2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h330ab80b59c11d7a23125435453a684ae488e124bdc53f86179dacbf77b15dd0801f3b645db6bcb0bc98e3118d385c473b2beea31eecb2789c463e9d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf40efe32866eb10b98f055184c9204036c5fcdc6980e9cb130eda442726a9253776d64cbbd9878bbc853819704cde0f44a22bc02364dd05c20bebff5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2431e22c3cbde4c9550f6b04fec986e4f360683e1d6b04cefc69f8f537a9b52908b5d9a168ac3ca98f54c1ec60299b684a00f0c0946c8d219399e8cb0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98664bac49677cad7dd65231b9de25107057c600a4d47912125586438b48dc42417f0447ee066ba914982b85b93eedc84e4fa9985d2d8da0e1edd1498;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb48a584e74dbfa8f5e3a2097ddf2e391395d0e066b5e3578105b05e0b336721b4d89d8d3a9ef5c47eccfdaa619f0b7e34081d91bb57d58e14bd3d5a67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27151f698677cd56d0d2d1cef9501cfebd12f6c40a785e35123c935437f2aa922bc741737b319a9eea1897be2c755cbf0a5505ec08fc49c4900c87a82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h517b18936d732a12603fe493a6ecdea4381976b84cca7e86efb40da3e5b09e099e2184893c9082d0034f129dc4f70ca2259dc558df6cde7258a4b23a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he28118d046e0a61a57a49ec4bac1a5c84530c48eb26a360b45816be0f4f45815554c8da82265a6372639f3e7104187c357ff9b3b0f1e0eed3b2e9775;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb2dd78674c247e923143acc53cdfb75f3af4f9ddb190ea533c838a66608f28fe739a0b4b1f97f43e1f96a8679394a97482447612bae7fbd142c294b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc04099c55477f58a236989cd9db0fb0d08742b3a3f02bf8a0ab26bce6bcae47fb550d148cb5b6aa27d2c708bce1c810182ed0592490b21f8edcc0096a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e83bf2b5fb510550f7ac02fd6ae7dc8cef0c2bf5246e1d6092349470af5656c60830414ac690f6f133c05211a80cecdd59772af9aa4527b2248b2367;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16b833f5c4e4a01f82aad0d2e72fb6e13c56333f48f362893727c56fa4c66298d62cf55aa8bcf8d4a20828438a771ea74ab3aa6309ab4360c2eba83d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10a11a431cfffc349b4068cbbf33f12fe6602757cf97be1d8b4e046e9afc09925eec7e643979a7466a4f8bba867f3ceae34a66999654b9b36bc1740e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd602fbcd17c79cee8146e4c0eb5b2ba1208741603a66397ca622dcbcf26021ffd3757ada9368e6e18edbc94fa7c0e17f325c2e04825eb6904cd79b200;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fc3f77498c3ecb0f71aa12c1db81222a3a235098f1c21c36c8853152a813dd24af53c95d3f0daf0e8f2de2d6fb3b8ba8409c0f04d14566a2c7c1c8c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32c8c8ebf9331da963394b1ec0db29c2d0a5941ce3b8bc7d32e8484a8001abb1520fee70390bfa6bd9e365748fd2d7253467d074a7fad0533ccf07bfd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf3ffd262b36638b3b7e8223e5de19fd350d3820a8a0877afb2deccbdd268474bf2ea4fb4f47f46bd449fab2e1e3627ce3bd6cba94b3e49f2a675658d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27f3fcddac7e7b8ae5c5b984ccc39bd61d1c706b37dd68c02a04f0335a4f2346849e25ccf06e754cf46302f15fd3d7ac78f783b1ead01a4a8b1b64fe1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85959c55938683edc809039b3a5283691fddd4cb39ff2a71480c7e598bb992913e0fe566ab25add57027a93a6d7639f80e9164e40044c97711065bab8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe4df62d4918e93b91867c4dee6be69cc577315d8d4c0b3643678b8e69f4fcf3171cc2342f483ad424a2f894856d109fd6a67a4ab16eafa912a4b7605;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba46d506b3636901a9e5ba256c6799b1ada17158916b02a8109874c86d215c40b94e839309b88cf46a816cf6021b8814777ae6d751ab72b896d1b4973;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha72c86b61d39da11bc44d47a93cebaac7bf9965551c04f00472bfca59690e7b151416e154cff4ff3be9a9aa52fc0696b2ad4051573d5ddaaa93184491;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdafedd4c4e147a541a4b4fa97cbce9b175a50d55ff106be841f44aebc6b0de839b3454c9b6d0c56b4e4c7ddf3ffd6b128076aab280369bc6b9e38a00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe548ddaa02ef87aa556fdfe6c27b3646682541040bbffd2423bbba147c5d778608ac945578a6cfe0339add4f6c0e4b9a24963e05cccbb9a871eb3d25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacd65ccba9dd9132d8ff553f77f0cbc8f4e3cf4fb097b38e258020bda2243ab7c2b3f4c4a7309206f93df3133590bbe8c693320d75c2d4ae8a18bba6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77b0e8a27bf97c249ec091cae2c7ccef53654ce542223902404686b49b4da2d2db1810b16e77a0f4d2f53309ba37ca13fd19aad12d7f2192188b3cc86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1348227fe017ce2d1512a0a830f3cbc98dc910946c44a476f8c9e20ba49f849b40711d1e2308724771142204fbb6a16e9200483c39e15f9c289c367e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4d10b09ef3c54b96b008f28c1db15ed85dd0b87866d5f87fc51fcb7cb2b6f9abb9fc08cc55011f645eaf01f5d3c26397bca8ee69bafa35d5abd18c7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9db10a95fc34e0a787d6a8f8aa38bb0f6dee3bdc8ba3cf4dde01355bdc1ee970cebeeb315ea08a7a82a5f2ac0519b275bb749f3043d8a034e4fef8617;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h867f2d39666089f9c31396091e4da9a5c0a86845a478288c0ac8144b1da39590b4b168049047b459f92bccc207c706331ee1bfd0cafa02e968e5bf17c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8652caccfc691fa24bfe4ef4e4c402a665c7e1ac1a41ab99bdfa011d6831e110c825b81deb9842b18900e2244220acb85139b815f24504abba5cbcc1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5624a036746ca4f3ae270efa81e3edece81df14113109a225a230d430a2cb249d97d3ae57d0a29ba7d7922a8544ef042b25ca987bf91acdf336d680e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d7c9650380a413e58d4e7664e24d8f5a858147ea45f8c6fabe837fd81391bc4ca46d0da692cb8754a1decab0f095116e7987f7ae620e793ea59c7285;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3324a2fa0fb20979130c87f078465822f1b473a54ace1ff75ec6639c209a45e50db1ab5f93f40fd28d9a65258412e0a06d59c9f478bb846bf8dbbdb97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fd12fe9e2d84e0b8c30942de0e0d16c03d96b6588129da8d97936ee7a607fd2f5fbbb507cfd356d317d82bd8f289a8b97338ef102115cc02fe708af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2576b59b432b63cb6ce3a0ec749c19fa3ff538e741b7d6b20f099d52e41dc2a9be5f124fa16f09f290051347f7fcf791c61c4bee6d2472bc7a2bdfbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40315b6d7fa8b46dcc5d02cdaae43e582a95c41b5eaf5a085a69a2213c75fb44c340486ddd97245c443c01cc4e41a51aeecb3c1c580d1610963dd2f4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9acc3a753dbcc515e81df08edacb2a26115da928a6516030a50110f28d59c1ef36a53a7a2f532525080f10b7b8c6b716e657d465a17eb26b9ca920b4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2397b311176c4f609137b4687f93e45c2f7cd66392270892fe607a8472e455a26b5d185cbd63e85bdad3b93e8d861e516eb85d36e63acc7b4ec089420;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f43c7ee5f7886883f3e6b9e2d2e37a63ea4cca084f797af24129696bf43f9e0ca0e235076e920f6a00d0e466d69293b94bc718221891a819521f77f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2ed15106f3a9bad8d4bb3ce85f36f555c129a9e965e7ed427380c1d0d579bc632d412a95a3b1cfa602c17cdfb8a9ab735a8e109e6de7c80a9b8d72b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc84b1c17448fc37a15a362b7ddfb2d4476bde2800f71d7addc3e0390cbd5e13d78602f920a0888474121a7d1f1988114f159755ef4d75fbed67fc2916;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc6ba33477a380c6bc692e9347f64e3f909249c64f1dbb4cc14866c3f1cfc138ce704f58b53e656a8b812b9b427f5616be82cef1786b4f69451886611;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h152cb7681a7cda6a61edc40c9482bf30ecabd0225bf1d434e57b4753e4877f3610d24b82d2c3ce8d43c6310c5129a682f4c72643d39c374cadf40848b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde712981e13bd306767610f7d664d6cbf178a4ac164c4671fbc4710cee906287f5cd01c3f090dd35edc4b8beb369cd97938cd47e40f2e91178a197e3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h444c4c11023c044e44994e603fa675a8a375c36e907cfbb07a7dd0d93634f7a299406fe2b438b1ae9a629df45552a4d3e7557ffbdec6e398cb8598f11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h595a153a72ce7fbde1fbad6b0256d175e41fd9fbf4bc4a973dc5682b8be9d41fa81e878a6618b5489ea7be9c06d5c66d21c16cf3d6d58e7f2b4f0cea7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7c6de3a403201579ee5aede362efca562c101ce3ba42f7a90ffe3373796adc3484b18ea8976a62267590d16741ec2698cd1254ec3b65807a44c8fe6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4693514ec83fa7105f7e9ecdcb0de0bbfe3c687607c13e2ec7ec1f6a978beb5ce8340b80daefe16c9947ff7d626e90f0b207fc31e721cada864c11f8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9226c1a325b374cf926e74bac2a08d043db9689b73899927fb250afe503bf17df5922b4bcedcffc5ad61956fe8f9616a9651e30718eb0c9c64c8a4f56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6d39ba855b64867337c1072840439dd179d9efc1c283a393ef592bd7863600a70b60854299d85f4f9a3be99e3efe581f706c0543b60eaa5100e53b0d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bab91003ed8663fab8c1363a1f5516ff5ed5dba795995250a500b69c454a73facd4054192c59456798cb7cd2701e7d73bd4cd9e662448c59f88c4100;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb77ddda96db6a587ca6a08f5152578ea6b13c0caf6a81323f2bdd5356feb02f0af601980b750131d002a0ecea9803486e55dcc5419a6bba6b8d992cb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7814c501842335c8ed23813e723cbc30db396079408995685d90fd56caecc96cdcccec047216e7602e8dcdc634430d61b17da7232f160727b4e60155c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7899ebce86d363311ecd3bf67f996b4e4b4f82b373eda035cce4928270ea37249f54ced6a8798633c88a59b28823854f856c882c685ef5157e06d601f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h128aabee04856dd5ec82b1412e8ccb01af2f4085d1b07fdb46eeffff59a3893fc6c621741a8988a50a583c580a1ba69531d6a4521c4bad1b902a4239;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha31db2c74dd5fdc5603a332996b6706a3e33e132b6a01d30592e1cf1360163d1d40fd6a192c69d4f012bc16a55f7d43dacbd4d55568f0b7b4ce318d93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c72097896cb50eb68e80c7dc70f46ec4863739b245f54715960abbb6286b69b9d274883476ef40b31dba165e9dc1b181178b8d3480fa11c595114ed5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce87b72186420cc2eb6a44aadc3c7e76536c21908c8e933252cf578d857c0eb560593b3c02d235e11003381ac6c86969331e228264a0e88ea399cf772;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cd7b8a73610e1da3bd12aa543c86a7ff2d35400852dfc76703548d49cf519a5ca93207424760972ab5dfd36e19c74d3420a6263030a6a419862acccf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9e6372199fc242b96624308d2c23e713d58e1599b6f4c0d81dd3b24efcca995699d1be0ecbb687ca355290ab8552735ddd127e5f4095d4008c24561e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91413479f663dfc911a080e37dbe21386649608273f1da6bf138c518522bfb868db2f2c0dd6dfe4e12a5284bc0608acd6a32e98ba3afee1e5941861c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d532924627bfd2827aa19807c3e9ff6322c9dd6963adb9ca0c8e80d6ff077990d4b801bd788f196955b5caa4373e04598f7061243695ea9d5927034c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29f769dcbe1b0f78d22aeeceee5c8edd64d8fa20a6bb85a94707a6c1f88ea0bf887c9686b851553af53592aa95e65244ab9c9b31b4291ca277c491a58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he888687edad1c02fb71ae8595615ffe7b20f78d4056abda76307bbfb20cecadf38c0d4dfc8754c5d7684f899d7aaaf325be85a32a7b261e199cd9bf64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e3f765d5bc8b60a82e956fa123878b9699dd4048e0ea2c46316082a69fba0d7a30b1a07a8f1ccb15588828aa03d5767d191f5720749e35fb334dd6d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5618cf968f2dadbec53f45504f19a659b0b9ed45b9e7f66774fb8fbce24a4fda3ecffc42fa50ba766c41225c17d641a8bdce2add233589a83e122f1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f470b9c9a8477cb44de12cf42c57625b36a5bc90234cacbb157f2594ecfb15b5ceb4373e6a8ca82c5ad4c13f8fc225af97b3f429d2693192722a9ddd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4959d1d2fac3122b455d9146e261867d0dfd2493af822fbf8abd6f93223ccc90fb443fa7b7278bead5c8fc321c7c34a3ae61d870a9993363fb8a30b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55964ca501416e09351aac725d003be6c6e97d2674f404f9648a477834e6c42301fdbf6a0c263341a7fa47b09892202804dcbfb347e7bbb6f52bc7b49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4309cbc6a7e58d3da84cf7b8913990841dd76d346a3166b9ed4d893fd732ec3d4aa51646612d290b591b108fb4779fbcd62528a6d0722a7b8dc2003fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44708bed076bdfec1ea6254a07a7f2435329c52c1b12703d10f84ce9168c1144db888519d676f79eeec953349ed94c6ca8648285833e11824c46cd0e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f3bcbddf591fd0651b0134d87e5920bf4d99a8f2a111a432f5cd2f6a06d0a8d485a7d5b23d25c0265c9b59c7b189f409f96d77bedabf8540b15e4fb4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60dfe31b6b71faea134ccc846a1047766f54baae9a449dc90814a8e7bff310984b2361a3345171e4b0b7748ca9fe294464881989911c4c77ef8dd2560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h266cd3d92bc26b0bd9ecad5734729bed6a06028e7d0ca49f40ed53ef13b4c993a09bb4818ed297bbdf4c3456f19f48db378438bb273398d305138efcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99ee13316814b89ab10a0629bc4c587622b0218d61707d81dd7ff49fe444d33d22de44cf9b61a566760776a313ecd2ff82e5da1d4f6f3d0463c3892bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7de8cda2b21c29c79c91e6c02c1bbe41f7236929d6fa6caa1d09c25aa5ace5c6396dcadcc77a6b913c863ab88613f15c86bc1a077fb6d58bbced9b189;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha657894dafbae1c61753289d4c5d13fcd2c5e72e7a74691790029c9f08a4031d8c9f2754d8aaca3a44b0c626942c75d96134c6a6d1091ca2fe020c23f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6bf7621761c80af6bb827d84c900ddb28edbc9662414cb9acd600ae80d8d5c0d92f0da8aab9be323e90a5de445d2ca43c95cc3feef46234cceb3f87d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f4d214d0f5695aa5d3417837535494293acd966157c5ea853b269fef99918bf2537f470542c217a32f3329f6abbe6dbf2f5138816953546aa5518ab3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3aa22eaa2d4e81beae067136f6416f903330e79aa68a6f8b9fe752f487e1f0637de61d688c6ab8584def50ccd2be72f6de0dd652b1084fb1a40e4a375;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc860f358838c3230785961767053834b2809ff3332ec3713209b5b4885a5acc9e58a21698130cf3dac08d443bb11bdb7f7ea1d2ba6e0f969c6fd13701;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89fd3054187e0f547fd1f832ae4a465664347f47f372f6c58b58fe8f28d9c273282f55d8b0eaa80148ef031991a259bdfaaf6aefde12335bd8b0ac31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9230c166083e4612ae8222cdec78fe98bdf3a38d45055c5a90a5903a4eaac6c4896daa9b900574e71bf00bb20a762b54da48e6254b5e7d9fe8c423fe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h884918e8e7e7f0188e77096b9538e747812be23055972c4dba8040021014f7b49b9b5759c19aa6a944f35ab87fd48212866659eb236ab705e5c088118;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1ddf8601a4762338d11aadc2dc6c5ec535d703640e3f9e542d06d17ebd7d29771124432290050026293c9f6f8259ca3e62b0915c2e94ab038025822;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0ccf9b6b02f960de6762cba736f0367036d0fbb2a32ab65ebbcaf3edece1b5e02cd9e1753a86194d18d5e832beeeda3dade6f615523b150b9d75296a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e2737b4c681437daf96ea1633679f1544cbae3226b40a4e4b1d48d2febed0b832e9eb49778db64c8444e1af38c5ead9ad50faa6cfe8a5bce35da8cd9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59852ea8b6868ab61c5b6c6389d603a1c2715d3791840605c4714930a5bca44e8c00094f043cb0d8522ea1005af0808b37d899e3058716a6bc0660ab1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cade51591862539ea0f84c3227fe449d973b78c5c907edda73ac628c15373439977e6e7acb371cacf1cda899787c1452829c294b9ac755f83d37ca47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51c36ef45301fbaeac5325376c406be894372fa4cf56945f47099a4650bcf847d7227a4c3634d140497df11bfc1174ac18605d39890130be9def9bb58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a8f6e7f6ed99fb3f32901929834727dcfd74d1992d972d02a84a11bc9b8e1c99b6aedbd3d88be5fbd1262ecba635fddcc3b55ce2c5f0e34af8025cf0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5febf04fe8ad2070fc77232804cb594b718dbf361b064935750de71c0f321f806cee876aec14f82b79a4a0c453b278a7bf4378a841ab5d54b0c58cce7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe19ec5910b53eb5a2cf21dc580029230a80d15d2947937ce133088df15703e0a3508a19d012e5dde762fa9e5783c3dbc593305c304241718778635c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c03f705f8ddcb21ca2440acc58939f8638834f3286f81642f03f3b6c781623382211243d03d78eecd36bc48daf7bbfe575d5a2c3d431f314b1a641c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h482de8f6607490e17d5f02b0668a6b348d7ee11ba587fa4b74ca3b97b0e4985bd972f3d98206ce181a4e6a81f4190833aefff6ae80cbd04188a3b9fab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95756cba1adb773b2234d19c4b14085106c3aac338bf9e79bf8d2bc3e1022495b979791114dbf94b4317628ad9f4c163e42a7596c0733fbbeccb7093f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3cca271f059edcae3a8043b600369a22e10ccf05f5b99c3d6dbcd7a8bd1385794790892f3cec8ea5b43370dd3ce1fe92cb1d775c7e6252f3d9bf6ad6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58e544cdcfa21609d5822623d0607589f87a83c00dec5b14490cb56dba5e6d69a66e128211c2092f62a0d94f7854affcc6077be00afc0adbd1f444926;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33ae094ccf5e52ab765365504adc00f5aae571b20894333ea32fbb88b06928a3b82f429be8a7faa15630c1445d870db5291a80213bf37432a39547162;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a1f8616038d6d8ff81c7765599393718ac8f26108b39af2c80c268b7cebc2af401271ffaef82252f9105d7789f425f6945a823db7095d8ec44f19dad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7e0b3065de6fb820696e39061f363abe9687294602a0328ebf79a475eb476e03f04c3d718fe603dcc821af51fcea6bb211d50b86b55391f6d2e66814;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedfc5ae29b29043e788f3f73a597e9da86ca844a55882ff9163175ba849007dc976037812a174ad0a043327c4835158aaf1deaf8875be0df9ae6800e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h611ece38624edac6a6993a7e76618d4dcc451b3894b4e0eea95f512399677bafaf2dd5162332c77bb3c75ee194511c22ec58e6cb41f77c31ab5e05a2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11327271ce43021b10c16d360e833af93534bf44f4c7c0234db058aa8cbc76eb9b7ff252f4b90a9c41b1be497c99dba9db919ca1a6a0132cc7019ec5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63d1f15e1809527194aafa4ff2cca1d597f60bf2a4b0eab973888a04e820087054cfe0a3df281981a08409af84e790d9d02147223b5069f9aa8a7849e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25583ba6d4538a4c40407f6097edde93e0f4c73739fac52983ffbcc5c2a3384f12eadab2a796d2b7e1c31bdedda7fd812995a506549602de02762bdaf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6825201133d094a0635e9cbdb6530b78471917b0ebe70fe6a1440659b3a90fb6eb65c9094baa4708ad3945f5cb64f53f7e560b645144e460e3046eea2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ff99fc807d2b87da1210722b3b275b5023c24c8491d06d8fc52fdaa665e2cc8478d112ff5bcd29d8782ef76b368a7b9f3f392677a9a8f0bab517e895;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h585e5e9bff3b98164cc26c3194434a73bb8d65d2330e4895ad1a654d2f1174dfdbfd499bad1b32273489a3d2ff7163e05f6947a1c100141f8ad97cf51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61739560eadf09fc49a313b903b947227e745447066f3e74218a102e2f83c7e15f7873a7f4e6d2970d8a64f420f815977c45f2a5a275407caac82f5b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8767a45318b16ff778591eedd0eed824d08778e07e2a08647ed96966cf918bea3349b29dfcbd071e7bd39ab84cf5907c35fb56ffc72e2be10d60e420;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h846645d20e173f997760481a70a12050eabb173b04921628eb10526d0284781727a36cd0191a9dc768b7dfcd583f65b795bbeefb33df418e5e56159bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a70711eebfdf90b9778633d37e3ed70d9b87018a911357bd162e5937c71b1cd67ba8d9b938b1a9f3f9efdb864efdb7069f279890b6b79aa9eb94061f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf79bccca2f5a3c6f85d8828a2ebcd999c39c77bd43985d8363d47869b5090dbb5e316c1e5f4c2d86e36d2b376758433d018b1c840f9942658f1662ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2611fd47cf4002aaf70a4b276e5c300fea500cee251f9c21d48df60386e41c14cdf6a8c9f952ad389d78663815e4ed9f402a7406a919728b4e21952a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2806e5dc5330c4f8b43c6809dd73aa3b1e6f478a3262727676eb997b014d15d08f7b0cfba17b97e4d2ce2b7939e02b4f39188e0f1daa3055a0596401b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc44934969c60e95777d2795a6bac2200091dfe01275b5027e5aec1b847d9a9f034d6a934fe6e2d72543349ff8ccc95dfb565b3045129b69fdd09cb9ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h450693c227fd2747c83cbb725ee0c5fd0e9135bacb5b487408628fe414319867d13fef0ee04efd636e38bd14e72069621296d5ded7d59b3de490317b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2923e1061f123f974f8a38c18ae05f728a9674ed4aa72b7ca9676c34daefcd320bf601149754cad9ea49e6e429502a224e556387fd97aff7a8ebb1c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h981a10c9e71fb95e23f8786749aa106b3268485904b93a0528736713bdd4fe346ab2712f63f06afaa0b4976cd721ec5c6aea6b1f4d1d3093d119f61aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c812eedeedd52938e63de5d9f2a143b8ac89515b4b11528f515cc33ee11e1f4a1bfea7669419c61d3bcb6dcaba4c7d7af9c4735e0cbd7e332505a0de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bd23c6ee30fdfd9fa1932f211079c151931196596288b62aab5d6bf04291351cb09dd4e24717f01484e402ffc82486920aaa78d994cc7bcfaea22ed2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h164318d925b3635c50b5100e0ade2dd4cab9d7f34d1c5af73c14ca6c5bb369ed9b03f5c4caf790e3ce7e2f5f005a77b6ceba9144f4f39221a9272599e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45913f965b564f1bac3cb795ef164f8e9bb8948c885df7f3fd8a12e83e2f08ac0f10da91d75d41eff877f5f913d5d3d3f32917b2dfdcaf3fc8b4f4f8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb24cc9b12ed090068edd8b7155e3dd813e4e3930201720455fb28ff6fa47c2145835a2de762bf3778d191e774288ab29aedd79aba29dc505b1950a40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf75dbb456d86a0b3785c05168f08348d1c79264333ca48e283c08ede128bc9b65ceb8498842bd89f62aee03876168522e5e36a1cf062f9c994b7bba9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf38563c94c6447d6f4711599f8d250bd2c1f243671d03aae4bc2e53a0362d3209cef3bb09f8eba40d50188c965ce4fc2bb3e28175dad775df2a4888bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6c2474523572a4e18b60c19d31b4aa40630d6415e37d12c08914efe77f8747ba7897508d9326b9fd0bba2a142b845ea52a85f9a0eee66d05dc3dbb7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4905921c6b5aa5bba96fd13a802d4c91bbebe0643506e43124b30e661507c108b920e53e74e656db0ece1c391bc9cc2cd17a0f9537f8e24fa39710562;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba7ff38bf9c6062d2edf0c57dab80dd47d9d159150eae3c73d568937242fceb2347061567b6492d816a746261991ab8a5e23bf9c0a5f64e472175e6bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde217de16c16fd138cd903361260335bbdf79194f53b190f372e5b55865e7a99fcb4c6603401224fcb23741490b3959ce9cc659116671672bf44ad68a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e139006898342b286698393a6c49f4e5d72443fb8f6e2e28e2be0189ec092f831704bc52f5af89c07d5f5fbfc7ad775992788b33ca2ee16cb94463e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4c15f47b29682291e3e1763cf37a6ed80ad7bf19bbc7aa48f34e0f9f7edf65bf835f1af8f6e1fe2a3464b3d1520e19c4a7197ecb9a6b8091134073f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h544f8e62109a0d3e3823f7b89bfdd91bfce8228eb2beab5bc91ba4cf9740bb4348fba383b5c060dd7c74190ee2c979947b1dfbf5e23dacc677fdcb43a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39bc9c4d39e89bc5bc59250b9b6f39f5156b602c4dba3a02d553f88d1e72a56bb7c1a39f7a62c1d9d3b33691d128d4b2dbc96a9fe2cffb605816442c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h430f9c6153c52b564d7f5cdd47a70be1b633b7c51a3f87e1c9d676e375c6a866380bf429cbdc6df2a30e532d52a919b256f129ad7a5522f94ad2c17a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2701d2c54586d3ec5d9d381619df5622700e471ad361cb406424dccc3fd7822b1544627f319c78a359f9a83771c76eae5d275473993ef4dd848df520;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba09c7126d19aca04c482a180771547659a684e33b23268ecde59c5176c154901f260f3d670cefaa7557f4b0f5e1928a2409f5e4e1c28dbc18ba503e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4baaeba79963e9538b42fd8b0713031d2b9103d1424f4edab04fa9b31bb9b55e4c746cbcff36b2e513c4051ffaef196b185e8e2322f6f7c127d526aae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdba574dd93ced2a8b461b15b222f17092a20a812aaee90c286300a704a5bd7dcb22cec269254a00173cb523e0ca06d87f3f82699380eade4792150aad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had020e0e08201fe98e8bc737c92baa2e757fd09b95f742a4f99bbc780a961118fc60c2d311ed14e4167110b5ce42742130d75576996507bdd36002759;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c1042b19d2352732ab44d4b98ec57c33bb3271272560df4a1079b5b0bb6985e5686a8982b8690c953bd11fdda5914d88d2627fb639cfe9c078fbd5dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8d49095d84d1c7714a49125a0780144317c5e85ebd7dede188339fa355ff17d6957b61fb41d08f0708fb1065eab1620b08d5de2bdaa569b0365291f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58cb633cd0bfc3c8d0f03ed44ca99552aa2b39714c6fdd270bf999a11f26311804a182488f0fe7ce92cad4def21c21c4ace8cdb71cad17f5a7f4b99c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3dc3f2492673895f32bb52904da38c713224923ae56291279d666dab2128d00cb2f51d69e464377d33f47c62ef0ce9a9c2dad394d72f690c3b995d3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ae6ba0dc6f230dd4914accaa47c3e57be294fb98179e1b0329b1827d56302bff1b1463c1dcf28f2e1743305b6acb926a45b00730f6f42fe77ea4d968;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf925a882cf744de49c8fd8f61b46b000ed495b4db35a606a2792a0eaf7964308d13db021cbaa7eda3178956ea02a0d3fd654951de08a85d2977fdbf26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c98eb4fbce2a469302b198e2c90192376b463187a9c2089ea77219c34bdb708897b30860f6d6ff73d4b36f4b1f1b772e744e6fed47121ce360ff79bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62e387264dd34c45351ddddf56219c9c25b0ed528a854f07f30c714adb6b9a2f2c797b5fdf42ba7975145756f9d92ff650a1924d511bb1e6505e1ba99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51157341952a9d4f8bbbc627c095aa307994e041c56789f0ae8a9b5cadbfd8b3489d1ed21df0816736fa7c626e3875ca1e52ed17bb6316852c25f9b46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb393c9ea372d1f6d02262d3f504505b6003e90c66ee5d0edd82f3f70f18e49a7bf247104b1ba30342a913430d02305fbb3ad16231f07e30c12b113507;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h669a7189e42ab59fa201331ea2bb201d07addebb1e4f462c5f8493500c02405db0cc13040f012b6645e7e186c5129664bab6c67873650804f9480baa9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ac1032dee3d4bb12799f6f51bd574743574b819a6fda496b35a3ef437248a943c8e730e10ce3d824d6e3f57798a3789db84c9a229cfcc490acb59bdd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h409354a1a265f3c8ece42397bac21225d4117bd1f9e287763d2c8f8576f0ea566f46601a376a3e2b575ee28b784ad08f9e199772a780d136dcca263f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he47f53de063bddf9db5feebafcbac15cd6e525a64bb6632aad023a76bb354380b5e1569738ae29f07f478b74257890fcce81a9e89898b7fefc007355f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d99a35f6434fd47fa33a8d76376ce774449f4551db288b527ede1c32754a14dfa41f89592a3544c2e88cd4bb8116fa149e5946c02ebf25e8b6a54caa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2230da113e7e7a3b59134e203b741c325969915487a03b6c55edb9bdbcbf14386250ae367516b341565f3b458525293906c94893e6c85af3f0940e0b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h641a2dfb0634a988c8807774d4e2b2fc15f8e16cb79c67b67f082770fb618776dcc930a35e4b5faf65306c63469401fbebdd9c1accb10ef952365500b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bc9eb3a46f55514e01bbc64eb50fe95e114eea20e7586d220a1d0959548f6d75c9403caf1fe32b8229c441227dcd04a6b5772d443764646eab14177a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h732543ed8c0ebf10146bde6e8c29dba58ae6ba4faecaa551bf16796d8b61c3bfbdca18b5852c01a5c9f285a88ab4868b49bffe7bdbb7d65e0d1fa19c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97b643bdb513c4db35365df0fc6a2bf9dc46c0235bc7ed7d01e64e79841233e9cb55b4326ec6c140de863e7bedb882c717bdfe6ed776d381cac8f11dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he764046ab7f09f94281e9f89cfbf9225ccb1f4bc1d6e93c0fb9e54ca2501a788ad1e56054225a3fecc3c9b5836f3d940c927b8b12d88fde3c1b1309a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8dd87f16dbd985536d14ceea92aa19c431221531236b0dac40a9f18af3a22a59355832d4c01e473e2c4fb0000b1c21e8300ecbc5038e4edd5c06e1989;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91b9c0b6f930704352d0470bca27e093111aec19db429f94c4f669d59fd1c53376f5aae935fe26d4f92d6ce8f2f26cff03c36699626160955bcc69a77;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcee7215d9a10483f9e854b7495e4d381812fa2bb299e32f50d365dd1bd9f394afb8693ae13679058b961c25a6580a98bbca2fc2f65c9e219584b18f44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87858d6567c3bcf6b33dc6d6de244548ca6408d18c7ae1aba2a7c70751d8159ead7469f1f4e5057d3359eba047eb753574733ef661d089287e25e5165;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f870332c1d5f76e3a410e353f4bf2ec6aaa21629166f325e83df31856c5e1f991a0b29995ac5d1a12c8ad5ffa30a40980833c22d75e2a4980091c105;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadfd2455aa56e4bd385d275b1f3bc55b10409d1f3ce60b9c6c2f317e504a5836eac9b0ff1369da4ce9b8ed262ab24b5bb2d57ebe352b1847ac1d49176;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd8ad11abdc7665a4e4c11113058ef1dca70c3620d4ab62f5ef0f07832907adf2244b62bdd5f7b3fb3c358c781be1fc10e9a82ae669da92255bde4d2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c9811a4dfec67bcd4ec974179714f66c590df4bb854f4c3de44d56d5bfd4eb1b8f53896874a96932261fbd3385ec8cc59dc07e4e8d1ed0c64a141ad7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86f5862e2fcefcaf1b90e5c17894c9ab6e58dc4509cd0679e50cda7898882c0329831d895287ed8c648fa1f9b83ed61368004bb7541927542fa693573;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h538bd912385721e2d68c2fb10f85ecf22e5611055d1920075b2b9c16ff550277547dfc0dee2b328d5e225cea88512f68a00951c736d8cb1293fb176f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h629fa4a9ab01031935cb3ecca0dd9968762ed2056819c8d8b0d2d6335c52f23c917f9bcb18b0436d1f30e750f7960b36ef9d30c02f5a1ba04553b6073;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef832b8a0c82f8cec3458faf2baa6dade64f44a04459b52f9b25514b4226b77898f912e06017517b45b68baa61af7c3337b4bd83eabdc04903cd525bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae737ea93701b937f056ff353176a42ab412a3ad83588bf0e46c9b599faea4090e88c9e42e254626500d694354b02328c97589703979cbe2062d2f21e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2122fad49c84cbe132741f5439349de352ab372b5e199a0c60947ff8d0ed348a2bf04021d1ed90238bdb3006bbdd9bd1b2ea62315542f5d8f2a709960;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b8189af81404b9feeef6e2310976457fefe17c410dd970ef62769db64db4d5469fa440d0142f966c5a0e051e9492f287ccde668fe4892d8bc83b025a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67f1d096a0a267b82bcd1a6611f5242c2862b8a417bd2338df3676cf73df24f3bc4313d82ebadf59e43272f4f3400528963b5a19ee8980b02c0d87867;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2219c0b463f0a32a8b28b96ae809c5ff316dc0cb003c52522bc79c7566ea7322f205963fcb078ff0706a7075ecd758f071de76f3ce234da9ae678314;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6586482ae435450be094dcca706d984fd6cd513bc189f3a1c47570616444a627cbd2effd62bd88afc7bb1e48d737b6cfd3a510190aa7b92210e16632;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcad99194098777b2ccb72bbfef05dc3bf8df336d4351998af221340222f7b70be0cd9270413fbf6031b5344e405d309db9fca8ee0afe364c2fe2094e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2aeea16076e0949854070c1b4e8f6fd50505a0b3096b9f9b958852c445e82d6a283f45fff9c895b8e117459b7e3d3f78f1339b62e333c7749fdb1980;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32f127bf81dc868972a269bd9d338ec02998750f47005f4ed07fb70eed6a82ffc51ae68dd0fb90a1264246a5ec34ef5a87a0f3a6e7f0f35b1239a3f23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6885aee601a59792b6b05dbe1da9a07975eea639d46047b2e59c0de139fcb65a94742ba29f1f0b17b416767f23141eea474c0e77d0cf220ed26aea016;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8830e54e8765fd9e8823611109007aafd0fceac1fc156183f258d108e687b222dd6b7135f376d1f27057cec06a38c803080c6661451ccb35b7dd4321;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h577f12ce3bf346dcc8399137013d02c102a5ec03e58a14959a71547eace214747be783385bd7bf7b9a58570295d591cef6490d6297d632b657474036b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c50fa14f9d74cdbf54ee92718806dd16fc68bd0213860211fa410cef74d48307b87990cac78b5cc53bbb8f62215408eb0778fded4481c3bc83704406;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87a0b678fb576d4ce166c10ceaebc93786f086bde64cf75aa2aa5767c5a66aa0774288b2772034fef8387b83119b50af6297855bf12d4dff95c0c45c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ff4cb9755e286e7d335db6f87e7ff620618a2d5921c16a6b74ccda1c4ade84e2a196ed0c12e2ccbbec9aca60d590acd086ae6013a4cdffb481950d6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha217ffe18d18cfc6b14b7d47e2950ee7a7afa031dbe29b5ba2c1dc6367f7b92a0c2eee5da3f214abc1961e1b88bf214082983f4412b7edd1a188f1cc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b029c53092663d64880bc735ed890378c713c263f53c392053aea608c4c872caf1b57f838af8d352511b750134fd1c53f1995f5b46bee48776e5e746;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55dfbdba7633274845fcfdf83c837071c3f733a07253075f63031c9e6f394c465601d5416c14ddea49a6599d1687f3847b92b2e748ad0dab6ff9bd236;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b6e5775c75a92f5ea51c022683a6e934b233ea25da98953b80e2caa8c6ee024f22c2262a21b51c6309fdd2cff0c4d3ad9cd5e9b0089d4ae1b632f61c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b8f1ad3051cf147d6d5f41e2a1897ebea33704bd3731e374f463ef8a784eeb41776c0c86351356b0cf707bba9818bc9f6d43c922a055b97361790bcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1736f11ccc902ac0064cbdd77781f02e3b479de85b49179963f8f1878f1150a03c711f182e6d12750e5e4d5e6fbb0b9fa19dcdd724f5257388edd981;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f863e5c96f446bad1a6a3303651b2dea09c09ce1ddb875feb0a13c291ab6ae0f9df5507fa2c6ff214c23021b40761fc66594f0360811c52ab5084bd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9818ff3d69b6a934570c5be224bc73f7da38ccdab3c208a2d071d7c7a3b683f7848f8cb731e14298a562e626ff97752f33c3396e398b1963f23c7a5d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd2afecd5dca06b6d69080e8f1a82a1d4026eab404f0961fe78e1f105437f5090a9084d0d50df2cc7df48b467f1a1062e179048106eaa96a3ece3f755;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h499c7e157c0d0f4a382b65e780bf5bbae42b3ae55e67d6ce3ed4261d7b8d3c433e15a2310689dec233b230059fb8c1ce6b53f3401d2801e6720b4258;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc13b498f349819c58d142a78978c632d8a9806dd0e9b488d409b29c78a670bf9d30d64f1b11582bb46c8e5154fa5a335029afaadf3a697cc2809d5418;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37e92d576f3912e68ac0160d730ce245b76fc6060500b0acc7c99221443bab9a3ce4ac3fada5230c60429346924151744f3d5fd1f252c0e153eae4068;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14b5be31cd8894bdb2dc00ec106921e68a24dcd05a1449fc3ebe1d50958308d722650ae094d00d63041c2d62ab7f97c854f0425588de79de69673619;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h325420d10b8a82a0050f0b8689ed367388011b20cb0e1d877e4b15efdd9146a23c729aa5eece11117def82e9554950bea1da15b724ed3adc10f487c91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7291ea0673d7990e251ea5a7ac1fb3d3b93b1fabc50b41a1fcbf97bced211a28db98c3bb05f2d2560a8381d0c6064b5e406adc816844e4fd5178f8fdb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha173f4bb1f66fd22c418de71a00bcb3b8dd410839bfb721d39baf4f71344d1360cc79db4ac5dd6c373568e5fa5d65b00e0cfbfc5c3bfe0c6467831b2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h878d48024c9b4e20dba12ae26ba536939bc39ced088b456b1c639e0a0425d1a9af780924b50bf50679dbe586c4e3ff9be24966d6a935e306f61e05a61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3184b16c8860e74df021fcab00c6312a04dde5a04cffbcadff19da907043372dda39006c65e9dfb5bbc10f975492d4eb036f749abec7effa943830da5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37c46db0f584326de6921d1b537d634d841e9c224f1b3166e7ae04f1b4c46e9fe22aebec38827516af5eff1c9ed224cf1d6fb73a8fb486741baec9c72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd206ab98e25a4ac483adb3c7b093f173dd950049c30a79398701d79453c995e0a6c866a12735b91fcd8773a3b73eff0e4ebb827c4bf778499d21805f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec14673830fbfd32516730ce73b3fa8600495deec6449ff2943faa95aa1a7c7e9ce693e2d9ec25d885814ad50bb5b41a1136cd48c263e01f451bc9de7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13dc92901b64429ca321f4ebfe6178f94a05411a4abd5030310b84a2da412d263fecfff2528ef36aa24a62c47e9e25704e7c9f5473adb869483b232a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h267564849338a2c90ea2fe3e45bb1bf77bf56febb626cb59754d1748af828bd841aea2d4376f3d9e2cdb1804484f41c5041cb45ac031b9d830c142ad8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55b6b685f9ad4a5ab71dbc197b59db6c3071a64333c49ab157374b881ace7effa31f4ba466fbb6cb81d64e66a88d3417be5a487b8223f2a93d26691b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89b6ba50c5a168c5e5197b78568fb041927189c16878f600a5467b66c9654802cd0e43a15c03dc00ca6aa1844d2a522cf4999af7c07076dc9bd32744d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc280f752b5d9eac4fd607422762ef4d983cdc7ba4a75474bf57ad6c9cc77218b334275c98492bd0c9e5b984c23f6413f7b3edd6f00f5ddf127cea02fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h782729010537471be72845349545f291d589ccf34f8581c05512137e8ca2346934eb79f2d5a7b0134ee8b7583faa3cf23367f33f3d5da0e87e450f509;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86359a7c33e653ca288659aacb0c43d06bc432c7be7963f5f320ded1bfdda9c120514da6a50768593eb5e648a1e3ca0331f89f567e2a62fee78d578ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5e34dff7cb085c876de635521ed944fb863fedb91a2fb93f04e19ec1da966b45dc680f37f14c8c2bb6209eb771d9e2dd030c84f736383a7b253ab2cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31c4238a54bbd3950aca6fcdc1520bb50250c5242af5eeabb4aefd35099d729bd094c653d920e3f5114574a552685e1d2ac1fd5063df37915d57ed9de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9eadf4be1fae010b55bfc284c2f4518300ab68432ce607d815319e8d5fcf76db62a2f2dddc9dbe39e550b20c8d31f0fc4bafe1cfb42532c2a59ee378f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bcdc8bea3538f67d2630b3de48ce7e8ad72eff3c3f87234b41653213668d67d3cdd33b7b21810bef35769579bae6936fffff5fe0d28b4d2d573d4dd8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h451f1f7c73ef2d7abd40e72c5a6c87d63f95d741080d065749231877365103c15df142ff184bf214924af9181fb274aba31db8f1ec535d715ec86c493;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96106354e5401060d4e8056ec5261085b5cf8943af9b877d5d742f656f6c94453878d0a138c5f6911372f245a40b8431efa2cbf353cb4244dd70b1f23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha50a8886b0342beb828244224b572217ea3ca2ffd6b69f1463a2973ef739e51d4387440f12bee239034b1767244e541541f9541cc61b6c94b08ffe6dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b73a74a03ba6365eb1a993fb708bec4b7eef6019063a9680ad4ff87fc431f3f6e61861bb36023316b38a99949d1ca6193be99da05b447f6ab77638ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90f555bcc05e671a227b5c9f7d30963e03b13b7f8aad69fa80384f10021ce29fcd37c27dce7117728de79cb155b812f53b80c8a6b54af371d12a74b2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63bd4d9c62345e116c48e59a828f7a621c5389e195852589c99827d7a27c8f3ea117588993be0b3cd32bf6efe47d8e2e7074a8ea1cf03887845da173a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1330b4f5831989e130b1af38bd0e548047232a3fa5aebf779e3139e8a43470b4639b3f66ea0092d939399ce3cb88a1e7666dcb2a8449d4a0658251512;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf37097358d432acfcb0ee18a1624cb5c0f546490c21ed43e7c15b6fc6d541a55a20b4f348042d6a5ecdcf40bb025a3ee740ff5c94b341fc09c4da8db2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec91984112efd617806c2310e60bcfec2c442afdec34d4be98f2908d949c81b44a3d24c440997dd62d316d2f1745a4d9bb62f12435d4d8fc8aeb90aa6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba3e8f66f71e5f9c7c1a643c4d9a2388b2538061ee51871ea4fb52fb9bbb9b185dcc54731df79717d9bec5aab581ca28254af4a4053147eb638d137eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf4a394f962b218e41afcd63a67e8687680e3f32616a3d6d089fd4c92118f2d12bd7c560e66428e7679aa38d3ae7170595a2c601d107fced49f999e11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddf421c838198d36f653e34664bfa96a4fd5b0438d8372b808a1908604009305501807c969dda8d8a5766406f0e1345215b071d36c8f0837271696143;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h255baf311a76aadd897e8a1d2aed7436c92ddf772c081eab87bd926e88da7e7161b125ef2fe762a935051fd788745e86d39ce6769d651382a2c0dfe5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2136bec763d5ddd86215e3a0c66cebe01b3f528c9e678763c3b03f403fd934cb0e9a95e49268dd1c42f5c7744c33eedb171e89cb7a78565a44b202375;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd64507f99b5613cca9405fe867ef83fd014cd17859ef80ef7d8d4cec8d6c48dd25d85407b416f55707b5cd0758712dce2815006bddd6fc70e7721da75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54782c3fee046f96cde3fcc0fd9e12f2e3af549ec10f26a160e7b4535969e8225c2b2460775f66b647c49a52a510327a5237b601e85ad110aa1be0310;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b91ce4bb638e5421faf06381eed38511e2303bb969a90c940266b97508a6878d68fd3675dd61859c78ca901e65289eb7f85efecc655b180187bd035e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72ce3e72ffeac2c5d813e4fb96a63775ce33b692068f5acd0c9cd88ed8a8931769f30f30ea49bbee1fe50d67f0e8d4b01ac92eec24796251ae0e1c951;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h538b8eaf416735332425e526382c5ecc881baddffcb2d1b2863042c59cc6422f618f0f9efef800453d47400316999dc7b1bff5a2c5092618e1be6a377;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf713696d562e49f8747449a64d06d8d31e5a7829e219448f5b3383c0437f24e6b1c36ec19f72bfb184b30054ec43ad13b2d52a2e85239af6864206e0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b153a5252556b3322933ae587a7d5b2c65b99be210bbf0644a084cfb7431f15eb267201d9bd122eac63eb8daf0c704ea5437b872ff289f0a391fc490;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5edc5ee0e234b831693baa8a8502300c3618e2c30d39180ea2961ef0c48f54353b4ea96213f09b58908a89747d49b20cbf6c1d28db4dce68b6dabf0e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f5719155d36ae7b2b89f4de33fcf098bedf61f989540cd30d53caaa6355a667320cb79040e29aedd98da37f2c359b287425260dd3df395054703a84f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha874636bcb0612f0191fe309a3e6a2b981e0fe2a371f16d5b1b056df366da2aff4cd02a337483ea6d8a9c78dd7755a7a8ae9347102063a84c471bfe57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6c0f04dca7657780d72e1e9a21039d828551bac2b5ef1081c9a6857415e2ce76a7358b556d2c993f3187b905264bc836ef2f56d000beba047759035a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99e93885e5da9140dcc1d06cf15021b066e4aa8614d987030453696ba25f9f73f720657ab7d94b1ae3c6108b5ef3f2cb8ff811991bec8ccc72fa16ba6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7639030f0eae7db96c2d15f252c51b11bd50224775155c56466d5ad5b87e869d6105ec1273969ed0799af139fb961107e18126a37e1cfe0ffc5c00f64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf32fb55082570c6f6e6ddb9a5347a6d5a9e17e0412a32fcdf6e00af73816272927a2921a50512bc534de42bd4edb90b01604bca4c5ce9a62cc9fd910;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89f327b3f54ff79d03290a41048b572cb0a7300cb450824fda1ff4e5a5a7e5c3fad0f15a2ac9c34bab68ad8e643983ca2f17883b0e4e58dcec1414adf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53e0c2f31604f6b820dda388b5f565faae23d04aa73ffed06a12afa64a3238bd2f9967455f26af97b35caf3282e64df4f64fb9a7451d73b2af5d2e005;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h473a6fd1ae1432c94c94f3af9a12a8c33d0dfaf263aa736538df70be24c5da58d532c9728101f1e62856f7d875649f76580fa05e08def8913041d1fb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94613e9cfa608416abe97f9439301a8e4881d1463d86bc862f7dbf938f2c216ebe5013ea144bc2beb7bc3ec017809fd45219dfacf44469ad18962b729;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3db4b0dfdf93c46ae4a160f4c536c8b6772d1b60593e21680e660c82d0d6d4f5eb8cd977be030dd0a5d88e1fd1c68376d5a3fd0053663b3a3ed1d9075;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h691b03a97b60b3a37ede14b7b80a5debc7de545fe70b5dd23f78dc9c18c893b50388719a4a755ca4e4b43507f0cb2110dc9224ce0988c47e36c871ff9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9640384baca66f5410873abae4c62382dcecd15aab27658ae3f3a2967e7ff9d707e1718fdeb22a8c437ff20be243b65e63d61180b93643d16e62ad856;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0fea4d047c26e42419145898f30f369c6f3fa31bc7fe6906b237eb5b65e04aa3c315618f66e15fd9e603842503d8b42e2fc80c5d9cb10c7e891a901;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fd7a76ddd59277393862ea63cfcc7bcb27b3a32348962c5f8bd8a3a574d99ee91b3f4624aa1bd5c687e5f2f0a7b4d1703ef2d8a4b560981320d6669a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa7c98b88c6e43bfa013bd2048c6e0da75e57b680d6b4f885a2b4616b481b07f8d1020adfcc49838810c926cc781821df0c7a03a07103eacdd7a1d9e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d3406e5803ad4d396f81204363c521981a41f840f986cdbc9dabffb311313fd39ae059ea82b325c56594688683ec8709a5640b9156b76d661aaccb97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he72260e607198a20442eefed50aa2ab9f077d0b60f488cb341db580e7e26cc603ae2628cfb5b5312170bbf30a47320d4bc277a0867f86b1c37d5f725e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb848bf8eef5f0e10485dbeccad4657c8630aa21ad68bf179fdcc897a4fce6e0dd0f2006dc82c7b53252f1ecbba04b40f02b6b9867244c9218f67e748;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h616c3c73ebafdf30dcb92feb5d602d9a872afb40ebc5b40c3d31466ab39959574e7abbc7bbd4e33adf85fa2aa619524e8a302aa8cfde20c33c7e46d2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a6a0bf254ebee16c34d35cfaa4cb465f0fa75d41a07d3b210cb42ab20fb75502e50ab862748c500e689a6ba8ad58fa05b9dc3fa52714d65562bd7ebe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38a7e355b422910f3b63fd3de86f2c37e0f61c683986d97fba846eede39ba53631c7bd0521f12a5ed6096dffa44990a288bce6483b6d382b5db2eba6e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e8ca654b2165dbbab99806829f75a8603779dfe867b59de258f877f71b8a084c3ee559846bd6b241467cb8bdb12e24b71bc29d6888cf9967fbdc2566;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2986fdbd051c2b71d19a9c1a6fbf721ed5cecb94721cfcd024e54065dee28c945ed5ea188e646158ee670886cad31f00b6200b6169906a5349416dc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5135d3f8352bf7adfac270f1340ed5e055ef2f0ccb1dfc6aaa6373439f98023d65090d00ef51e02baf9e42f7305446bf91c49447d5cc5ad094043e586;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc79a08e4fcea9ef8c89ae90a3514b5629db9121c0750d2e2272c71acabeddbe46e7b1d30323124cb6a992668fed14d62eda464ae120324397ae45f91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h693c0cf436ecafc1085ba339cff01ca9cffbe2aa4f95c4294f84e893634e3d61256578a6854de5a30ff761ab8c78712f01eee62e441f858d12085fc1c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb063b398b8061ddf9c61921e767028bee31009a1a42d9f750178cf5ef747eebc5e88a8e708b0d91f634e4f5da10fecae702d8007b9b798290cf99e2a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h897ad91b719776a076357679cb166bb147d8b50ff7ea66f60627c3e1c7ebe5d52092466c233b0cfb4a75021e9640c0b953a5d42917c38d17fbac1a649;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d2e7dfed3542ba6891791fa16afe739e134c9e8a5a0f20f187781d062ffe1ae6d32d7095ef16d646182e36623aa603156882f32f1e4ff40f3290fa9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5a6d140ee0250a0ba532c56f8cf06ddaeed69ac21dd278eba2e78944ce4bd36a1bf3dfec7a80e3f9dbf56aa898a369cf30c1f05f4c934840114b3718;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb90cd4b384882643b268d1c35e2f5071e7ace156e55c4d66518601703ef68f7208f0b58294259ed0e018c759b8043adf265c405f3a4d57d889d6266e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h141820d83325b79a52032b12e6ee7622a1dce78e00da39140ad18f70874bfaf98ce645ff14ee729e884448c8910d8ef3a5f3129b2a62351309cbe919d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb278b3286b0c407adf17d8db17fa977949a464c7030a9794feea22e045ec02be409b2519c7f3aeb7d6618ad1e1f1b06fb64039f3543caecda461f3e4a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc50ea62f09cb4aa708117e3b50aa1d29bffcb00a8c19796792dc1ddcbfa556a33eb23723dbae0c45dc90a068431d2d105796ce4437f7074ea4a382e2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h262589fbb6ca29602a21801f2a94157ad39c8ce67cd6588e9f3c99fd25c499d9af5cc6622338742e96ffc308a5d42e9830976650d3c9938e258d8758c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebe8a87b17487dace4c271051b0940100014bcb87d87567d2d3940d83f672cfe3cd4d2e7cf5a9b8139f516361e3f40ad639bc868472c42a71ee030f5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee697dc40b73f79c2f06f89173ab96c9d0a440b8b80f3388235f9bb9e985b2506f3dd2e9432fd6c8bb97d3314d5c53cd554c1ba17b3f65ba5f6062ca2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a6d315df11ad8bbb7c9463cb93c648315a36c3f171f2b81681c6040306fc973a208e165ab1d67495bed99a481dee09b291c1ce1e37e61977d415d6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64ebe88682c4ca4540f0c87501b91e386edbaa7e7c79b04d30153e2189caea3444befc1bb185837ec1239a898affc8194c550cba2b787835ca9f0763d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bf820fc01db6dd5fb5b3a69ddcbef31da85e6f861629ea63abd3df5b0d57fb14ee0ba4f3dea9fabd3efcc7b90b3a56c48bfdbe7ec157e970ec5c3e25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadf6175b4b1fddeb353d85e68b32af51c7cc742e0a0dd9a34597dbd8758c76056197f91613918141300f7a5f7a22977a2794ae1b12c82f054d743cb00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1a8a771e72d7cddbfa99e5680992b5f0f0233cae0ef4496875d1ad6d7bac070e505f732f9c237eb7ffc8217b33d8539090ac01e094e5d5a2486845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f064588ac72709dd2c45bcd6256f2dcd97e32b2a2496edb91d0b30c3148cd28bb17720cd415bae78ee10682022230494e1d5cad7ff2f4dea1fd05eb4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb914e128e4b1b3919e3e7f77b030553162e01a5ca509a9a363ce57cda1b56684e06dc5239960dcbe49cc8ebe3c2d844aa0537a973fa66f5de965e308b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb693d647eee5185e23caff0da708ec88422c567de16236e623b3b9e0741c312c241213bb51bf62f00fef42818b998d727eb070d9399ca05c3a35c3668;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16ca3e91f0855ed6c90227d702cfce3c01728c8bf253b890b86374b40f6511b7b41b8a2a67090ae0dd2ca1e7fe4530e3190eda3be09fb2028c9842b09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29e4dd0edca95992ef78527590afe703b715487d825748dd8834de263624239d4a7f8fed4198b370ca0e5830489840456134e57ebd2c8ec1e2e33e34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e0341479bd1dd99e2c985ad63225cd175fb229ae009f04237c9b1ceba37526e1e7f12af0ef53511efec850ce2c9eb795f1e571803033327644c1c98b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h256d8dc3fc0e6940582d30e3f03c3590525a935a7f9e5470e8f4eacefcf7aada0f87df69cc1021085a9bd8203c244b2868f932361dea153b89b751619;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e75de59cc96d26becf6bdffe3bed8dfa00d8a6ffc773a61681f2deebc8dce53dd3787192d621d1deeef78a7fe8a38455084c1e94c12c910ecf92ccbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h605c7c79fdc01431f3819f2f96de4ca002024b6a17147e76ef85821be4b419fe734fc684e9712c8ce5db63bd498290dc91cfb12df543c8ded0dce7008;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9a835e7438bad0adc0000427f47a9b51690f0b0a3feeecdffed1fdbd6bd6465e7e0c2f60ee5da1b7d51995b4f75c5298f9a09feb4f6ffeb4bd7d3c2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h950b9e2f902ed304f41116d12d3d2933855ec31572ebd2f98f264569f22a71774f2f46449f254b6250375ed36d15a2067e2f7de030b84b3e99dc66b09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13a86edab98f8e878e3f51aba34de306b861b64324ffdd37c9a7f5137194e6300cbc7e5b6c7952e6c774a75aa09c89f1b632e38bbc4d1a9794a7b8aca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55807581cbb069d22a8ef7e6716c2910a07eb490151c27f794d44efc55052753c54250753d35ca30e18be2356a2e06a9f1d537f6943f64137479c0074;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd5222602716dbae357fd5a10e5986a3f72eaff14eff0ed4c428387578b116823a6b71b4782408689ca0f292a14cb13ca24b6ced91d38d60e9414880f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8343bfcd9eff431d31b16ada3c9490e8cd186f1cef04d73e754d5ff0fbde05be1f70fd49c957b9bfafc0add12ed4800e79a012f71c39b2cab4a7160c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbff5a9b76fc0b05e29011ffc6c42d8313f46924858f9a092401cdd4c7c3f0f996837d72ffd685537997295263512c0e45b50b2ee1fa91a45b8a0070f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc382f03220360474ab7b61c0a0134e70b4cd35424c0d3e3389bf87dc48faf9055de678d7b6cf2ecdea489ea0516d2f2a5cb36b870c70ba2186857f93a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52711c03970d1ed802a4761486e030560e94c98f07dada3552d51b9ffd94952fd83686eb3380596ce665789bcd265aecc12c2af8cc9256447e706f253;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5380f7b9856e14e274d8cc7855687a7f66c854cef0f08de94d3e09ae98cf673ef850f95478aab03bd7fc79ddad1dfff24b6982fc123e05f121d3337b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cb4682aba88b682ce36f03acf3ca12aeada98938c014ed75de8501504a15898e410a341ef17c6092bd2a65d81d841cef4a3ea800b323fd8e93848bff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bad372ca26ab28c6e7b41dce48050a37b8afd69f900ac94770d48cd4e1d1d7479d308f8974393c22610746658a8ecd0a166caa935205faa2fdfb1306;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c440f7799e72576a4bbf06e4c2d5d1b3708f3557ee091256afbb40828a1ae10bf0de87164a96c8a6f56ca5a5f4d007e5c2f81683317d1373d688371d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e60f0fef523c20751a9061e658704340b559f128d507f6786b5da820d4429cbdcc1ebf5f8d6e9db91dfe9c1ff819280995c6ee09495995054545c562;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5060d602daa11f950143fd1a7df13a1eb050fdc4e3e3eed4595ca3ff26172ac9982c2dc4607d09a3c0b3a0a88df1fa9480690a119b92fb7871e2fa7aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h474cae4ccf5c47e9b846b789a84e36dc2bdf76fed7ab309663aaee7c4989645f9b1af6bd5a53e90bac67d7c9c61db5bef0e2abe4cb1ff27140fb45f37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9699a7b2455c263cb0e806a1d65fd5c7b12ef311363b24b9c11ba72aa6f21c228bae2d72335f14806ee20db331cbfc6291c2db89d6c951c6d1a8c1b05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b3e7a5142946a6cfd7eb1bf00cdd3261d6f33f5d9628d2c0a106a1119de767f450bc9f45be940bc589d72b8d602f7145564bd5bd15bd966a7f2be9d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7470da576e54fbe3e0b13a4c33eea5568a0535be7f06da3f21ddc8cdb68a4552824bdceb3e73ead2fa418dffcd75d4b978198a92ff449f00cdc1398;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde3e7b7cecd66757de00acadf9ee6f782230f99eb8fc0c5602c29ac2e2e9c01aef5e0ec88aa286209a8d96e209909afb9b59a9fd6354deab09e10767;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94ff03fba5358e8023ba45f1405b2d348fa74c88c1cd2011a06ef63f424fdf52e4069da387749836139c72648c71d2620da120a317bdef022e9bb34d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h128a754f1fc1fa02e2588a2763ea62c4582db48283f52bcc40fc4f6ed057d3d7c287931ed03da70f8b3b0fd46116de65568825fc32d3cc7cdecb3336;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he53a980197298e4b9066b09938ecf439cba7b15b32dbd53250d824308cd08750c42d55fba528ed9583309e4988c0a4e7b992cd7565096b636ba7b540c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9479472936170cf813945932298d108da28d5776597bcdd8ecaf381aa1181d55ba3a594a7252b8efd44450f15fc331bc760aaeaa4d5918ef1c57fa6f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9475a67726bf74a680b61c2f26d80081a6a17095e0e556849366a94cc755eda50600f5cc6ccff77c9cb658368cb103596b45b9f6df0a821beed03667e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7328d0a2d5700e40c1a5e5497f4d95f423f732ede3fefeaad616bb4ba97f2d833a30ee259e7af23273a4b48437e81ace3d5436b2d283a5e0025f39566;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81fd27dacb7401634d127b5a0c5ad18d834070622cb83a319b4ad3c837a40c4bc4d443c7618495c5ebbc2a7380618dfa5097320c11b896b98130e5a57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bfe84efe9724eef4cfbb66809660aff417ddf1a535270233c913a09dab96b7d081f9efddb1df0c9392c9ac5a98888d38028326450d56ceaf7655e96e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5cefe1b79d76a381d0b10474b3e7a2b85706d6fd15405db0ac6ce44041e596e6857b8f113617df27860780c1e4ce5ae4049d10ed28ef65e048bcafc1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54a7efd2eba16c07f82e931d6d3e05717e3a4b190e5e1b3ec873d2dba563573b5fca56ea80e7b93343355577a034c54323b8ae9e576155e8c2f697a4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82fa52c754199a41215e93be20bd352f44f1c4ac739a0c6ce9e1bead18e8bf7015a6bf141314333dae6a2a2d8f12c4d1b5796e0ba13e360004bdbe7c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef8544bba18a99ccd6fc24f19939cd2f9f91149c337e76d03b868eebb365dfd0654f5786f4622001f6a4f5a99604f1806be88b825de8e3f6259401009;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc25234b01392f9eb3d8123f5dc50ef7104bde40b9a65509d31b0355566c7c91dce8d55e721258a8af2192263f5b13d48320d1a2448f566e4d56e32ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4015923449a05432776bbb253b6e48a5286f4bea693492ed89174e348eeaf347b1af800e1e38b192928d3f8e8ad2ede79bef821fa1d91f4f2502896cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8384b379b2e5b20cd3ba8011bba51c80b42dea7f1f66412a34aa4c18040527bcb6f9a5614101beba3719bf3bc28cd9665a1004af7564886992e95161;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4556e1bcc514c5ce3b16b69fd1c272ee86c156d82a1e17aeaf6e946c815ad717145da3ac18b0c2a75910e4d40c417f8fb3cff24bb7e6ae7afcd7e0274;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde263c1c119db07fe07cad343047baf5ad549bba3bc5f62b176fbb07c52c1ed80d261323c7adf37586062ef87241368e080e158eda538b849ad33d358;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb71ca917a0c2b710fd0d57e246661fd0c719e7ef4698f9cafe8e098580562cda6e42b10ab356436a811403801ddb3e1e7b580fd857ca59ceb0fa7fbae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e1dd2fc0b2cd5421bb8efe61c4879f9d6d73d392aa56d1e15f41be36f6abe6ae1564713289a6fcb254bf6bc686ac0be88c45e4f51298b8de49d9f51a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bba4d0d35dad6a221e0d1f943f92062dac4047a295947b8b5f732c801113ae5310bfd53e4de6da88bd51636d49798dced7b58b9d95c4fef3b93bc84d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h883628948cdbba70bf48cdb64053ff5dac3030508a2b8390ab2c3bcb2809f17ea5cad342412c704184cd12c3b7c6b4ee07df0565f32312e942f4a2765;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3d1c97292808f4af15705866d2c373f453852bae6ce6cc62acf8366458346a70b0c55a6223769a8650a76e3f07e4847aea261736c92abb6ac5495e57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59992b5061d8f72c43e2204359f8a24ca36148a3e4610452d540c6a6362444508c1f1519c25e6199c276ca6eaaf7c150ddc7ea5d27707d2d04dc36dd7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee349bbb0136c4eb63accf133f0f155c935637b9491d7887161dbe4d9c11639dc159707d001ff83cc61c84c5d87085aa96b4dda12128338285618ad3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28ea97e2e48622157453b79b164856f2151c10fea9a1c90999e3613e4401a54122ab72b5b95bac7a475c6dfb5367c6bd4ab7def2ef76a5ca7123b2eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4c3e7e1d403605109f917d871ac8589b438ca56e79c53298f1f175ef9ef020d4e491c088a5c1b858d2c90b1630a9960c9e1eb5b4c0c4b11ed9f1be78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6f6b24a7660cf8616a5a5059cd5a02041484d375edbda255d3e37e9fc64e7ae7fbb770b82a2b667496af25f5c23d364ea54b31ecb63ab247be010752;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90e8ed49c761fb28c8260ada284d359ac1d06021b260fd3e36d012b0f3178f62b5ad78b662bab1d6eb2f62f0f7f88cb969dac1b64b635b008333fbb69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb10deb1071caa097a7a7d44c6362999776081929384413ae319bf33c58158a4230b6dec3d2092a98772dcde7a079bc946c4b0be6a621f21b72c3862ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he49a9b09090846dcbf157d4cf7b981cb65ee7b5eb85c49e2c821f50941885f6026c1a3aef333145de09b4c44c0e096cf6d645eff116fa2049543f5c60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a08b886b49aa80cd8dc1bb34b6787c83a43c492919a822bdf2191746331d3b1221c4cf3eb0e43657e971db59631a17c65d0ba591f8beca33f50e0b41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60b6c3057d1861b843ead618a542f16d67dc5831ca9ec06ce87970048230db475f9597e9327c96e5f076470ca09adf8af60748cca3c23464c81d2dbaf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf9c97228e7b01085a3d5dfdd5bc6db2d2b975d6ed2dfa721ba257d0a083937d88730fa810d83f46a01ea061e024b61891827c588888f5fa0ae0fce3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde8f067f04798e13e2faa081312d692c9bb61e4138cf8335470bb03b6249258d0b61058c4067648251fc29705cfa8333dd1014682274414fd8760ca8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf21fc3fc4ec04ee8a194bd1015e06921d909054ea6a4e4ba040bde7ef7d507f3497ad6ac2346834a7f7c633b7f1b2775109553985a3aac9a27039308f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39a8e1dfdb7133c63efbdbc4de445829f2d518bc964c4644f04dae1299692322b0690b8609850881f41860a632d3777c0304d5aeef1c12987e1eb767;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85a145d19b0bf8cf605d3633894c46b785aa3ff7215619e3237adc930d39613fdde83e6599f4fa5a8450b1d6ee27a25b01794fb869a8db21814af8f68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf01c5ac9170fe69d8fd9b0c19726fc7f805eea5e07990963dcb2cdd1426d4e9fad64db9ed7fa40fe8bd929e9605c5b60a1fec208e42f45066fb16a306;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8cfc55731429010364322e0a828433ae0ce73cbebf2823428ad92283d0f07cf7542fe9b4f0a2f69ec1ae19750ab0cb2c79bbe867b5a9ac9c548db14e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50e850c0f294ef699b2e38c521286f46f89bf983d7236fe3cf0219d5727bb8bd71cd71c7e343762531117b5ea392d1c67301dfd1285b326f25c25339b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a158cbc4ebc5050469ba5a1fc36280b849e1075d36b46f7e15309c8c4102adae0d1a11091834617e52d3e2880ba0253346686864f6971c6f6a33170f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f660e6597be2f1e95144d5aec095cadcf754d742eaf1cd1c0621d492c8e7598a27798dc4e053e9f9fd8cd8bb9601b7cbe9a07296e1815aba565c9345;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ca36f4dcab54fb1496b5ac57616b9197a4d2677602100446714146191a31f24aff9fc739844b549de6be4d126c915223e93df03d40c13f3e321b3472;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5315419af2df8aedcaf437985ac5625475ed1d916579b4e794b0747b8ef35c076cfc0bb1b4cf261458321ec236702905413dc6b8ee27845ebaf5e1368;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc778bc79a5be014e95261d5717ae7637a4aed4c1ccad2747349a7a03ada1a7c4f483eb0382a4ac3188029fd76a0dcad625125fd01e1712fd51ed1ed1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a18185c266d3e10802c39717e94a8684d1f03f6d8b3561ad9b2fccd70341a5e22dd7efa7f47742835db88452ec86ec692b455179d9cd0257c7b6837;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h854342cdcb5eaa7435ef71ec7d63866940c2c0a4c9907dc6280e0cd84dd3d043996dcedddb4d64875dfab823e14ebe1d80c15bcdff45e261efedb0439;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ca34a0426df93a80393af400843dda6976fcc32e768688465be1e3d71056b8882aae902501cc2f2993366789ebab21c71a70371df1a12018e6ed650b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fbd3b748300a81e75ee728301fff9207494509084ba8778b9d101d4e09b2fa79b49d47b1134967add241b8f1dbbf87d2415d1e1364391bd44d29ddae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf36fdc14d91bc5530cb43ea1550419c42b83ae15a96771872a66df7bb1ec0fcc2c71f6f997928efec6b593eb7911ac79ecadca08f4908222b7ec0b9b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37e5a5113eed1b6b468630c116e6fbcf2c7fd987388a6393c7695a0eabcd0e9a8f671ec81fa712bb21e3a2d82188ead40d954b4450fc34c70cdb3912;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc6499e1ef1921e159d883f84ee803b3e9e228ddcfc65ba71368a1fb060f1cb15bb0d656878fa4736d973bb6a3157ad6b3e3ae4ac9ee5944bd3d0ce5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5da865067e95d4c5366e78680321dc99e0c8b234a22d9d257de9259315bdcbbdca540938cf1379254148305f19ced4386c34ba43671884d41e6fff645;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5acbc876daa16a7059c53c84022d071bdb4433acc5d806337f6df165bfd6c972c13f4258740c551db9f1a1b0b492da20ec58289a1aefe18bbbe8b34c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h645656fc0947b95df4c3c92d6554de008b56231aa6091c41f0bb3c8ca05a136aafc1fb2024e42776bd1c482a3e00d0baff78bb88db33b8e653522fcd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b64f1bba106a735fd2fab9f75ceb3da340f01fe775693edc250f4027c6e167a3ec7e6bf94c022f34961dad6a6e1e915ed0030efcc8eac7aa3e66ec93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8011adcb094966ff68d3c74dc29ee6419ea6a9889d7e03b17f21e77f2c9ec35c550d8849bb4954630ca81b01be6450a964181057c6e08ef4d1c79cff0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h947c614e870f140f9e6dc86553da0652ef35772cf1b1040e415276e4ae8ff27d22984ec3520acf67e07ba4c0085cd6b600816bca68e3726fdd7879f7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0db5c2ee508ab780fbc36099d5cca0ef5f70ce3ad325bb457b1fd5a48d42fc4696f8dcfd9f96fa25cd9a51c20646c8542f713c1fbf714ba3ad2d4cf7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e2e8ec3dee0b693043bbfeef817a20f8d951512575566dafe342f7d0be3f6cec4b341735e17fa60444cb75c55cd6cc66e1fd23b30b078e845462c835;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68e9490c9a3c77a9a4715bdbfaa87faef7bf8c1e1502754def5552df03e15d9fb645a1c89b3361ac39cb5b1efe1a4419c02241fad2845e50823e7dab4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he98355934863a1af0c8c8510f7929c5ec4cb7be1d3a0e61b472f393bb7e3c20d12279bfc4958cd0e8d616b575cfcb836d53b935c80c560e614f47d4b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fff1ee4a8d0d048811806e21ea3cc19fa8eb5dc04cbb1def7cb40bbaef927a50b30e5e8843ca4e22b16e73f923a008419afab2ad105fc6afab874685;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80e122cacbdcd8484f419496780676ac4c6f3062b86e74ac9222b849a292ae565bcaf02b4000a10c786bc0d727e3e2286fbfff4bd9339a6116af4f039;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd4e09da61cbdd787d25861315288b51fb95b0543910a02cf5acf80d674f018d643857fe3b30398176a58a8cccfa3b12b800a07982dad334f0a7c1de8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h875e86675614ec4ac54d94d20a7e8f558345677687f5b44a756369816dd9bbe784818a2061c63096d130499fb18c927e5dca21f700672aa22a7240a3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2212c89e279b68e743f772c7c308a0ca211ab344592dad9123afb52750bd4c46a5e5eb5c07ff5043234514e55871a4b95da04cf69abdd04ab4b97db17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d7e6a64a52ae5aafefab2633eae1d5a616507e59d1d1271c6cf0054c80b1661f10563ca35d8d2ab9a6925d5cf6ba8de411089d7550cdc9420d9e282a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbba612508d268a2bee8b41246e79975136f0c86ba6ef36bcc49b3a6ebd2dba3cc7f72c5cab866970cdb8d90bd2b2cd1d0635f4c6e788986e39e8e35f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9abb943dfdb18d141736f5a6d40c3d9b948185667eb901d53e1ec9af2c30e3ba671451ce2d835bbc2a5d3187626ddc3c66581af3bae4d152f8942925c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd0f3f0674fa517838fbd03cb47cc796a2785e125a11c9b17d6b9762baa3fbf1e16043beb28a5896e9368559f6520ea57a9ff7fbf4ac3f437dc5865cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf79d2456585b4029477e28182d05a2a3bcd033ce306bef552f9492d6adfbf8a4c4ec743805146d7abd8256999c51105e1be499419c322dd646c7d27e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4908771ebcb2442f874e74eae2d0eeb232389cf6c0159162456e04ce75ae33d86bcd04d924df60f88541c1b7ad15edc50dcd6b686c1cbd382bd3df06c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb5f73d47fe9840e46161fb907241f89867a3a76c81b29137bd7dd94e16bb28054adb6a2eaec25122b5bf17baa862626c947476a84a7fa8eacbb61e7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91342876152813f2b4948f69aaa2db22d4f91120d6c3a5c9a61e6d626552b0ceb085c9587e84f77b32cbe00dafb2c74d175b6745c02a2f2d42755e91a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41f516ea817aaff4166e66e9e1b9b732fc7421366b9e1e1337472942e35c01bf2fe9df9eec2b82d407b930efc8745eb2fc1d57780f52a7226d3ce22da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcdcd3d998f40f394a62be1b69f44e2b2a46b8fd984257bb21c215d4df587a1f5c759c0f44382db07bc105e84d044d19f8fbb4559b1580745c685d14b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8fb8d25d9adbc8dbcdbad59706b2243c8e6fa3adfb489cd7efe9ee2da60520076fcfa01711ff463d3b9f82b6fb74419ca4dae9cf85d6bb9c17b20029;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9d11534296ccaae319a2d4c01f0c9a8d3c933dc30705dfeeabea3f6afe0a6a10c65a43a80a59be7f77b3bf0ecd82bf9d5199b8ad4a54a544eb601726;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b6aebda7e418ff6cced616411c929310e32c2f23ecdb2fb11ee879f191fd7948fbb51eee8b045cc523e39bfb9197bdcfdc5a07e03c3ea1e9110376b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39a319c8a39396d46b3982f897322f3cd48a22488637d5ffadad2384726caf5bd005e92653bd9ad0dc8871e7aa5ea6ebdd46db5dfd3ad454a8a24777f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c36b7518eb6a91621099b8d29d4907eb8be9a7e019a615172a0c13dc5dd9d02a33f09244edf124899c13075b07b5c0905cc478f90502579443f0d661;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h378b771299bdc2210ca7c01c358842b2bc95119ec1a3f95ce34feb283354e6fd9cf678256eb8e6975c30106d5078d78ad59b97c7acff0a4718bbbe614;
        #1
        $finish();
    end
endmodule
