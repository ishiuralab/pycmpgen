module testbench();
    reg [28:0] src0;
    reg [28:0] src1;
    reg [28:0] src2;
    reg [28:0] src3;
    reg [28:0] src4;
    reg [28:0] src5;
    reg [28:0] src6;
    reg [28:0] src7;
    reg [28:0] src8;
    reg [28:0] src9;
    reg [28:0] src10;
    reg [28:0] src11;
    reg [28:0] src12;
    reg [28:0] src13;
    reg [28:0] src14;
    reg [28:0] src15;
    reg [28:0] src16;
    reg [28:0] src17;
    reg [28:0] src18;
    reg [28:0] src19;
    reg [28:0] src20;
    reg [28:0] src21;
    reg [28:0] src22;
    reg [28:0] src23;
    reg [28:0] src24;
    reg [28:0] src25;
    reg [28:0] src26;
    reg [28:0] src27;
    reg [28:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c935a817a9312f9f7982040732f886cbc4e6b7e79d2332592227041ed76f9311eff42c528fd44fdf40378ff3ee7d853d1266d44fc2d45b9794b91a04afe79411e99a49a1390dc07e8871e2a4d6d129873d9e0e121534a56fa5e515b6a9bf96045ce01ca6bc69190b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha623be4e1df591c7e62a5a99ee7943bbf7ea1a59162f7abe0c4958a388d8b102c412b84bf25f514a383958b4119f6ec32a601ceedbd461903ae929644bc3080788d6d1103a0ee5db2624e6485a0904a25507aefb27f6e197bf6359f3ecf9656535dc30390bdd20338a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a538c5614717409e409f28af6b06ee149d6be2244ad0e6c63e057d04401adb4d7382983ec2c313abd939c4d73d2f75558ab910e14ab3fb11be4330dbfeead60d03f6e3d079ec8bbb3fd22597083cab8bf041a20ff9fc168ac8dff9ae3e3753178c8d233b7e25b58d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb3caead6c8e722410d68e936575c759df257ef7319519f9f7b313e13c0841b5ee04b3f7ff39348bd651b4771c9d07d078dd8a1f723e749bbc0cbca4ad4d50525b97a208e7b2593cbe8178a1416d5360ddb912a7533ed0e9cb4e7cb7452dcaea8f9297f0a8566184e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10969658f5a346549d27f3c874fe54ed7243733329023f744e61530aabe1541453d86db6c375cfe91d23795e24b9b7a6e34001edaba3b800330c613a36e50a4eea09df8b94b214409d887c5c7c1bcc1e59f390371031030d2b46b5958b3aa9e7b16eb7093ba6e4d433d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ea8aa1f8c1ccc2aec53db58c33ea03cebe93e900fa6dd024f1bf6ac27914e4cd1bec28da82ae8e3ef045825c201eeedfb502cf3e1c33da909cacc002e0d7582f985cd875103fd509531fbfb862c205b895b922aa36add806f9d6b3320dcabacba5078a331b67cf60a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h29bfaabe159c821875e51564a012b26a5f603b6ad5e689928cd210f68254cc407080b338b68c0a6d6b517293846dbd7bff711f19fc833812008de45997396a5c54531653dde000f88963c673e1699e8528222076e6f6afe67e9ed4091b473e54a8c3561c11de26d326;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb02628dba09f109188c7e85a43d63d40470cb55a0f4e5e4f4ba2fe60d15866f86623f6f4df725b4db74d76b83344def15914f9c9f1a052024457cbc81a4bdb4b404d85a3bc746f389a03921ed35af8225fabb61b05dc5966ac05b1428b641146c2932b9da0b2f31c96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a665463ab738c660c2748475897dd45bc317964f8bd507076f9e624e7b06dad99ec79c03006faf66d0775adf1e672a7a8f044c2ed42e35681b4171882d10e37980393a09e31c147385becec197c3f2f287aad58b68f84fbcf5242ea0a876595d4618e82231de952da8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bf33ce730a3ad225d244a32228e6a374cde0974a79ede054fc67d53deae5faeb34d7c870497efde0b4af496ddb45a1175e139071d7bf3ae5d61c9fcd41277e681b2b0287c744a30ea398a16a0a1ac71bf8d45288b91737f1cb027c6044020af92d8515c7fceb65fed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc01b6bd3c41d8425e8d2100563852e3b97f4d48c5fa619600b508465dddc451ffe046cad901fee2340d9cb4c88e00e7b0b413efd263158e3a71ae4943360c4e341f9f1f9c1ea6f0815fa795242d8584333a25a088d46627065b39f34f93137653ff3e2d9ab4e874ff2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195a38f5aa91c1cf1ebf47e12c636dbab72886856b370eca5d25c31684e0605908604a91cdaa3cfedf32b3f5462e11ba7a7b01afb80080f9c0686a33d0a74861e35d35ad941c38598019b20b5a6c350c1f69805ab29fa982d0a5f00c05454d7613778978c21b359dcfd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a967a43ea67f12512e4256d19d8848040e1c856127eebdf328aed6cb4f9a176ce64893ae80da2c9411a7e25251821375f17db8832e941d9714e63e8b33d6143e05d41f8a72efcd2faf8f26db972f0a0c0755f9cd6422b00212d22f4e11447caf4262669053f8bc57d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd36bb9d4444c4aecf88aa30f1c576e994ba81710a98b887573452a54bf8b17a41f753d841cfa76f03b87731d8f1406a64c4cd70222b83620756514948f7b92164bdcfd4ca8b7691623f6d81978a5404c6c8844d16244a6d7b1b52162684ead2c2b2537bd300f934509;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a4beb4c93ee2b37687b89b16ffd7859b79b1e85d3df68f6d5e92f71dd677fe2944aa6938cd118ebd20c15c5e7ff1f2050f6b3531e38bc3867d1951ea82f1cc8c169b135a1671c84308f84fb3696aaa8e533298f0ec1c899b4b0110d9a10365693bd2d750935086bcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbcee6be5695f02806ea44d90506d68e835e65e0a414e423fe510586ca11bec8358445290fe9180d672a182af71b27542e6cd532361649be8417b445c3208bfcf5e145cc80fa8b92a1baf41d935041ddca91cc6d28f6d0f43ab92e2ac522a8046ea7ccbb17d21c1565;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161a5f5973bd1083b2f113ecec39825454946faa8ce8e70d3910ba702dc6b56740469b013af8f50ed20367105e7b22bc7ec4aef5e5fc6e6dc7d68a7d7d437d4c0460870814dd67a09aec6da9476c6feecacddae61cb870a52cf75bf110fdd843cac9982e4378e44afa4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ac30b0dade58af711597fbd02ac486e610d1f171649867c3f8257cf8787cfc99c5e016f70bc4fd22557741f7b653f1680be6a4811e91c09b3b93e2d96f6219225fb2734a17261b00094a38912f5c8320c5a7443a4749a26809145891349e005c2ad0d5fa7e92ff84d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c2bea4b7eb124fed33416ab249b5230ac9fae5049456bff1fdd462ae305480d2690b38e09b3cb6cbfb7095a38add4b78881eabba3588ee5b314116d5205e6571c06c848e41c62d0f2a0b92a795781b55505f17824564bebcb1667723ba63687ddad02f158296d0e38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdbe1cd9acd483dd8cae1de2052686483e39104c8c102244cfde151379c42a6e1c6120f7ea27f9a973bf706e07cea00ca3e7cd9bedabe798def65f1b7f5b78f7de8e03befebc34b79a939fc73afc28faff0385ee547d5c2a2f736b504235393043639a703d07e93e0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb8743d6e261605b67ac692f200eed5ed14b17b34709a7e52ca6d515364cc364ade2dbb4c1a225eb82e34f0dfdf35731b75c9d39db11cac1b02778cf7d9f2be9bbdfa926957a9f5a321251cb4ddec8d4f4e87097b3ccfbd366ac6fc399b7526f195a8f2fd1bfebe37f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b846c20d41ca9f5526327199a4200411e1777465ab8824496e49cba83a17f2b9a15dde21d3560a4cdf9ef846999d8a22fde7ea080b328caf6dd7fa044dfad0d0d61ead0c2680ae26982cace403e7a901c4de4cf7c1981a5bc14c674fcceda1d97d9a5d326b0985354;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6028f01125806f04deee0bfe7353fa93c7c3052d50b7f82b2f3a6fd0c9d5840f5853ab0c4d5736b06b67e5a684a369c6fa2df39abdcc390e1b961dcbc0736dd2c380f6df43c2f06ed634fbdbb27f1a6d11692ea0a2f45dd38ac918c67e04304156fdf383267aadb3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166726d9870c57f5ed9952362beff3ee5a0183819b871691a51fd793120ba6c3fc8e9af10d6cfaa61262df4b7f130ea9faa9f3ffe513b49cd87caab97120f2c1af53c150377d322e3e616344fb8794ba09982f813ad2c76d8f6385366f66324f73597b6b5d29d61e1a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6a8212934554e775677cb37a6933d6477444275f9451ea39eda65d8e8c65adae25a1c5194be03655c4a8a2046715585fbc6a40252f56a54d74e0b4d0ec176d2237b5eca02a442c0f88f27228ad0adfb4458028d5b56cb0d37c86c3caf44bbdc85c551592be1577be6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ce488feb4cb6d5bb9570ae774d5a2a3348bddd85acd28a3de147f01ef8941c66809a79353fe1bfcc1ab3e12cac89048cd89ac5d25f952fb180afc6e22c61c603c83974f9a2338abb8bdf3d450c5b6a2dd957159fa1c03f34310066057fd3aed6704cbceaf7cff9417;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc97ae43dab91f51df110c69c2251239ecfa7d4078a9828c0aca162493ee3f126f26ec48598cc55395616f6c4066e9361f971a1757eec02bcdfc59cde7e0741a251bc88263b4509a48bc10ab73b7bcac7f238ebdea36ed506fbc63dccec7968f18fc660b2b6488f28a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d3f40c5093b117dd725f45836fe9632c497ff3fc1df35f5f68f5bfc03373ae9f627ca72a5706b80bfd14148046d1195d42a78cc5c563b1dd7581eb1f6796ccaba6a656666421a364af7477037dad7ba86f22cf8977ba707aca8f7fd5cf7917867dd840b7efa29ab5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e92c2c8b93ec4623342ee12170780a88a6eab4add03c5cc9a48647b8939f7bc2543f326092fe993cf0899bcefb74892d5e080a027bad50d152dd100ba7a25051fd0c1399564b59ad11e75dcc71b07fa2209203702051d231a9eb68de2ba91515492830d107733430a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12523b4dc1de516847ee3f27ba855756aeb34d6eb9eda3c42ca24da56126b9f70ad01c181f488940dbdb670c073695ab681dafa9075cfb1ee0352c4eeb206440559cab75033268bb6bd5125d6b1c4216f95f2998b1e2e342f35a2c57a854bb443680e35007cfd5592fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98a486749ecf69a092ae8addc023cc9b9bf0d80ca78609677b78b7dcdb0da05f179a438fdb280e49b5d129fded15adcf981cafbd4bb9ec8f2066f686a13f3ee26632560c502b340b08ff96a7c5f582e9c6e199402abbed52d4519f4d54c5330833e624bb15194f84d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36d1a4b024ccd501cebe2290ff2088b86951ebdb34fb24f45fc516a2c8fcaa11e180cb721f54bd0034720cdb187901ed699cee765233dd1239030352e48d4c1090b0265a8d4fc288422097e3353290207b2d07b8bf6d2262cd20634e2ab16bbc8d6ba4924a31123500;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7855295cb7f11e433128d16f3cf72780574309538a5f248af3a0ca5cbbb38ab4d0cb34d2d58f91509ec6037e165b5ccf7901e3420d3d93cd3e4111fe3f892afb7377992391ffd74dc392bfe53c5b388b2439f85bf2ed6e58de9484006224d30c9f2861dcef98434539;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f53988ac15e72179dba00386a78770d0807e5e7f411400c1e70bce1afebc2f020f9161b2f9cf8641818d70a275c17c354a6daf90bef26b68a6bdfd924713acef3216f7d13bb45099f742702c5ad81d230eac38eab54ac662f61945c0c62ecbbde88d9d7664190f756;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h929a1c62efb12b9b109ac08250376f6d68b810d5ac934df3af97999e97417be663830f0ce580bea35eb5950d1ad5654d75050b8d515383c879980332ddbddf1f52355e29d176fd760343fe4a5090130a21791121c2bfc440f374bfa29475ba1c30cabbb4fa3f936ac7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h347425353145f41f7dd7f4c16ac22dd35893263b99485280c355c2e768f5389a1408e3a8d65f41a7e5191b1a0defbada99547b5e719795c78051117d6d15cbb728ceb9bfb9b0bad1700502c37e74f4490a20b79edb6bb1da84f2a71fb211d8014b9c7158396656c016;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b7235f2dffa8f28085a79bf4aae0c5d58db0f5817d61762b24275a22b35ad687479e73249c221d69bfc143f4342f1766901d3a8bd4b460a8f8996ebeb9bc74ddfbc0ab3024332f1e37fd3301f7dd1389cae5c1a00628405fa51cb0fe8422624006b510ceed87afed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104520af335d0d3cdf4aadfa6bbf94eb596feb913a6bc623e429a9c1e9471a80db221bd9978705bc24b802f340fb864dd57d292d5ab761e0a9bb1f850a71c9a75acfcdfd8dd6e3f1880544391f08ba62b332065810a582e4307c200a2a63e9112a0e113b8aec425bf7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb82fda265a8192932e558c8269e20bbed526ac4574814d039729baac3f00c28b17ec0c04205f87f107b8be6cb73b165214e73e397eb7acef40dacc21ac2a04fbe4b66630ca30194d59180251458635db569bbf616c57ac260ccfa2576ab7113653b0567cb437c4d35c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c469062745a75ba9b341ea7f84279e5f45e45e320bdbe881db180930208a66d55091692b22f9df58affd9aba495f0dd3d93f8a34ad29ed3e7e2dbebcb7c229a295e0f99acdd8c5f22e7866aa4811645f4538abdf6fa4c7a9232e95dd413c0e5cfc9501f7bc2093d951;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12074c68d760ba381f4628c57cbbfb52b7ba1bd23b5d1674e47a233db0bceddf8be205d88df684d6b7ef7cc88051eb90a95de797fb93094786017f93840266b69923fcbf86336dcea5dd1116df3a831b8f3cfcb8734bfc546f91523bee3e41bf7990cfb6be6f72ac370;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ab4acc3bcbb8520f26dc025ab31828ea4febf51800e9587f17898729478b7f34f90e5d91f8fe6135fd8dbf7a5414076e9240303af824b031529905f047149a77e970bdcd6a534599259401f666e1afc718be9d6c5463cce382047a1898348f297b0e8652ddc71cfc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64944998df94c171e1d4b9cefde76622e13efa354d78b4f329a070efd5ea19ff4da355e766acdbf21c856fe6e7b649287d1b0c0a2b5ed0b96a7787d2edbca5970f28f3b31b356921c5c5f35fbdfb86243e44f096528f8e25e3f14593d9e6bc31721c4039a082105c26;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a34ea9530e4f8e8c5328df13196c203a6892650ac499d65c22c60d62ee2e626433efa6d78ebcee8208dbeb1cea551d693b0b1491c929cdbbb7e4d0a01e7e148df47ca65e1ab8a59ab86495ad9d08e37c5b8bb44e36beb463b7f01699cf413bb768b7de0d4af2c77cfd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2becee6ee764efd6322244ebaccdf99dfde65b19a40652ecbb8f2cb82f7e5acd8c79fddf96d2f7e78fdfa112a27feb499f9f9348489b1f149736bf74fdf8d3a528661da19d1242fdad7eb7cbb0d756ae7b6c671f04edde244891f03342dcf94a1f595c5bdb3f51b13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d640c5046ff3bfe5a55c3a9397d9841949b25949c9867feb1484ea98f452d62fa434430fb1deed4f35c93d4789847ae666233b0d7bc2d328d11ec78d3c9939fda73ec0012fbda6a0231b4084f712093af9fa966b9acf04f527c88807bd8f72ef83ab9ae72ba636bea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcbd0fbde172e27f8737010950b80fd423d166c49f2bf7ca5a79d67848533bde7f7cdc36250da9a4331fd803a0e9f9de33818e016f9d06cec90ad0b167adfface5c6348343b2aa4e66628000633c63786e84259f193447bce1a72d9b30876f20fe6ce7400491cc0c962;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacb4f9e47e24d32e93b664313e33397025d7f2f1b4c660d43282e9405bf6c19c3b40916ecece067758cdac2f089a5961ed5781c4a83ba2563f35f23fe57051ea8e1db90aba8fe7f0f50c95deac2d2c4524c644893c0b49f2ebcec3f890a8bcc507d10941b1dd26dbef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5fcb368f781f913d0c3e6847774ffb52f5964bf36a3cb0c9e1349dbf751f80a4b31095bddb6b742aa1d56f2a3b9d6e5c80e0489d5ccbcd7a0277efdcd025d9a46d07b2a58b6e9263ee07bbe715c30d0b74effcea62e42d7551594d676027404f50d3d54da568a7d4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e7de3f81a72f2012f6ee753d30d8dee0331f7728e74c63f89b1080b39833548053d3419ed10eef5c4bb6a629c464feff4c29c2afa77e3ae6417d69dc89a1038ee03898955cae4ec3157a1d1913b95b97e2d8b648aa44690cc10a018841a48f441440cf616c516d792;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d08e4d15304d95ac54e2d62c2f43b5efd32a5d249ecbf808d92ab62edd42d47055326995c01e4c32dc8267103a3ed9edb29abad62ed0c11dcdea3b108158b76809fcc4324ad4a23586e17c0b855d44ad12b9a30b1321c3f309122aa3e552acbf588429c008fe132cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c78a6015aac9a714280e3ee9d76dca05f335ad1ad4c58331ddfad32a9f03febed0f8395dc909440a2baf1224a447994dac210dbcc589e1700f6b3d8139f7b9f4e095826a969b26181252c853a3636b508ca44c0a487a3c974bf8637fbae2ea4c485c4f0db1737416c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1104cc11696a7f790f2640c36bcd0febf6291b280b86749580a2fb565f5f753af205b30fa44e4100263954eea3fb7b290c97bbd4fcbb2b356eee7343757158a18d1bfcaa9110069ba758e424ddecaf3c2bb44957929a2ae5f2b0fc640442337b3c8bb5aea82777ed847;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c16aca7be3ac2ce7ce3043ff020012abe91c548aee4ebd64f5785e1b233fea4cef5e3e5e0a52799dfb5f50c26e1d4fa0bdc49439539cf2f9af0db1fd4b9911c782c05f34d2318882afda3a0bc4c71c712c062cd4d472203c453d7745c6ebcf9aa0df31c942490071c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9552609941b93d36e84a4fadbfbc700deae4be073e5170d1ff37cc4b1f83024c78b6f5a040290d0aee6f4529024f659604836eaa42e78d0c3d0074ff5ed6a0d9246187d80ba4720ca2d2cfdcc87f5e67e8d0e7485b05eff4c8f97edbb028a4b8de2cc5f08f7aeb572;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1def1b1c474667863b61eeb7542ac31241119f9e73296ca32b23f8f601dcea23a57b7d76003ddfdbffe26e618f5eaa5416e305e07d6c0d5b7d8e542e0fee7141995578f6bcadc7f3f65c6a70c2e1414ecd630877e1bcc066bdebd77af74c717924ee8f035fbf85fa11a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172f4ec5cb8844fa200e3e861f596d3b7bded718bcda65fbba6b540cf7189ad346f6a434cff540ce2c16e5e42b1d2a74e15026177e8f64b2fb978f57c21a134b3c3a11df630a1abb6227372f27dcd519872f4e97244359eb74b5bdcc1acfa3981d44086b648a5fca9d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a798fd885d9721de78912a0d3f5061845276aa91ee2b2cc6279f4ae27ecdc6084dfbc85e98e8e2e1d42acd637a2450a8f88df9665069d8cf577127479bfc949bd07524ec56f5fc3a3a79c47d74e943c4038567354bc8fbea3a93fd4a4d6022d5a3a343b7d20ee99ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118d0164c376ba5037dd20139e5118fd75bb61a358a1601fc762151fdc81454844bfe885ead85933f1fc5054e47ba39c4d9653da65fb5f3491906765d153f212d1325b9eac37247e7df5431e0817272ffa81ae7d965d50a480d0168b4d83983f3dae65e68170f7abe00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcfe386459f9dfe1734e6b804fc5762955f78a5e0b04e9db7b2f52f95402df63d27286e48da2730dba0ba3562f4731903c66be50a203846ef4ef12ae24ca65fd12bf221388722b4bcb64f72f74af853c4398c76bef9a1e707811471a3680ed8733574ec85483dfa6802;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9375f46129d5274d74dc0b1782fd32fcb7cccf6e1a7b3025a9385d81986b10116ff898e10456e7b8fe58fef64497c6493aaedd40794d9cc36d8bbc4e08d6306ac834ccc44dc52d21232c1714e6e8afc155df7c3207dae152eaa170a10299f63b91c02fd67413d6a13f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6ac60d565806374f814b087b299f7523554f6a832317daed35d26e49092887f05d9c47fee0111a15b71d04041c12997155d7df7487326980f182c70705fcc626530089fef43415c3a39d75e646a4f090d4f2cc4860981b419dcbca74a25ccead4a8911ed47a91905;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166c29866446956debcfbf6f921f4a15cfc3e6e9774e1015f89077a0c89960c20786414cd92c5b4fd0bbf536af593042c8d5f405e7d5d8b841e8366c155ea551b24b5e4e0aab8fc9a89bf7562be86aa0d007b09995087556dfbd84045c949822f78b23878854255213d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h610dcc960b188e811150610ee3f2162f36532dce6ef3ef9baeb7b6f4b8a5ac6da35e793066f9fc48744bf055069534d9ea5307b2abc77166543dcdacb3c682a09337bbfd6fe1e57fa0b8dc128ed273869f3103a489fa2731413e02b2c3630f7711873655266d48871a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he734d145d514a1a7ca0845d528029bed45bc8c5d58ef8920a7166b36f0ba9853ae203d505762125d0bad90ba8354811c439fb13183b36abdf610a3d6f527ab6a9d788d216d735a4e8754154465163882013625f67c643904e5fdd6163eb76f3e2a720e1c0851c1616f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67dd4e575f935db485fee7b6f8d6643b389f689cb80a948bbccbc7368c51e531a1de461d66957f08ba93c7a42dc3e728a91231ef47a06e283a13447312fb1d6d9c19868aeab3f0350786afc3a405ae7f099802f85d03043600900199fa3b560e658134aae3e408f040;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7758fd1cf976f16fcbf61eb920607787c09c9515034db4f4a5302526453f0ebcd9836c1d735f37ce0d1e983f7385f2429bfee751be3828a682365ea62d58cd7c340547077719512f5eb968eccafb1fe6fe0345ef849960e434c84658c66523ec295b190082d455bd9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a746c55c5948b357c16246e8df9ca46b5af1a2c6fb7a9540f211e50eab60ad221449fc06f7c7d58bc68d2d2540286964319ece9895eea3b9c40b71e1425a60699063699b67e7e146ffd0b254204c2e241f6b47479480c2232f7b3280327b7ac6ea90da24171b15b169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haeafcc41ef3ec36fdbea2c76db465416f980a62728b4a7ca93b1b2d6d99acc1f1426209028f59e8c4aff66e4bee9ad633db1dfc9547326df90cae0a192e30dd79931d8ff117bba55df8226b817dcdd95b3746015a2998eaf7b50ec6f91216d8b75cffb5b78698b5057;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1376d629c6843de6ff6abb5048903a055284e78b400e52e6f2486e8dc288c0eb13a01bae4703a13ca1000457fb5eac7822468afa151f50bb3fbe6d68679063bebc79298624e749d339ef7de2523b4d03c0a172dbfa483b7a4614931c97677319f498c3027d9aad201c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6040a3b0f6347b82f1a61ba5c1f13c4a6d6bb6d845da686e87285ab18e89d49ad37fee311a6d20ef6e4efca87ec85b148adf88811cd6fc02aa291f434d319244a07ad15c95d24a1d7d018ad30f54fa1b1086f9ef12039a02e09b92f6c9610563d54f656e229fc91ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h683aee89e971827767acb05839035920156a1144282896b775240647051b17e747514b0125b810e0a46820ff79e007f13d6c0ca157995f364e9e0351ef7efa2bdbf145f0a478260ff7c00b6396f7a21fc41bd140b5974fed530a7ccab00ea100afc82b7d89b5ee5f5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d35f118bc8dfa5867f4be7ad5e4a68181896f17e99d79e3289bbe4aef333e1d1b4cdee80d3413f041b36362af39c13c0f7ad9deedac0ecf8e421a892c78079f55f70750fb16c76c25936193d8fe0a77bc76fd6d59a9ce1ac901aa32b153978c6e00b5d4087abef6151;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16dc140351b53e6faf8c44ce8b398bfb89eda52357bc5df4eb97e8ad2db0b6117ea04febe943df2d592571c32b94a4858ea27bc6ebca9b8b96bcb54420363a6cc9195a8d5f276654231d8adae1ef30009eaa5af657f5c297dda6d025cc577a989ae0ad8eef2895ad55f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfaed3640c933dd14fe3d2ae1a5f50675a67f0508444babc7408e526834410236061fc702b8e7eeb4ac415d58b1784eaf59857b4fde96a5b0dc92f4a573ce4b018cda275b893145ffdd509b70c585df5f3122946fccc45e283a72efc95edbff184b1fc08a425c8343b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf6182637c4eeb290d76eda80f453fd39c86264fa90a3cc46db525a6cfdadb23bce456afce209d893afabf26aa664b4e345e697f084e67c80541dde2d4e34b5217c22cf1b00febbc77ee9162391facbb0cffdbaba39b885f66d2bc65edca994e895baf214524257e9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ec259681766ebe6f7084d2351d649e517dd861aee97242e11742ee30970b5547cab36579ce78fdd7878241d3c1eec04507757bf327701a353e2a3b28c71f6e1f491420c41548e4c1c28f5a7949fba13686e486dd9c8c760d9b5e6b87542133d2a63a501459b39db44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0e6dd3f9ff695d8167403fb0a8a445945f36b0efcd093ba33f324181625fddc4d18a8a59a6f04d250b700db1f18c5abab90068afa9ca941e3725ee682f1db3a959fa6cad4ff4b55e91819af87127a819504c28f6109a9b9a43320a28ed42ef47e48f5112f81febcd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d091ab4b4549a04c63cd76b11e95f3f46d4ba2173fc604b11832b3bdced6edf0dd2e8b142acca43ebee0d67fa6106e3748f180eb67fa9e76163f14247bac3765d7d4c7e1d7d105bbb509d712b6f04e01f19d1211f0567cfcc67bcecdf0ecccd6dfb0194f537ca079f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4c27caf45c8b48f820c726a91021293284a8ba78cf5de5a0cd5664b57fd0546123405a86611765999b2aff37063fefc967e22cc54a72ed78729027355b647f91110553395b5c2b4b54a3ca30c22dea4906041e73a07467cdb121da5b53d25d70b7358706b7807feb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13bcc9c8afee79482855224c0f34be7e996e04dfe5f2db5c2d1917d1cf462a5bf2998e17b00c2c93d8633161cf2c89f42cf50cc46f0ffd882ed6347da566a047ac095c186021852d3b172c27f710d334fa23602846c5736f82b5e1f45b1492a558fb6080aaf8aee1fe4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdc5f869cd0f644e7c404534f320cad6348ba93a45353b3d55d57381ece53adb27c7a006b20d1827d52e068e173ac54aa184878b40e9bcee065ed299f87d628dd0ddcd61c169edba95327628e76113c7e9bc284df7bea8ca11d19c63b6d82a1e5b52c4b61a35a0c150;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdef72ce496cb8d5cf1e498d69759e29853b7eaf4edaa2af803a871a7502ce3498b51207b533b9e0a769d3444fb3197839f97bd78927930cc11b7786bceb6892da1f12950c454375c8e5f463004e07e39a59a58029e747c6b9e61f30badadb560d0eaa687717ba747ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdaaf71790a686cad92327e3a088293c38cc0dd1a78a2836b815a33f6c2a40ceab450bb47becf571d4d26416c378df07555efaf453b35e2b0b27f7b546652ef43eef6d6ec72d53654e23d4587901e30c8ba265354605355e01724911187188fa371e3640245e6664f6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3dc849c6dadfcfd523c5b7b944c61fbe0a0777f7461cd21834f3c467e4a772107e1741f5af111d36a9c62f20802529466143b22d3230f3b105a894ab26e4096ad5bf3f6880abfa8187cd50087a4787cd67873db335b65f454d230859bc8810a39dfaf3cb8987fd379;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc295304b04af26d01eb19266b3ec93570b5a1d7b5d675fa35a6bdde966b875847f9384a7a8290ab9c57cfd4d06dd69b4b48ee0f2ef3066f9f2dccb87b8b364833311a0ab9c8f9d7bb1ea6575b850882f7e5cb9f1257a7138db9706a736f98c396d5997a8d2b7c2522;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7442312cacc8b6b276881658f564cc8708500772847c9190220e3748d116a62c02ebb5ebe6e35fc8d7cae58a722e5a95980ab433d6ea12f0fd48a90a085750408fff41dd47c61bc8e9dc6e28e63bc8a9b77a7db2aa478e1cb6bb4db8f4fc16df1684e65654b0c815a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecae8c373c9e1c7589c76f1a497384ed4f195bf8130788250f1fa88307775780777aa11c5b8112117504061a560b9b1621fabb3dc51701aaa5ffcca968a0c4a988c5ec883cdaf138298080cbebb7b778fdf098a9ceb14e66805ed6fddf98f81bbe9f29b3b83b49fe1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h581bc36c3180eb9a38ea18c96f82e027ae89fb79965e6735db75bbc62e7df0b630eff84e581778c575b842dcef462d2fa33139f6360155b7cf12486ce0ce5ab5b0ea1b4a311d37158247e3c915beca2e8351e756bf5e8c8a0f47d35fabfd5a97dd22fe78f714c7e8f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef78d8ff421e34d5cf6dabbbae02a213c58f28907011372c50cd5be7db3452980da86e11b7892cad10736637f36e8b11daa58f48b01304c5d27b6d107dc2f7bd01847baf4c11f741848ad6ed478a1c5369277f12950629b42239f171dbbea9c402b8f0179fc446219b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105c9b76448769b75e57b4a0442a1a751dffb853cdaadabcc5a725339882002cf874e81528912d3b8c5d4a92069f45399a4dcc5cb9b2464daeaa10a290676d09bd22bca1557658650bbddc17e044539f6c55aade559abe161aa47b6ebc38640ac2cad06c41c05ee0071;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf649f1074371ac9468476feb2bdcfec2165c2e8585139548378d8e08305a81e862040162d8f2810b97a3193b344ff51a0e4646e6ac02119acee50a83e0477a94d9dbcaabf5983135ec43aacb0a6750cd5fd763c7e4df07c5be2270d549e8dfa5739655aca5b51a86e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10dbfa0b906130f54d221fc948a7a337378b9d83ce8af9257415d772525e131bc9748dab660cba7410453bc941ffbb71700eb62f5038ea169888c7f5b0ce3a5e1a0a8758ac41187acdc70a512c3419bbb098178fed566def0f381c85418a85eb028edd0a108e2f7702e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h714648762e302a03a38dd3740b4f9e514c7ec188d316a1351a06a09a1ab4752b18e9c803e8323899b25e984db90543dd993cc47d56fb247c47d4799f8608330e9ce4ea060c5db8036618b2695f9dbf99e7422a9d075e8179385aade5dfff8de45b5e9300f382ec86c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18349f9cf15bcd4f79ecc91126081d56c92c33366e00c2bc940f8675238c1c89366863b2ce972647b8e13bfac5ed888e390a7c417b16880e0e5a944d2dfe7e2d3680e458b567e599fe53515a211b48863c8ead0f1234e2f4e75dfb12675e0c1608ed9d56bcb8324f69d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14267d392d6036247a7619c34e6fc157433c85efd3f90a757fea69053660777881a02ac78f246701d81f5cdb260688346d05ebf3865fc3fad355501c69aaceb944f470f62becc3df3355c5080ad80fcacc345e571977fcfa94c717075e57844578e7f402db7feb9c59a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b73139440b1f3e90fd5ffe7a7e657720d7bafdc284cbcc844c98a9bbaacd0c428de03630b27f40b217b3d3718d9eb97665e00b0e2fba586fc0a69bce9edca241f173ddca318426a0db4e0eaab0088434aa8a86720ec9eda4691ec2045d5ca77bc1913e3dd238713499;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11863c3b7f0b8495105ceccba3db5dfb8804bbcabd72bdf9a3094fe527d1668f804727b3cbcd2720d5dd998390025abb9210b976c2005eef4fb114c7bfbe05d1d2d713c7ed5c96288d3d5687c67c2c987e2be672ed4d8dcedabcc2adb7fd71b4f22b1cd541626a25f31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f9a30dcff54e1e52a5d5e54029bcf39f6dfaae3dd1aa2fa2dc282e674ed06d3534702cf45fa85f1418bd26385fdb4010d88d0489547cf86d95b235a1ddeda8297ddc3e890467502c4d902d4c6ee5d07030e081dc4e96583f60e4c47fbff4bd37210316c6129256dde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb383efb416e803feb0e0bc5c34c4778c76e51f801dbfaf19f43e5958f6c671be480e9aae01b75c9caa8dcd20c3a914d1f8c31bd8f969a002a0cf081a200c5e0d498b158386e9b3001508ea841244065f01fe78f7764c03e6209e085d7bd8f01067dfdca8a78cecce8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e406a75faf25caf05fa0f9fc1a1977e1395096dd45c48ef1805352100a3eea2a54efd782109da1eac7ede6d8c5ebbc5435bf5018f2b456ddb27a2e0c42b300c375dc57247e2e5af12b04c87a51ad31a09a4e41c7365754f8bf86c9e33c387a72cf33ef29d5e7c5f91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ad1cd4e8438f3005820416195d2025c7cb1c77ac4dc1f55204d231464eaca1bb1e11e9033264f7c72271b4e9cb0f68201b2ca436de6a74c69f66a2e283e77e3ead434b3a9ea24fe2ac58e49a571e29399cbdafbc0e6a1b1ae9a0723dd8d32796fc8302acfe92812f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76eb170753333e0cce82848e4be38cb37bf2abbff8530f8b9df78ffbae25ee8767877d52d3093edfa66d2e607ba79b04ae849c8b8394436b558495d0b03be59e71448019e54d4ebb389aac8220ecd689fa4d479adede679e1d5bddade0c34ab40d15124274ef13f1eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25fd17df7567c53753b61de68e007448f34ccf11b1e42b9271bf9f25385f1c0520bb5ec946608d618992e52fce0bdb7f18890d73c62586b8723f209673a5c90eb0e5f3fd65fa32c46dd933a1e7400c4963e47ea31ba2d7437ea05b8822e7ea4ffa57d15a1695d36770;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27199992d8340a67b149d3baf546a50bcd005fe113d2a855ee1c69a27223ef07a70ce939599123a1447e62aba1ba6cfdb0d4599054c910bd8d90a0b96ccc94c299ebec7b932702c0851bca786d3eca758c873d966a29acf599a98e957c0d43abbfbf0f20c077cd6772;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcaf938b44a3b43aa440419c26c69e1f99fad6c41b5356b3022e8c4c98eba30ec3a995da4e67d582abe69dc38b1e5a26d007df1cc92926b761d81ed8d8b6ad470eda6d0984dce3f241ecbaeac6492d9567ec23492efa544e90cee0e1c38b05b4c61723ca699e862fc1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f7e0d3f9f45eaae1d5de54a6e93327f2abc7b798aff8b6189b1e86c0d11c66cbd8d1f2fb72a8075d06ca4f53e52e47c13e19c37d484f2290c286eb392ecdc190a27e80bd8d05831294dac5441fbf6cc5f5411379134a07fa62d23f6b323608dd2b26146bbd62016d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee1a7fe759f9f0a532b931d14431598b108a72c5c263c1150a0a33b1566f7e2d987e2668a353ab2901e161d49e00dca42ae7268048655276be50c5d06ea78b46f77c33f99e2215dfdc7baaedd912b6b724fcc187a8e1ba5248a3e10efac30d4d88a2a7a618aab7aec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dec1aab5c21287f51bd6fe9c70f37f2a20400ab5770e4573a0a6afbf7ce9996248d631466c5f886d61bed51a63859995f2f237d093b81d0fd9247709806d8583b966c12ef5fc31d1684c0069cca22dd7e0e8c4d8626659692b50fcba73ac3b73129b6d2bd9928b710c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ea24b76d0be7b635a1e23a0a3afe3491207a8f081670877bd5640ca48820a995f311faaecb448905ec796afa0714ca2d5b8a6aef63e4eb32b5b388219532d519c8915e7ae215d6255054b5a41178083d692047aa331617842aae8a1c8dc8988bbb1291380f3340f63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbd045030fff993fe0ea1880af8e2ad252b13e229cbad9f2bcffbe81b73f55ba9a6b2a09a1ca29a0d2888243f7e697fcaff0114cddb6f9c5d691b2a1b4762be6d9fab02a280525c06c6b057283eb3d9eaf85954c6ef231a3dbf2a6383c78a982d47f992bb125affc45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93893657188045858bb5f25759f1064d1d8b887ef343edd99ef08d3b01184b3f2cd983dcd248acae0aa1a6daa40e9904f5653932a9ba4c7252cb2f6034f886e1e308a4a78037c3d2e3ae9ff7d9c0d2123b42b591c700269165adcffdacc7de355db2402577f36c6fc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115accb5b07a899c708c511ef46099c0332dfcf591d0dbad456295d703a9b75f3ad0afd7da061012739aeb0b664d77c3750f65e2aae6dfc24600e02c6371a2af7b4ca262328378f7084bb58f6c03c8052aa1291741ec76975ee37eeb24a1d00484e5c2e07416ad9a2e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e4ebb5360d1df8c1057665c7045593df30a9cbc12ce5737a21b8925063021b01f608f917108047d3417867334f306d1542be043528f05f4f710fa375c46709660e7bbc89b81ef74a16f2ad0fde7cbc417267bfb13be21b307e8ba5065c7d134285aa3d4f7b9aca654;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c36d0ea4fdfb73458cd7ac28adb35fc227275126f134a4924b2139cc28475bd616c5026c3ff4077bda7b6d28cf7b781a17f5d0a40acc6be141581b7bfb497c8e9cac2f43d08ff0d69ad8865a1fed9da8a43b3005854636f72434f43917e2cb630d170d751dfed4ec68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c92b5dbc65a35fe06fe882055c891f928280675b511a947e03b865d7e4543b4c025e050abe3dc091dfabe39460fa9fa5b0c3133da29fd3368bbab1212004ad24cc167c34b0dfedc1ec5b7a0d66619bcd6e1933eb009f035b6041ab4a7466adb4f1cf378202ce635320;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153d9ebdbb7963267787db39e88104d597f3b25767feaf53073f098a008cb73be9be460e02113acc114b45bcb2274290f529b18d2c6da1964dd0048934ec6f55df2ec2856b11ecf31f6850c6996d56f3f0b557377bea7ed60dcc21c5e9eca6a4a912af3836980e91e12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10178cdb176665ceded5cbd8ccc739c725994b2dbf9370604a43a3b598138173111688556d124f076d950ddfb5ef81162b3ea9261add36a4399abbbcfb069a93f5f30b04e3375b3f9cdc99adc8f8e610fe7049b103f692ef75fea63a5fc86af0a21076aa753806f5456;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157a4e1dc33c30ab45195f8e13d5f7a12ada91cc1055f69fa129baa0b68357d194108e3a95297596310d9951f6a298df768957cd7aea1739bb164b9c3a3a223fdb555b7167a2baee5b34bad823577cf668762f5ec3604131affcdffb03f7ab6793226fbba06686beead;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f08548db8f72986caa84f2f7e88fa8ba2969b34452dd12e14262fac47adbeaf42b25b9e4237c1d06e5f05b09701b75d0b7613840df973f40830944c75e2f35e11e6207f28ba28cf0ff1c8d5fbdb0ac973efda545d5cae0058a9ab3876286378dad7868c45641dc34c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136f6021b841f1c4a65d8e8280bbc98d1c34845a53bfd5ea14147a946b7c57b227e930cdbf05edf78aae9f37bbaf672a4557b707f3668ad7b5c9c89e95376ab86b8abe5b2aeee540853423cbe08a7797be68b274a891a1b97b6e0997c1420cdf2f61f782f22010bcec7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3891e618b5a91b959f18006028a067a0be538e13d188b6883077ec89e12cbd1ad526f594ad100c256324e8d6ca95cc2eddbf16fad39791f53d55bddd36263984ca4132e2ca32eedb05f4c9c6a9fc6cbc16cb2c691015cf249b2ed1d6d6004bab1cdfca7686bd81c3aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1837967d81a4cc0079ea0587393bb6dff7e11d9510c515cd7a5d81e58881a0fc74bf80f38b40f3bb1b20c6c5bbbda3f636987ab13824477abd30d844973e45dca5121da71b914b5a2a27df1eb86d1db8189ccafce43973a7f422e4aa740b98021cd744c1691c9eef69b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c32a2df86d99aa633fd774676586837e77020a60407888129754824349f83e5c18d98635bdaf7002219d1e5c134cb68a7a9062b9bcfa5b412c6f4b6db1336bfab65ec6a97853fc080be5bc461a64cc7e4b6d96c3a6c2d5bf574ba93997dd8254ee309c419d73e8c66d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c11a40e20d8bed35ba678b689a5ef86daad0cf39fd4bfafa0f0cd827e3d2d701c451f4fe1168b2e83fd1edee34853d56f04605db102294e4fa74379e11a1e3a273c97f26bc4412c8a8191749cb81e3140c91aa630f877d41fe52bd38295fb3a4262fb589cebcb02f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1321a58ada8188087eb6dac6b72ba06c539709e7976dac0c7b3b7465d763b6c8f4d12fd9a8e3e7823af64bb0eaf77e205ded15df81ed8280b13754cb5692828ac548caffd588380caf578d1d58f5b3547fb365014cab746c4101a1d66a056f38688535d69e1df94d05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc46660edb3e46561ff823b5cfda86811ea0f9a2f59d631fd930b38885e22aa9e999f1d72b076458edce5ad66146368de1feabe57d0756d9b3839412ed4f6c008dd765aeaf2203d8c8aa6bd333c654f4347583337139437bd2243301b6ba5aed3d503356447bc35f23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af2420cd620b302005acc0c55a677f8f9a11a16bd1fc5fc78b9f6818e370896bf81245ed8be9df73beb8bda7ce7a37d03a355934ea99b1c4b22cbdf8ac4818696f54039a1fbbfbce3009da02001b66f1d58058a7e78521b1c9763c8e8f6a0be026eaffe886e3293f20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2bcec2889c2eeb09fd71c44b1f8855f1a625e4901ad0981ac52efd6a0bc280a29f862b915ab1e2852efa73f8ddc873c0da302a4e45c69fed9c2559a0078ca4b2ad4cdee7ea4417210294fb1e760cc46afe95cbd0d5cd21a1ffe2805f112f9fcf9b5ff5381f9d69b05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4be12aaa0d70eefb8f3546837a7060a9f4deff27dbbccca54ad1cbb67f0ae88a7d4c863fe6d9a9b8821e26dbea1ec828ca97aabbb42eb75eabe2739e6779e3b73e0e768f7c38028fd441361696808f9d962992df37d06bea67db5cb642f164b1f3c391cf3b040b7892;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c910324b5a7b08a65f8f64cc01f5c80f0a802d4d98e837eff7f7ce1a2c60aa0405ab2bad9c9945a5e9a5ae316290e29cb9dee05470b4112e3c08af927618b6c5c621184fd0371b543ce2a4bb2c8e2e9288de4b4008d937471fe7a10eadbdbe8a233d8f8a1947b9187;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180355a339c5e81c412391a314049cea2a3f67342699ae47dec8f491cefa9d2e62816d6872302753d6de8aabaf4159d0ffce0b61dc7011b930ee9bd382dd14cb14dd5dfb62725db1fed161cac34e77522d0d4beb2757a326754fe8a41abf17a03c076475d88b4b4a868;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bd1269331ec532c508d5db428c8787058d869be8803d8bab445574b95c36d81c293b927fe24819e2f53354e44e2e7cc2fc9a221af569b1505eb0cf69ad4f17131d6704bac586c621196b581a57964ea4d9b10ecb2abf6a05248e421d83f424231b24639f1e54bd56f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b54a893d72c3e80ebdcd09fb7b6bb0c59f2a9da3dc42e45b71bb647a938047ed60a235dd42be519ce476cfa2e6ace20c856de6c4abe04f2f05018147b127bfe11b859b61b4abe71708b2a086976c0d3fcc5d7c91a77efd01a01bd76bfb8549efc0afd9991536b3aeb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb0310cf5eefccb1d9f02875bac399d50adee968ca1bca809a8521ff8d5c6c5f1891bf317918e571b4fdb0df94bf7decd0e323b3cd01d9e673540f889ef6ccef7486d8043da59f447fdec455042485d3190ac44181d79ee897bfb9b0f3de47f7cb8be9ee8f4f2ae5e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21780c917023324a6d6a2a917e8bbfd87492de6819ef05bb7a79ec7887a2f91363ab0c90ed0620f81d4c9653702a0e3fe4d27a03fa8fca0f8d6ea58df4de4370239d714f8d935a577c05afa949f3bc6b2edd03380bc1180b52239d081c221eda4174d2cf0fd7f75a4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7019e2dabddbe1985a0a80bd372b407e6a97e801ee16277e41681fd55b14c2cbb78f78b8a0d7ed97420774e89212f6f829e2cee882a3fbf5d726419592e4432c8907723c3fb2a3e8b3b17708a041bc9ebb1fb948014ee7b5453b1426745de7e20c2df26a4fb99b8f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7ce15c128088ecdf0fa770f45227b73665f85d9f437a995816db43b57638c667c7e507c04d4716c332aff4f4f882af1987cb7e604cf704dd90cd2b4965aa7d55f1b8f504d7d8d70e690677f4a15b1f152b2b5de9a06e2138f6018e1b796560837d322f5ff2146faef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ba9dc835118ace3a3bdc083344246dab85b3cbedf976970f860bcb45f05ed974750ecbbd93f9687648d7f2b25ec431b89a0266fb17c41dab99cfff6843dde19ef8ec7c458378711660a10ea080f0e77b00813e384edddae4dd35a3c455b9112beffe192a5829a86ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaf005903ac82f3ae8152fe4a9b5cd6c6c3b3b8d6dc40ea228263d6d4f1d9ce8cff0aebe926ba52ce28829a54422ed72f1b2465794a782660346e7153ecdf86c8b8597da67381f1ad98656ef03910cbb78255db60afa90c9efbc22a9d5185ae84e6c1689da96a28c39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha73c5621b116fb6714bf7078e16284ac054656f1b60c120a22a47d26975117140ab16d370b325b5f85fa430ae3115d94b4377298b954b5f62824c232a5908a8a3c8d3556eb09f3f0fa69876d6ea1fd3455b7f8be99a82f1a48c0fc21a69f10786b8e6b0e07c055f400;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b221841f0533fcd3f0ac6984306887e7e72127edb0b9bd803c9039754558686286b8b50e111802e1319208ca2803f20897f001ef05c87c06f24c5eb100b4cc60999176c55368d7993cb25e5bef517b0e3d43107a8d0708d486e2fcfd430257e75577d410734a2ac1fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd2eef791d4f866cfb13b3b8dfc70981301a73c67b6ab2c11c737f3777bbc67b1ce17923e51152a9ef9706e538a1536aed17284eb3a9ba103fc317795041dec5838d1098e53f6b0716609f73673f8f7c6153800d0cb1b98c949ac5aa34270cc6fc9da605c643feb918;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95c1f7cf19e41ad9d5a35a4475772ee4fd5a9c7f2bc0248698a3450baf6fdfbb24a4ace4800cb7a24d853e5b2f93a439661ef1cd2471948675d2e35837cdf7b5761996febd01db6cbbe95f606ba8112ee3477ef5003d900ae24d2c2683b24edaa633e22e40e3acd03f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b9cf61cda9065bf4168e2c605258929728e0ad9947b4ac3169aa08c76f8ad6a3cf4942ab26e9e9f48a7183f5965d4762eddb245bdca85cc69e4d734a0ff381de42f3653370b6eb44cec37c5a8f4071fd81fc28edaddc0a7962313c137acd41b468ebb1a78e771b4e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a29e57d79b21e49b64c582e09cd7388c31d5b814ddcdcf749f879262f8b1e0256535f36a34ac7b29e58615328678281be983342cdeee94bb06edc6fbc9c6c781fd7bee05bf6251300450c1ba88f92be757c2a23080e2fb3df5f3dab5af120e24c0667f0e5aaf7eab08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab82d82ab0cebeaa8f925f01332bdd85fdfe72066e10f0a2b097532f7fee15d7a8b3ee7392f2e69396646ea00233b6f5ffedd0c1167e1c50f7a52501e1aff7d759142ae48e26b6eea9d11847bfb54076b525e493a851745015022ff7036e417e2db9c4e46efd2fcf47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189f0c13d1d7152a585601cc35c1fc917bbc4165f3f1cf9760c9fc7e60ae584e5fd72da2b86abeba504278a74e121c46efa57552517b0eb75a41c2545349cddaaec27e42e19235aa47c45ade8d1bb14cd633630cde20c3e4e12042f5c0487a4c229aa2079a3ed6f6eed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha813910f4a55a97eb426b42da6f149680026af3bd59e38aed90406e7ac5f5abfd868019348f20047976a3a7fb00399bd464335fdde2605f14945f08d83f89e32b3530fc1a98b25d75afe9608629eb84ba879a4c01d842881a10cbbdda062c40c6a80583c7eab4a4da6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115ea8c61a29b94ef3695949c09eccd0a53936cc44edce5cc82defd2d706061ba3ddc4fc434d83bf59c41acbd8159fc27a59c5582f4a293827a8099eade37aaf3100bf3fafe322ba60fecee22ca8caaf2a80cfa0a0aed401d8e5d6b2f0df14e3363206b59a57b8c2f6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbcf038c0cff1c63be56d702143e70bf6ea464e7308ae7a793000e3eafeaf1840c5ab5ebb1d895a90c367c7a256fcba9f151872956c7f97c272c43fd0676bf5377eecac4b2e2502d1ca407c88ebc60eb4f2d7db32998a3d29aac00bb92d6e7fbeee875ea6f187c599f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8ff5a20c823ede7e58f3c72fb72a5b2831c26cb13c3c0e277377e49fcf1bdf6e2d43e53d199a9b64e25a8562ad311dfb66fb1b3b8ce746b8cf2ae6c99332860641fbb46bb06f1b2950e320ddf7d4b199f91d05196a152d88e9bc1b701ef14fd158a90804fdce1730c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd4f4e24f480a65d20a51ecef2ea28a1d95e9721f5c8fe8f6fb3d0126e87ba5c9eaa350edfa7c756ad95237892f56302e305cd1914192871be8ac0b77a102dc0fbb435961468c349fb774579dadc2bf81bd3c8b2d4ff484f198dc5434ae852663d6c8ebe3cf9d935873;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eafa4f6bf16d6a2e5285f74582e70be08a7df092fa18f8a7371806019ddcf13e53a4220bd1ca536aaf9a01c5e0172e2d1b594f85d4c99be17703a9200853c0af5f1b2273504a34fa949667fde87472f4e2f40fd0d24ce7b3802b35ee2b95be237ab23fb0bb34cb08c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1025f5af7d7712196e973e5cb9b430eb360ab1159ce96e4d01222719452cfecd7a01e94490ef446a04d27371bc10b48410559121e859e37f88b2302540759a4eacef33aef283fbd292b9ecb549cbe1f89d95ddaa6902138a9fc05e85ca132e25f70054b10e09b0b667a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he43bdbb36bde0d169153242cacc3e504b30d54e4ef22e5c0d3455cce4e28ac2d06369ea6197267031ad3e0f8e805ee0ab2d8c91e959f85c4dce8ee3dac2ae386e1d2c65f59132cc110c46ffd811dda0fa21e0d20143804ffe58ec721e9e15d9741f398565ca8fd0f35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d387a6dc085c9d4302663fc834117e44aaf3beef49f88792d7d75f38093d347f72adb5dc0bfaa401208349759f9d4d02302bd6c798d657b4e4db011d780129e522fa5d0d9b86846e00fd6d2eb44e37b884ff6306c272f1783052660cf0d3584485e10a1a858d4f07a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76f30646f290184a1f6437ee68fdee862ba2e1cb02f4aaeef3311552b30a38df0042b4bd8ec13c7db0015ceb20da6a5ea03c0e8849a6ac9e7fba4ba256c0d5df3903d7697546bf8d812e6fe0522187ad732909555016991a04ad7343965ebe596b40e5f2fec27f2aba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164a08ff706929d255daa85c34dd1224f94811167ce97c062fafedff2f505062bf9d9979184b09f6ef5db162c1d67cdf67de76877e04703b11b12725e420ae2d0d1afba854d8ea1e99b565a7da677b83621ac3e5844dbd36212d9809b9fff6bf28948cbb684e2dec939;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3db79209f60b06ff9cbf6b42afebf404588b880f7d396509d07af12ae77944d245ae80f3db4215a976f0eaf7fed4e43f4a03c999dc03c4ffeb98e63fae768989ac1d2e21a000c4b2398116fb736ac8e968543bbfddf6ab481694c0ea70a7c94f6d7af5ffd7a5788c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132431fade16c078636777166b2c86eb345d9f8552df803290b85991f7e01a7fd3fd12ba94e17d45b2ac53c4c65d03224edb8aa3e179e29b4abbe49ab19ce4cbb7cfa5048ad85c59155f8fc56d505baa9d5bf38cf381dc68281a8acc4dc9f27a4bba2b5416a0e13fd0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfd57e29e47c04770bb618a27edf58003cfc36725027ada68a11938ac1edaedd8e21feaa6a3be6016f24346ff8da753660cd1e81f95f1b51f015d7fada401dfe6201bbce7a3b1b0da9113cdb39c9a363ae14dd939866a419aa8678b2bbaf014f790cf00db16ef2f1cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb22570f947ba4d813179d54878ad875eb027a808263eefbb055bce51957878399a6eccfee285b7ebba4b9686b03148a0fbecf5287f4277783c32feed3ee01d5774eab28471958f846d8284ec9ef25c8ba7c87f917203c9796fd6ff77514592f51e161dbf3581bae62c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d45c2f500c58e5df4125bb0e0bba7c57e2705ca8380aa09a09dd79bdff855e36f55baf4d09e8b75feb41ee681340ba67366af5676247bbd982bf43e95d79526b1f2242dd046f01fd4d1625b16759713e5322765c64d690bb3abced56b141f0ec1398ebdfb74d39b1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46c6503996ef071e1b90990042701177b1c67899e15afced9b6c1490db521d24fc7d784b8ed2e8f121c42ff7a40d8062fb97dcbb1ba433aef075a95ed1757f85ebffa40ff9be80a373f8456e07e6bad86b647f3462773305f1ef3b730cc39f569adc4bbc6a392e1935;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a052507025e7e95f33dd176c05583dd50a18daa8bd10cd3d117fa0849f2235a4e81c3c03bd84af86c6bc6f0039f1919e5191084d483ea33208866b880ba2339518fee5ab28ce4682676d632735a535f35e839a5c737516226f884d10b23f6b218c162aaa1cf249d4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35d6b72c374260d3da2f9f5c26c5210fe99ba82cdac2567e70dd86afa1ef82b35c3c2d9705073a4efbeaf59865a7255b18ca20815f5f074895eefe2904d4e4135164fffdd22a07fd22d7a3b14fe89b7686a448a91fcaac6856322d3943a2f1a479e40223bfaf79dd41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha340eb0d467be941547bdd091ce4d91e912129a77559857a2aeb869c7ca2b0e9942e1fed916438f90329f52aaf4423d8eb03f7cf44c36fe54ca5ca24469d55f46ba345cafc764f60d3970381487520424405cd78a9c7502abb53533fe766db45096746ddf637d59bbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4051cbb3775916adf6df8e9c27ffaa1233fa156cd6a4b825efb75f1140bfc6914d106d42ca762737481ddaab1893d920d21d1c7cca4e400e75f65ee1b65fb527eafa486552c5934f734c9437123523cae44f5e5e0bca687ead0429b45ab2d56a7c87e9471e82fc550;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cde3a820f0e11aec885e428455a138183b80a7f312751101cb02343f2399b0a6ac6524c424d8e962b7b0c0249002309688c375f4321f0d4f8b6d8f00c0d2ca98afedb7f89fb5d6c5b8815d342b6ce222047adb5e8bf8fe08a08dc62da2ac8a76f5b0046836d0ad501a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c62119132b227cff9e450f64b506e572c6755e366491183c687f3d9630253d0ccd198a4e173b5e03c284c26447c3cd20b0acac30eedde8a8156384841ae149deeafac8dff371e7acd8b25def00ebc7d8334b41cf28f17fe6d67af0b445f60aea0b86ecdab69cf18511;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e07da5a940fc40628bb6216167af43518c48abdb183c1af203b1b35cd9351927bc0a7410a96f9f28bf65764ab92e907391a0266a5666ac6f8c40ca8d7af1a92f5dc344f3e39eb9de38713cc0965b7e00a2a8daaccbc7893b9446e6a7748a6a455a9baa4fa5fa80dc43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef4d3007e5d2679e5ff5df9b26234bfd35f1183080076da3db9ca82a5514279a007981dac6630639aec518aad2f15272d6421c76a87e14a7e0c2ba030b70d6b4d55b0e35d6419c54a475e545bec5d410551d07ff84b7d59383f5a3d486029d3f74dadbe8a455ac58ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9d6d344f256669a3927fa5673a8e38c9edbde6ec7ff88548b3d7882fa5ae4254209f4368002fb2500aea93407a582169ea5e26a6de5eeec67782193fe545c91187262a30319422f5c16a7317bcb53f6220b04b5c7583b4a53c6bc654a54f1f80f4cd342c1663706f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h837f1dde780f2ccf8cb331f9d9f846181ec02f0eed4ce0df8dfefee9233023b60230bce82159306eec881107bed712c0b404ab7ed6bd5ddde6177b6066f73da93821b117b84ebef21d70b5d0d103c4597d436d18520fb78d43b4c9d71106cf1b431571fe8dcab22c6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da3756905fb3411c20d094d7377f7cf375ddca6e72933e06f481b1e367c258bbcaa4f98cec8b592eae69e4851555245b3c522cbd4e7d8cfd860011058ee14af52d871b01c4563a502e46021e699030878a62b715e019dd5dd8a88cea56141e9c8034d54e46ffa47abd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96116c636855ba79bc7894b3ece687ec23af5808d32d8a61df9b8550ec8aa7f7aa1af13120ffab84634735a6fc7735903a1b6cb5e4d05e004c9406fcf792b5a748535d6d4518de3fd4ca60e2c4b0d7258bda73985f8cdc576b9d3d7117a949de0493c648869a64579b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddc4903526ed361b2d20728eee4fcd31f535819234c524e4e010005946d734b61d987cccd3d48cca52dcfecaf4ffe4c587e3c163d478f681ba09ca2a44753b8af1c74ec20822c0ae5c436fa1542bd60a9a84150d1159d90a6adefb3cc75c2e15b004dffceb23fa3c8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h585961d31f7d849b77b65873c5035431cd281ff717d4de6481b2a27760e0b5c48036f644ac4b036b8027bff17ff99795a74db667f7b46a5a7a0d725a009a53ba983cfdb642dee8da5f8c0ec8a105488603bc508513c535a6cf2e7d44bf8071cc29fa1b3cf281fae3af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb61b1f1e5c340c501e4ba610303023c9db7c7e1e9b14cb191ae75ded6a722d916dc1d3a701ce6a5cb1fd0cb3676920f2d187d5c7365ef05b88190e00ad6d3b41efd6591b36add2f714a21d8178eb25c853a0659b45064e679a2f8699d6835628c2d2e7a4b93d3b07b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4cab22133c6dbc293ac182d8c9b334e740a480187951c4bffe25126b5fd653920a92f48c564f662a30e632b0b0590880349f3dd8d4789c4ec216838daa687482d12a7c52ad01fe529f49ada96e082555b96221ec36d6413bd3e7811194b3463a8f2a58a02f53409a17;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e9b5a7a907ea5c8fde105f4896f416b9587238f2fbf896482d09943c7e3e77b60113458e4cfb9936b9788e959718b90696319197585bf1677f1db8b72815a887f781cf336443e0caec3a70556c1f06cf8f75076016b8b01db95acf4a55ca51639875a4d6b42c66e31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3116e5c26380e239c2af80109f2543473a0a9183baab9dd4dbfc10a1d060eb7d1e19f61712a2f73d681d2b1661218618ce7c68446869c8adca139295de70f2f088d9d7f7f75c33853640ed36851d6c03206232735907ae9e59599e5977f05b58affd6bbbbafe068e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e846298e86889aac78e8cf8d33d2a86c82015d87f678c97968daad7f51fa15ac9ebece2d104e613df91df3a1e84658d07546a7edb51bbc9465eb6d49c9752e3f5a2a9be6a291bd119b29e288204f9fdc7b3edd2ac6c709d7125fbe955352485cd6b117ae12f98257e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd46dc93d050eb5ad773c42d95faa027847b5ff16c9ea3a0f5417a1d6df75e5984a0378a65ac2a890cf20f9b2c39065becdb912057b0f18d2e077af1773217398610766e3f4caea143972ff0efd14048bab7724fa3674b0b840dbc1dc05bad83f78cf54354f194b1d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1248cadfd46aab542c554f7c28cd5054f97b2037aa3351d7796d2ad2b391f605c3e5985545897542bb368df46dd303b939b07b2dcf381392a3aa9dfe192b3494ce9e87c487cf2ca9eebeb17d3c31600f68b582dd41600aeb47932f2f3a85cd9fa964040a5f89ea2c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c438bc5555fe1e73aa7e1b728ed9815cea17353695781917b38c5fe422f1400337541dae34c0cd74efd74276bedc79086096a6dd18488aae7db7a4ea72c3cb1a38f01743128f0764933ef387f7a924797a347e362bbfba6486955dc86f249a41a78953687f1091e609;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abdd57c6aa275d7ffc3a11d2e5260dde42ee7b3ea71a0bea8e50182f3a767ed54faf008ebdc04840410a0c708145288a5a61e0129cb45c6dbd82244b50f265acdb1fc9619947933f9f4cbff3691935d5913f14f2775fdca2ae46ce9a21d47700503a99846d10440c88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a11acb76b3bfefbbe5c4cc2f7a3072c5a9903a0b7ea7c59e15034ebc1e35a0b5dc10e0b7b6b56bb73fa368200e5048215e9af1ac8fe419f339443a0f345da28e56d17feb578a85797dc2484e3d9e9ee29e57968929a323a2dfcd42ae52fb56f159b96fb87f1661772;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c7e5791a91325b804a9d20b1cdec3da7deb4998c7da8cefbbddc7aff079d7742f9d076ec6fb056636b7f1ae4de8a99aa2ba96f4567129e6d8c8c550b1e8d2d96daac1dd9f5156cc96fd9ed8b7ba68755b7bf63e0fbc393ee38530943e174e323c7c7bd781162eb6f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'habcebdf412d3329be8f52241f2b301400f13a34540699e00a2a4d7a893e2e21f7fb749714dd1ea8228b50d5ce59a922aa9d170b28c97af5b01615d6e0808a8db00337bc64b813aec54bfc68c7066748240013908c4fc817f31580df8ec8d5a3314d68876354c5831f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9d2974e73e39b76dc749a9f8898dbe103e193ed9944fdabb484c3774c3ca77439e01268fe694e1b727bb0873d8f4d7ec521a5ffaf3d809aaa7d016af71d0b4c4bd6cdef0061ea47ac27d1b59f2266bca210cb288b2e42207b6b39de6672d9ea439a673a75556a890f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf615cd865cc5cb2389326e009dd0e6fba5756fc0db939513ee5fdd012ad059d1e3583d4accbad08c2d5ec1ced0a0d78dfc656a2df2f272f51ac53a0a8a5f697ae1c2f18fb534e14ade5affd35e3c2f343848ad042139b5655809f8fcb42df1eaf0f76f869a9664fbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3279e70836a5c90143949736fd59f680f74867cc57063f111c3150eeb45cff7d28bdf058f173305e7e6515dcadef7908ae52456d0faae8d5cee11c82c98dd1cb9825b5b287a8fd7d92ff12ed8071d182d7a2f0631faed1ef9335868b1a32721b3550897c8f78a04e60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c1ad532c65d525d78f7507c5b56be148845264d0014aaf4ec87e5300ea56a9e09bfa6ee3fc7cc7297c795a79119b3f25ef5fcafcd703ffb9890cfaad025dd67fc705d9118397b258fc572dc10bfce9bfa54a6af243592f421563c40ca7b96a83479029553d21198ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11965ee8bbf2a704d3447766aee1190bdd936cb13baef662c3cb470b26b651c13dab779453a7c003707bc11dfa9d45ad58d2bf3e938997d5486b3443a1d0bfe9a92c9d7f22e7e977cd8af685476b700e39f63bc8a65e264b67f89c74e5eef226bdb102fda9791cac636;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5bd6e6881427861b313d1475c46c1b31deaed63874262dc88721fb2b538deaf38a1740fd889a219f0501de007696467fe6beef0388af642fc116703ab246983f6bd4dc37343f25e48c7c40a4a2fb1aaf01d72e8223136e37747f2cf80fff99ac7cade7db97a0a8d9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154b44d53c801076242d21e6ce10cb56a49f889fbf125a160e16392f66b1f922ce15c890e674ab8fc28d518bbfc898b8d250b5fd32f47ef7dbbd5ae7375100a91d0695844b4145f9a51ab57706ac094452232e7a07fc98004b9c761aa11ca29302fc7d5508de0dfc483;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadd40574aadf1deb5ba77c93520a10b37d0e8246d8533163a24c6ac087cbfd54f32f1ff937d581f6d4c6edf001e7eb31717635fa7c896bfd2c5b4d1c98077ec37f33f8f374465b7700c77f52cbdc51dca971ce64eee5891dbe4de88ff989ff9a12007a2abc109d445c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1656322221383be7d9c36888c6a6d613b32e27c71d71746b215a89c250e253e58d0dd930b79ab661317d64a476a211341a53c9c4265d299100f21a6e0feafb3fd260849f5fefbc95f64e55338d5402ca86db541071ede9dccd208c9e03e13f36ee775930d544981f13e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed6417268ddb17fe948570f5d44d29841098fb045c98809d3aa00121c59ea93d7b15ff475d909f0804f6be90ca19a3ab793bf2a22667da0b6015b730690724ccba12dfdae67910550d4f582a9be48fab1b74cd3db371996ded50a3b3e42aa30a781d862a47c8034a68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1e5cfa8ad8e3dd2ce87002fe2d74cef254ef1b5d1a523453a5675f803a1fc53b9575d2f87d73219f3d769008379c536a4e1274dd6702246ad280277a55e7185b8a67e1c9f16c3ab2090a45ad15d7d327786ca4a6078d1c97dcc82822d393f5e1da0d1046979c222c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c0d80815b22707c4f08b83ab84f010fa4a8d61fa6a1d027ca16d183a294c42459ce142d7494192b7cb0b978b4844f21d137e640d0533d2d8e76c2da80d25a977399ace30dd5a623e029a5995855dc092531e22d186e05c0b449c267d34c8ab276c753cf47a85c080f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bc7b4057f5ae48234ae4c41858b965642366c18aa98af77e48ac65fbae98d811a3459512dc7cf9f1701c12a5743540af2c28c642e08d9f5ea5a4e031b670786ea5eb35db59cea0b745ab321fc92cd8cc622cf21b4f0539e9d581530ecddaccad500c19b6502492cbb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13829d4b5b95896c811f33433c6c74ccdbc729e7887fdd0764fb0c3ccf68bd68158abffbcdd391709839335222e9896061c5840982f953ff935402988681aca084a2983bbcecad425e992d379fda6e0e51fb904cd8c0bcb1ff0c38ac8d868126e7ca8995f37736c5271;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bbacba9596e48b3ceb58fc18761d7e9b4bf10d49e35ccf3b3a5e4a216876107bd69c2a220d96c6a5cc959250f3a7a1838c4abede9916e91619afdf75fa1b71e7b9261bd62acbe6e78aa47b4dbf1aa27779aac0c57af7ec8bf33c70303beac66b1fbd6cbfed8ec8c4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b1c10007ba2dae4c45d132d294b4f9a9bdda6dfaab74eb884f7785e149a90c1b23601e47bb60e84393b3bc2cee595681cca55fe2434ca80aa77760b7283f5a7f2e8b8c037dbd285b6eaba6f29de08e035447e8e38e3dea1940c39ed47f78c04af7ae28c7c595ca1fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ecb55bd5e5ea050e9df4f3c6b6583b4430b15b7541598b905319a6d786f1b204943caa687b8539bccff42ba19f74ab9cba1a394ec8666ebbaead51901b7ca689601be135b9dbbc9a7cfa425b9e2f441f81ae49d2374e803dd11b9582cc2f76531b09cbecafc3e7ce3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h812a451fbd02c9c3bd7ea68243898a3e201d1b1b43d0da5f848803cc246728d1a7e83190313cf7cd3840766c0834ed766e93a90a72e4a8644fd78ad5c9475376bf5d117fb9af3268b17dcf361760216b39a0725663fa2e43cef74f71a64035647ca0a8c2d73eaca611;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdde15d09465a51a721c28a313f493b3e2110e763b973fc3863da820905795a89e33fc55332c315fc729b9eec064657712be56f96a8df5cc75307faa6651b2f20bc22753fb9ec4bb94faa19917e3437582b2c4ac92ce0e2e57a2f05e085211742b7e8ed48992f257d62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0d22424c34477a00c82c202746716267314e83ae09f9f5b4bee7bc14e80284c15bf39010b8060dedadd232fd339b5700ace6e12284c470c55548d6ca3bdd56342c075b589a5b562559215f4264fd1e27441b3924702736b3d884bae2deab8749084969885cc549cc2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90730905a28dc29a478c254e8d6a364628a366c33d8911f7509251a8bfd5153201479446a7ee8e73be8a52218d8a7724e6947b5ad16061e9873a0206a5286b1a2a92037c530bae2d29c8112b0091263be1bbe67940893db154d8374f608377cf4d5c4cd22cdae7913e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2b7ae5c02bbc2651878625198bf505c0b2af8ed114e4d1a1539d97a2cce63fa33b1c91f0bfcd9eb51efdc634912af9c979276ea29340f52e8696b07b905929bb472ab12a6e11da4e4f6ac9f6f79644b80f1ca5f336c5d0fd297cf049a6f1406c5e54791ddb550dd76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38aa15227110292de8b43175837c78831d1a39301880e263c13f3c958ab5ee04346d4a118dfa1b11044e23a527a440f8f8cf9b3899fef1c4db1d05f0073bc2e7aa3b2e425700181d10c2f1c5a75d4bcbbccc2e7d000e9e3acfc1a5e9df9505721d9447e25e43e7f080;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a7180acfea6e389592ae6258f09fa7bfae31d782ac94516101022f050fed52cc7cbeb9f3f09b58078b2a3d70c37cd043fb500714613ce631a884e418d417af6d9925d6cc6fa746e10cddc0c97e348c7ecbe44afd265e2a5e1a2bbe629ae1916c1abf809b00baaf40e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143a0658a14aa7e817434f74d4a5e5820d8e0bf697a653677950e6f512da8c00b69e19e14860db75561bc095601185b88fe06b239e2a9cf4d0bf495c3ee95a3c91d87885aab8f26b4c3a899fbf89294fa2b84d6d98b3bc5eab25d9395d602de5ffdbdf56e1eca5a8228;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118e4299da3cb4542340c81c243a4dd52256482f6ff47521696904ddecacb193eee51d286401bdb03fbe717d2426881a3d13743ec0a2ca40d5ed40281b85eec8d4290dc57e61e33f554104c455bd7cca7c1620913608c5cef055ec500d1e71d5aa936cc5cd87b0e25a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b066c1fe2d3803ce9775e7495c341176521ae7c4b8149914ccf83fdb479d2b12134f600135cec8601a5f749df988faac7a59b7ccad142e093117c799ff2823dc55fdc2832b0b4949ab540b8d34f2cc008ee14f91cf07cc5b44550ddc6e2a63fb6e536fdaabfc396c6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101e5d6a518f11f60b75ea858806c8b933ac9d80035b8d10543b94a8396c5e6546f07662e4562c37c5a5fec534bf7b34bc7841be6d480300b1784a469aa522eff3f78e4e705c8445d8e7fc6480dd6e9610162dc4d0e10fa41f3891def038e36a33b789fa65a1a71134;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121168eae9f0f43c7ae0b6d449a6d91eee38fecb08a613df9691c21ac0a54f794dd1b2cc14bfefabe3416b8cd4b155e2b5bf79dbdb908cf3371c7bfcbe367a625a976042e5d749b6fa01ce1d28069515ad5a1934efd7bdeaf6ee702c301e81ee13baa22a50c3288388b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185e03137f23b282cf7fcbda24ac8b2e5e7505778c02e4e2e26cf82a4d5733434a063e4c51d2d58bb898b2fd2d3d30cbf9ee59806e534e9d3de06a883f3bf73a8a02b1ab9313262af325ebde33bf5ecb0f89274721a249fae805462b145ead2fc1e73b0b36b59a08f47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he61ecabf8d6c6dcf1ccc89b4d17683b963995b13e2d7581bd821d0c203a3ceff981d0a78f4e3ae7644bcaf7f656959681223f1e54acc1b1827ac6cb98d7d958e8d9c1137dd12a10592227f134592558f2f6245b2931e1635dcbb49da3c20113409f6e1bfdc5418d65c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c8f53d288d93ed281b165464b60594ed32075fd1e4b5da674ff466f96880d7b3255bae2ef0bcd7e8a942428d3bc6795d0af1487e2cf97919a5d9234acfcf957159a9d44974a337ef8d140742215941df6ce8ffed54018407f6c06457a2d63a779860db2d7ab2ac1b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b50877f175b5ea1f9fc7576fbb966dca6fde036abc0c33ffecd13c8b49fc3f6cc4abbcde0974b2a6bb9a9547dcb6cdd495898ad81f6c7b0fd69bfe6a3831ea107722f6b0b07399049ee18e69889adbd6beef976d4b4726c68dbc4407460c6a61d8b7355cadd16c9d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e92fdcc5b11745e32033e8083069ea94080bfafb767eb5b8668c7668b657eae17c135aa27ca035b1348b2c22a697f945f48cf1822300fdaf0fcb92b969bb614073cc6939c99efe66cba0350fbf667333591aea7679546e32c19949163ce3b61412279a9d31a22ae04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10728f42284b56f2733365f3c3d5354bcc3ea55ea7fd0585c360aa1e945bf33670bf38fc06d3ad88698dc0bc3d1c29709de933f217939d50f5a7a61060c8a2b532d105b4b70deeca3463cab58cffb2ad70ce30d85e6103d9b86e1308badc12065f62274978e5b50ff91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e8c7dcc393848f2e69c053f8eac864dbbda2fc458b1e08fe7b63717e2c54e58ff81f20a00630ac212866931d986a9bdcd071a87335133b8625c4059ffaf0a0d702c904d7c35d3eec79f655f173cfc9319dad92d1087afc14fc4b865c93fd206fe2c6826f96cacf8c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d329ded61d63a53ec64690a5da411b2635de203db576dccb49a9d4d4537cffca9b9f33ef023f2240b29e05383635c3fbfe68286fdcc50ac27751433232720c8d1098b12449afd390715b5bbd1598d14a4fb590bd37d8ab69f959da8aa414dab4cc26f155b85c16b9cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4659e7bfc7a41eab0eede291a70e007166bfd443557e7e73eae795dec2fe6571d0a38bd63d94028919b1852fa949cbc5c133bd4049703f113b3846b5198b9beb6aa2cb6f67b19e39e670e68fc7132d73e9a95414ae0e70467220c4f5f65bcf2e5a016160a0cd0c7a6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afbb1ad6c2270c47af10794de41461f664ca878e2550bbd7926d890f83fc004f23c9e508ba4c015eea9343ae019deb0b45f6ffc31bbead81718648c042fc834956deb373f82d7fc07908fd496cec3a07a983bb31971fd852bfeb3835a35674aa235f0d21e2653f95d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167635c034038a484505e473538f9bd9d95c7a81a95614d27e67ac022b7ad7a5ae6aba30de01fb90e0732b3a714ed5af99b44144a82b30ac20759c8e111ed4122ad52bbc9bebe45ed066b34afc923ee22e50665d021edb1f68a3127d367a2398ebcb56cbca948dca795;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf03cf78d5d0840d464fc53e655ba69f21d7c139a24d5260720256a80ddad7bc59cb022f331aeb51ecb856ebaf136aba00e88081333f5009942533c4c15bfc134580751d33f838c5fda75404a2f72be59a4e9f1e725062f318596bef47deefbac66449d2118bd2c6b33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4eee1a5531b713eb473b16b5566b902171b265bb21cfec4850823180ddc4bbb9b451c3369e84c2bd3735741e8218527bee74f5af3801ad423597a245fb9aa9d9923569e66798d3d3d408e0afdce15f42a3005214f50104f743de8a847d7c6a08e443c11d5e5aba95dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36710a73daf9e71fbea749c596e61b2abaecf952c7f20435a65e6aea53d8c344a495819577f5c4cc01c6d5f15bc73044c843ba993b1781695487bec5efb1fd5b9af9f5d535fd627e1d9a953312223bf37320d8b8c8d93facc0f5a87e92098523d1cf1230fdd8e108e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a9b2df0447ae520e6d983d5e2d1d2e5690dd73097c8cb7e08fa93d7260aab36816df267c38823e2555f1146bd24f56b32978e78cacfc323ca15cc178f4fa752ff74760d60e0678fe09b718ec5874070992303690bbfef3f6744dd299fee4245d4fb3fb34f0ecb123e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef46e7c6f51f1a3c11bd9f4bb71e752a4d48cb090e5e4192d020dcd848dca5e6e2d3f42c86222e8144149dfcdfef67648c7634fd187e284fe6e472ad40b9be01985df554f4b741196dee704ea68156becaa66835fdf617cf28c8f457fcb83b94bcd7c945a5089c94a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53c0e42cc3657628a1fc41c82be527ab7063617bf28a121a76bd0a29788b1a10df3cbeb210b2c53cbf7f673f013dbdbcbe42e9e087e024ee6c117957ca68414c76fd6a9c542ac2b22f5fb4f548eee8199aad1f8a171cd22c80bc6a140b9b7da606bb2417bc63287e92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f90b74bb31788f4b96ed9b5e256cd8a86a5ca2787e25f27f5702499b311a7f3c24af404c26a1588b63e5028330ca5c51443c7f7e2dbf851c80b300e8e4e6b86791efe9bba294dc9b3e4ab356b28136b5cf6f5abb5768ef41e59e2482936af559a527632c2bb9610ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58c1d4df59018f96acd3f525aef3c272cc21dc3b820446b8f6ea69d74adf04dd11ac3f7fcbf209f00e428349033febc2af2d8d3c6e31e34dccfa8c5c4ac73168100b2289abcb8b7c14e11bbf1c03497726a1071a9540ea1ad177473dc1c05aed0470c37982524b93eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118ae159db0e075b1791542725ead4015c8a7212d9fef80e56e37f92bdccc4bb83d63f283c313e47077bf7e0d2b2ef4b58e5d3c1f3a18617a26cc2bdde8f409019c0c08e5d6b919589dc05e4684b8272a21a72052ed2b5a815cc7094f31fbd201505c1e20c2ab20046;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176a200a423e7aa133695c1a9b68ab46935954d195ab8461d2babc9cc5bbebdf38ead6b2400840c279670cd4d5abdf59b41ba340b52ee6a5895c36ffc8dbee5c91d606174f7685a9835b371b006fa989158acb6256f11fc1a18ec41b42444cb79f88d194c2d6b1b7941;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1593cf9b6eff462fe4aa1196275a365f964d861424c8306454f9225f410d2f824bfc8b0c645891876c13f29ab4e054f544132adced43db6e2fcb2db8f9af984d6967ecd58dcdae7cac4ada75ef228e5a2ad00a86bca04d44c985f820e2f4788153f71b2181b475cb1f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1511ad31548a5487d3a4999317bbffc3b044265167dfd6d35542d571d7b2d8c94575ab43cea9952299ccb61a614bfee8cabdf5d4b4af107a03650113e70c78c19430880504d29ab6e0951b4d91da7412a60d56f81c7f5f89c43f0b743501db344ca83df8db50c6334c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1450d8bf01cbf170a421f731aa09256a9321a751fe171c5fd52874fa6aa5f0b872b708d1aae47b1c2ec816f843c986d03d978fc83621c6abba9b46f68a083f0d619ddc36067b6e3f0a38f412504d69f193fb13fc831961e08a98c09c0bfa05f9995d7114d2e732768bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1947e9698e6245365e887c7e3e503597382420c2f9eb0ac84462baccc1ebe6aeed2d21ae43a23ce6e10cd05ceb5424a710d31349e5b4181b17742eed10d2eef868461881b685800fc9661f15bd5217e19809e663e741fe84ffc23e8fc2d5cc6bbb51dcc8e8e49766e45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9a638e01d036688c6759d19375ef78d89e8367ef6e188f600766f15bb499b6b9ac3f2461e56bfb993a0087ad587b4b682e5c051652ae3dc300dbaf63c62e942aad56dafdf5b395ef03aaedafd901c2298cd4cde5d7a8f2bb5c7ae8360af81e1260f1419c47765a25a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8626e1f1d90e215e63ebe13188dbee2837a64925bc8b701aef900b75a5fa10aba3df5f21f57b15b5e82b1aadeb0cc03f6fce47582a559eabb24f670f9fb6b48824145265f5c2377894606a9fb6f747994bd985757aa580c711d49dab3c03faba1d68c1576734b7459f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140243c661f6d2dea15ce210823cc956c44be37360cba0b9c2206b3cd387eb16856ab09a014513f37e710b35d536c3cd0ddb239aea8082ac99d42676ad29bc0cbcb5565e8794e9b6484e6f5430156aa7bb1bbf6a9d22ba6b780de3b3113d3c2059b4e7f37e6044d2046;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4955e81fe46984849cba70ef59bd7f03cc05cb679553195b67ab28405a47999388769481869cde1288524e80fdcf9b6da4113191495ca269dd8d41d83e86fc835443f87a4d411a887a8882198ca1a30ae6a338614296889dd8af383895f47cd9dda5927521b3fe6d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf373811be9449a2aee317a7ca1a6728009b11fdb1791735c994f36244af7c78f2259714220ce3262ac25346c60ad21448fae32721ea3624e39a3f0ad879e4fa67f8b21ce5eefceeb0845e4f50cc3b507977ffd3a19d532d50cfd6a91baab47baebc0472483c9a60820;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33f15c59b6ed910ce9db1f47589ef3ea7a316a2412a36edac48b2c5eacebc76c8153d5b9a703520b410c45c18f1bb7df01a2391a759571e295cb073f127ef55e92324d1ae851b13a2df0c0dfc0c1967a07c14b62aaa0a9d84ef9317ac345b53790e4f85423ec3059ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112fd7063d3f8898c112c5decdc50904e968281c206a5e33c5db9336a31134122a26ba5d09ed22c3e0c03f768ca099783c36d53e6f5889961a5fb8edaf83d23987fb9b2d4419dc671d0401cbf43b64b0635607034c373219f3feae93226215f88481df4ab768bc779e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55504923cd1a4666c3ec5375014fdc8f93488e4511c53218bb6fe9f6499bb5331a2f95fffb44447fab9f9c7bc4213eea0bd1b4d56474aacea007c4d74d23fea5a7ddf028fe4e0a260475212b38c003be7da82b976f541d9d94e85204bb368863e8c56d3584c49790ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1985c7d472a7f015dec03c3bd5a1cfa8ce3f3fb91ddcb210cf35e56aee9b43de57cba8c42ca1eaf6e131d05fe9377ebbeb41fe66cdbe2f2e9533b1fb611a8a950580daefa6f206817d15404280ed32bf2c9dea248966f9a740d01a5dd5c73df227fee72bafc76e7d741;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6921d659a8dab98ffd529e32831f776a4a0840e39d159053e59b6481455647db7a64da0bb6197d4fa2626b8b689b7c2a7390821d9cf46bde1ab2ed52596a2c346d22edff25c57ff716843f2a350b65fc3636b718da214077b3699cc422004fedf0e55f59d85fce2a74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1863ca15d3046b3e31efaa4ac94e80c4649803008c789b70874b7a1f94fd1f432b9670dd997cb36fc73caff5fefa9127041b703968b768206d001eb9529b78e126fb7447e8912a8e0bbbd6fa02db73bdbcf5efe29c37a457227aa0d835ec3dedbc038cb0d29bb8ea444;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196a7c910a26b0c4621615b7bf38c8fe81000892d3564d3c63f73e0593b9bbbf2d95cd00812eec8f1e4860420ebf472faab753c3cbac339a9f0ec52944165e6e9b5245b4bbc1c0738879b1d0531ed507bc2eebcad981fe1127c081d6ba44ee31f7dc1b8823cab68c1ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e57bd90ab4deefa29db052b89a88b09ecb24caa6e3c58666e35ce1e2015470c64eb34d3ab8dc93b0aa0fdd6aa0339e2844fd5c7972fc9219e1cb597be43d951ce347ec297bfe3c8fc8f319f0ae531dac1ab58c7134b18086c79e7979e0072c3badc750bcfb0deaec46;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19adca3286c0c96aa7423dae335d930ed236adadaaed64847807f010e81b0bbd629c2d1ec9b9c3337f6d2d5f5da20b4afb73e73e0dd50e613c715fbdd862e89edc102009d5c97dac1542a25c245a02ee8419aa02bd9eece4d122454af669ac1fb4faa70e477e0422620;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf90caca5246089b6242b28219a87c19a6be72c8f0ae04efddaf84433c41a24adcb82723ada59745e0fbfc4894c3ce6c89e449120a7928b294a3035f6a7d096ada32bd14f602237d0db416a1a5800cb873b710dc4cc31a84ec719c660079e3df7caea5e0edbc161dc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73e26d45c89cb372aec5a35d554e1c12c27aa4d37df53cc09e53f9c16e6472b3395e481d291862bb8eb67520fd73bd85484d5692d52b5674142067a8b8f2e053a7455395fab94d0dd883977488fc87e7badeb4661f9fbbe84ce43e38e170e5548eef77c810cd4b8824;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7d5f2d2cd1d6e3690a4f1a886cd2d53065ff359e27ab0c675f77148073758270308b3b78cc85f67451df290ddf4af5f95c1c7b3a3b7dc891a2c6a02f932c210b58b94df4d07fef0a58dee418adc84a15d80055abe476f5924896e28e47a367a8417fb1edfe0612a65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddbc19a87923c2fc849e558e2c6e7247007bf70e6bf6a24e48dbb1355fc6b59b3c8d64dd7f6e8500d2118cecb53976efe094b38a3b5917de8cadab0eb81e9e393e6c29c5ea66ff50dfdf3d29c128ccb1b042c090df44bdd3268acbdca13b33b9b058562c1318b4b21b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a222afb88dc51cc1832c458e0ed5b5f1379dc46066b6a83b7ff328417220f9df18596c3c22ef8d91bd7b6019ab183cc78dc4e1778cc19a736d88df4474846f51132597c820b93aa9917a5963a392728d19b0e05da82c38ab42c46651ec446461dbbebc6a9058bdae72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127686a6c2c8def1a128a6ec1dd47f16daa942138c15d2b216be21968caffc54845974115be4b069cef23fca181d2cd78d25999c02c3509f496ab5607527a5f3f3d81e683ec6910c308aeb33f5a33548951e00d84ed25929f39ec782db9216b5abed3eb2e4d53640e63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c8c4d1fb0a45040118e958d083fddfead56793bf2f7f2a4126231b0efa785932049676edc1c6aba55b363df7ff574a1aa84350894a33a788b851ebc9ec8c0144ebaf3fce98bb39ceb67caf4c7c085e3d0619bce98b8de8e937fc7fffa5816ffe3581d4aa24fbf37e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e4311ec52d4ad50eef6bd7ee50b9ce4c527f9596fd0eff1a1da23f0fd1aa0008b16cab7f7e8448601fd6213325d52397a172fe3a53eb924551251d625daf2148d347bae4e4300590cea28a33451b98e61537766edaa14af9bad7b04a7dc6a43b6c9a6ccde930cbd3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa89f5427620298e78319374cbae19ad2a167dcccdfdfb1b978de538177cf4fa021951ca1dd97186168e05e998bc1a1853f1f0bee304a920d17fb861ee7f7e11fb9c073b65a41f7039c10f9d0e91038a09dad453759086092630788fd3a620c290f7ce90b4a5232c56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162c86ef639c83e2eb3d616144945b6760d5274e82c8878518090e0dcf02267879d3f5cafdf7989319dff7bd9e123ad97f3e34c312514064c7397d56fbbd298cd8f24674246013bc479b2610c63a40705b69e8fdb35928ffc09d60e8489e4384a2379d6c11555e0b4ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a175001bf5d3ce0d11b3cfb416078117e5574fe3ab938f85a817ae8cabede33fb0c04911bff2a01e3197814b16041d976c0a8eaec326b9e7ab6a9ded4fc4b7bf1c717ae5774093481aefd2f1b7b14177f05b572861b9d072d163148beb3e74f02dba2eca2da328f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c095a18b7ef674526c64adbc5fa97c967e7de4b783ca6bcb39c4b4dc6e76a290594027c487c9116a359014570fe07d12f98beeff376c0cb8e1c72ddd0e2c8dec429adf06e341f7d4096e13a3adea990aeeae89258e1b5f5168daf7f08f5c1d23d1a2f83a05f970199;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec2cb5fd22662690086ac0bf665358a982ff80ad63243f1ee38863b707e7adf078923e5dcd1cb7ac53cb3fc8e3b9d49ef3dd95780cebabef86c1126317427bf58eb0a5edbaf972214cec84add8572c20ea4bcbb5b3b2447dd3ec54def94f18acdd17666f90df538561;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc5c5e89bd12c8348f467f4433c6315614afccefe5d4934df43c579d955c343e2aee7494045a812be6bbf503ca5ddb6a5fb59c3400830f61c2085c32748cee41fbd6d9e8474f8c418a540f2fc79ee94453404fbe6aa3cca6ac2315e6754d09961c666e0cb14bb0a29f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c24cfa2bafe25b32159c5898c81f01da74f4a56f2586e891165f06da05cf148f6c2511b449cd8b398823edaf593099df8d3165bcfb50c99ae780b7126bd6a863566272f557bf78122caf9fa19079f04bd9f35bd02b519f2fd7c5db42e91026fdeb8e1ed3f72be32e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbedebd46e4bb3fe2c82ed97845338cd60243747cb4a1f810270c77cacf6fc438e4a2bb3c5654a2a0166205bd02b4c810f31764c4f351d1b116bf1ea8a912374719c8555ccc9a1ac136dda4b29376a9fd8762c3c227b9d4a5707f7ccad53ed9962b22ff06fe1734ea49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae85083e5876ee83830fe7f05032c770588e938c6be6e851675d07cba690e80b22957e4721cb5924a131e710f3193834961ed735f644e4c9030daa8acebd6102e1d48ca8e2224c6186bff85e2d6e44c208f66e9138afbcc3c19ecfc3628c9f32750368534a35f7364c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b85b222d157bb31b50308341f48201445747857187d7b47ae5c6baadc6cc64c4fb9140851c77bc02a8d4452598d5de9113c8d46e84500135f8f2ae40aa68c24b4624ce6a2215a349461cb55e65fa2c198c0e9e7a29522b6f02a86fdb49ca255ee4e156710c421bf91c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a0d5b30e99e757ad797368ccea9b4aa4460dfb1d0d6b9f0375e5dac2aed2e5a3eace2777b87105e5d9bc3e236ccf7fc4e146994f41189d88cd17882697934c4b4fe836f991d9e82e205e0576297c73b3bdccf23e0de534237a8fdcae4752aa7eadb55f1a5238517c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3be5984db217146b16d602f313c3085ad2272435c5c49bae749e6600c7f9c1db8dec7d5ee7f2e41121639f17f5b080541721e09a5b728bfb4c193baf2090ed82bdab130cee37878e0e3383d0fbdf0b7a46f4cd2053d2877d40c65aad707835c79c0f56a21b05a55d1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h232c87edbcdeb8611ff876e66d5341da4e49264be34e7b1210b5b0e7b5ed9da21cdceeff462999923cfdbb5a6e98dab12a2046e1a953802bcdab1c0f66180593cf44ac2d256424e58889f42c8e36c11ba74045c77faef086f2b0120fa57cc7410d2fb3866683e3a64a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3afa6c8da989ddef10a9188a42309c24deb22eb995a4cccfe4ce6d04ca9787f2149bd540c13f1a37c174b92dc6bb23673ed0809eba6489733272f461f4087e0810b11999a1e429650722dc9228d3b8d95610f836fc5811b991110ca71b638d1d09a0b8dbf43c2125e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h519a450a9604109914e5f9142e6bf5d126b0a8ff886cd13a4b359f01a3dc9df3cef505187b311610f82ea6b38edb73190af035c8793a95868b10f67fd446d052f479e97c534bc8599c31039a5fc88c92210062787be436f39ad2eb9f624489c32a2895f49c6cb08b4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1966822ca3c5d5fda0967c71c25dfd1efc9d2917a5eb86f61041ff0cff4f0e75d77ee85e095b80156a937442491fb502f7f5f0b095d0717a94db0d8985e25f14a8b9f376e9623f9badf2d3f6d0e7f849414b4fc417e17b6371138f284cbe78a21e9ce4732463a7462e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfecddd6a245fcdd74230202e0052b402035f8fedbedd4d5b9798334624637dddcc59f997bc405f2b6f35764dac0d01f04d218643842d00a888d50a3645e68fd0150364ad5f178dc0ee5a95145a310a08bc5b9f066e522f31f313cde9465295eba96260b3efb07f10e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179ed4a29c014d896f2d57a0ee48f8458a835e092c1bd9c65d913ec9811661fde7c787eaa676534b262751e7958e5d9075e31be47077bcf6a69a0283fed03d25ab509d6219de905f30b455774268be5e58127073e3b8d6187476ec0ecc3a27acc30a96949d57de327d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c0753e2eeb4ddc05a87774078b6c6164386372fed0f314e91c31f9dad26d38fdbb34be8a73ccb87afbbe807ac44056296f83cf2149f46bc2b2e04b0b24c0d98d36f18e5dfd117355c0f65e02feb407ccb6c32cb8a9fecb3dec04b896c904add1d0eea0c5f12e6e1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83aebda18f2623a1974c8dcbf1d913c36595c5c63e3550c5e0f81d7186124084658882e18aee080adde884e0c79d9c91b634f32827316ffee16a5b82cf4f8d482b12334e739a634cd47570fb19614f716b54a297da419a86c78ed07e31b4a605e25af611174c9edf13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef15d78e2cbed6ad63ad09f7e2a93a8b6ca2e56694e6116f7f48a4feca83677198c853b7188796fdf66b541e9c34658d5222539a1e929a3d14d85261c3e4731dbdabb6f5fb194933f9e8a804bf5ac43e09890737ba946a994122f0f86106ded62c2c96738cac78a185;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1292bf327999650ca93bda94ffab601b4f7d8e0216d2ae4599a0894e1f8e09d84b365c429c44e27e872c839f493c8918c716aeb20074aee8d895a8b44236c88db845b345be0fe5513a58ba06b945d0aee691006591a254698768b6bef8f7a564063d59a4e54ecbe0e2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e257733db780381370c0e6da02fff282e1a9fa447b82c33eb5c14f278bfc710dc01acb933f31973f8af1b73b1caea8898b3176df15a5ab8a47b5a8baa9611dd3d6b40c17089889e8cf3b5dac7a9b73e2e6939213e1885059243693194b31774f2f86e072913446d3f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c130cb0c98a260d1ec236a40cd612c4dfa25a9ca9543b52abbe65d19a7d898f320becf9a03d0d54883507006d607f3f35321fadc7a585f5bd7a2ac504998620559786550558a5d49a9799b6d4f05dee6e6b78c875945798f1021c25f727906ec1a6fbc68ba79449fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h279d4cb40d98fd191bcc00db8e6d39ac7abde1e8fd43c6c4bbd78e27e95c2b30d19e9194e4cbeaa72b6403415eb86be8725f22e311e3a21be8426ae94862b592603fb8f119b9573866461b1176c775161fc6de00d7d0d0b362147ffbde2cbe0771ba16ce021649d8d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h778450a633d48756389c43560d5933d48be45fa925db52f9fe93d3d959c05c7a6fc5f49c3d5d4fafa87b49e033d6c4c9733a6f8a7ec06ec2e58e551f1803f3f24170512a54c887fcb789d4037e24956a371e591c9868fd46a08b76348222a2938ba0a2df47a38d02c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33a24b2b43ee33d6ac3c094590adbc73a20015d97b3436108e8c23ecb0726ba65c2ee10eecf8e7066c0fd1a01af4edac2e8fae9850a80d4c83eeebc41fd958ba1ca8b96b62325a4f01401e508d607829f0bdbc0e444058c26cfcfba9c7798b2233d6c3d154ceaf54f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1202d5a6bdffbd25c9165286e7f769d671ba16154ab125ac4a90e4713614eee674100dbb1df674b19f5e37fa4d5922d28bac8be14e9b30fdb0305ba46d8becace97a6b449eb578255a154305007e6d2a58fa50e134dc7134d6e0d993c8e3820f04fe857ff4e9f4ebcec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f62ec31e80e3cc7fb9800c460cc068ac33a9089e2c19b52b264e6b10e48c60a3509d3e0423b81916f16cc06a3f0f9e4b9e2d4b37995b81e16f6368a129042fed722dcfa15f0880750ff444becf9ae8a1e8a63ec168983a0ea921ecf763816744f5abbbfcf317b4c386;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf03abca8b74c323e7dfe19b277dceef78e2556248cc878b87389518ab871d2e058b688c85a74ce33891e2b117312253f9166350bd2a51809640fd7442d5c8a33573981bb86c77903426af271369a6adddc967303320d063149893edf6c6ff4eac2d358f50e8aafe8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12df062ac2d663c58ace284800c23fbf9d9513d3e20c6a2b4a03a3a3050185f4b71bd0285649d33fb984c06b1df26871d028da8928af4448c9c84e83f896f2a1be2ee02f7fe2fb57ddd1ced3a4311cf5f9c73e426a9cb09354f23cbbc52d5301a34493f688b68817ea2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125b05e6e732e08927df9c5930c67de3bc8bb72ec3b6354308d0c68557edf9a0571e5a825f008e7e349743d3cd789f6f8762d80342d8c1f2406be4ad790023eae57bb754979d04e2d86b739a0688497a8f9d188a7fbaa97bafa43cfb2b51bf8adcc1edd9716a179fde1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1001194fc20bb7399465ede568c95a2f3315e4322a63736ab0860336810edeb00b99aa50f7b0a61311f8aadd2dbac8eb6e289a934610019faae19af642688a079ef2836b67055446b6d47988117d9148ad69a9b92aebb920a0df0b7e334939d8018e9126ca2c3c60126;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14283b9355fb619a1872289f57fca59bc797a0f824c0778daa870704b11abc42c252e39a6e57f0f13f55a77fd1d875e316b1b29759ea07ba2199857368aa01cea3f2be6483be5f5ac1e9430f15bcf2daa8fd9887ad372ba5cfb6af8851f273e6e2476c37914d60df024;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf988cc6357931103be603ade48d16c8504002509a4f1fb372d82d5df252d0bfddb81861768dcf62310650470e07e9afa86795cec0f9ff15c574c95c0557cbe5017808583713601d03671992540d154073cbcf89ac3e9804420a84f4d1edf857288055e1e77a2aab8c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30af4289b73685b1cd5f20e029bda6d475f809d68b9fdca95047596e98b22492e935e8fe7a3d3b9375c41272ac3378d6c426be889c6d35a41f47c9f4fcbf3f328688126d15bc06e9d545dc9b00f8f49bad6637e9485330680f7970441bda471f355e315773cf6348ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148bda1925fbb8cd437d48b1bf8fa67066a7c3834c64399f6c54c8c30fbfe3b4b1b35bf45e32a010b319211a10158493d71adba4fa7e58e4e1055203c07576d665f0dec2eb2283edce2d6c7d996426566349725128a4c651fb459d3ad1abe29f2e798e0f4c23a301758;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48e61259a84319e6d75947ec089730a9b49c50b5df92ac931acf3b2a63e70e1deb9d499bbe20d0729d3f15322566a58bb85d1d5bde012edfd60e28913c68958e81a5684cbbfb706ac0a796effe7fce5d119cce613bc723c0c86529be93c71a97fff9a21b3766b0722f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd7f01d94855d0faa085c6d847e9b488454db879dd258f57e557f7eaeb0dfae60d57f5d8d938c16d232695dc5d3d43dea0e61793548ef67b76c34a66c31bd1fd0ff310f20b287e3172fe840a9869565ef5e84fb64ecc57e9cf074624f0820a2358a75f9e31380975f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1357f71451871702852b16b87097b32ac026e9572a78dd3d3f68082dbf77570eacf1448d23d7462d7f991a41850e16003d721d780de1dc34ace66bd7a94e70ec36ab7fb791a98783be7fe6c9a5fa53ab4a8d39afc01a3d1c3011685a5724d3b584ce94cc2372c541acf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcfc91d3c9a52bfe9ef26b085eb8a0e102350277b2ac6b83be42288ed1a1339099db44193bcb641de61e228580db4237b92edbd6e289513ad27574d89f27637e331b5572b5226e2c53341e5e853d958ae7061ad65bdd1c29503b736d4743d4ce05482280671f6e2755;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5ab0f805782e3309a4463cf7a51cf86a2c5c09b402e0e5023fccca002449c74b152a40bf83e9fb1f636dd3696308df5ef607fce002bbe2781bcb6117326206f3136c937a89d87a408da027002cf437550b71a29401b4d05b87c2e8576abd63bb285ba69e0e62817fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha83f99660233a5f5ef4ed5514974e1ed11d4c30164c959f0ebee4eebd392c125024096bd221b0c8c94c29e16b7d56f589e6647d9ce86eaa6c3621974d1a395e964b96efb717355cce4c9590c524450d880e1df2933fa83a8727cff8961156930a504e25a7d8b3ed22d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1873f0e5cde66d9c4a757a8a01c48ea674479d1cf1d9434525c0b29d79aeb145bb93e29ab35d753c112c664099b5fda47e2e17eaa3830a37df99fb9f2b75cb5ec4c6e24c47f800c80d0cad1e8dabd51311314e5f17e5081a059f1c75aed71d121a2962bef93101f3e5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea24d050fd20ab2c73353f84e2fd0dc0643d6a5b4c5a244ef2adf2e2f56d0a44cfc87a059bc74b49ef4d50ffafed9bc7a094db966a265fc4ded2979227efa5c984e562b9c3ca413f478876fb37cc7a920935ff3fc423b2b3eebd5cbbdd4392416cd3edd6f22418bf71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha40e3e59ae5ba2404e6798516c7f852f27cac5e4ad436995ca80f326137b2694d33242c99254fb29800a2023c785b22921211d7c67932db48703f468280c761b9eeff7acca486955b1b3d84847a849b1372a57c857c538a556c466bfe00f6d424286c4b15a52de878d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8157a8966ac3d5e0ba0ad71c77d222628200ed0bd2fd7e52e0f8d8176d21b5a1934b47e0247f881c72c037d9d3f9122e72b2aa03bac6f64db4c0a90fc68cf46e61a5acc58c64ea13aaf1378d1a894866f9fdfcd942aec01ffa4afc7ad82439d64e78510e24f301ec6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2e52f41224883d733a81d069370b90573056cd05401d528e30f2b02738bdf4cd0ea77ee2f55080098c58496a1dd332641411ee34739ce8760f409f66b52af388fb76183fc46b3f1beb98e5dde3cf9177ce55ef534bf1f9ab4fa2fad81361f76465bf920e4df43019f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32fc3e9c2031a082140a4a9327e2c5787f67147aab10768f49b82ed39cd5a2fecfe2f0e29d7866a42fbdea00c8b922d83b889f71df9e1a8111a0f3cc7fed33662a61a8ddab75ae4e3a19afb168d1d4e199a5b85d3cdf57e99f3a856296a844445b75b619c05d472647;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1942731c4d41c051ae978e1337194e2f2cc059b0aa3043e5d59e288839cfb4c87e03ac8987b84a723073a73090599e4f6774aa6aade87b0e236c4f937e7ac6000a7280ddd7082ff049b6683dcd5dae1cbe3040756afb8dab8d24dbcb74b638cd680dafaba08d637334c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd43199e2af4134cd3f359de70acd191c6031bc4fa46d8e29fcb942d6467ed8ef351b0ecebe63643a3435e76d50a0dc9fb8952b1327a5f96137aa8fbe3ac8bd334e9fc7e29da7320771d60af8596a566f3892b797730208aa6966df8ee3f61efc571548bcf968769464;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3d9cda79087e92fe135816f365b87cbe6dba651e6e5980ac3c1ae3ce85ef0cf0c3df721b96975d03047e1d8a9d47408fbb39b94739b0fc639ee5db9717cd706404892f0bfcd951cd133045a2cc26a8d0f7cd91abb7ed539a1670e413464d8cb512f874d3a112ca8e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ed20649ac29eb5b876ea900e610e164ed43d33940983a350ee03c43eb62da3c5a709a6bc73e7ae5f0a3fbcf9e563144dfe64fbf21aebf7cc97979f520b3c88cfe9c6cb5eceea710b7f0cf2090557e1920ae27cc9ff808ee5a85f4659edff894634b9b5ddc1e0239ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183826d4a96fbcfbd5fde69cb6ea9d5f7612d33fb438cbc0ab7b9164a575c5ed0ff3917cca13db49c9d66911201824c73580c0feea2c56c95769d9fe12d6eb8fdc3c3e8261eafbcf19ea021c8e215b4518e6ea91f43485f6aba70619a33911515e7b12916bf623c8679;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18abb7907eb94f86f54107e9bb8a34c6c16b8dbf43b3107811a4df6c759745968cf584c782a733c609eb9d3f615704a001561d544dc3283bff4e12d6b1d2e8c503746692d22c8c16f32e0c79dc82834b4504f5ab2b65ddb9266f1e8d5949a5410fa81d0fe7074f9a654;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16633785f077496aad18230acefbc4278c56437f2b7831869c89c007c547b4f47c1710ee8df3ccf690c0d050970d222f34340237a82a71c816deed914356c8f9787c017c85080b9839396a975a5c9ffbcd2cade8d8c9c514f39b0a04aaede28ac5b8d80195e2fb915dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1a79f7c71706be602b57f417e92769c22246003c31c8e0110e9e1e62ea8da50038ba89abba46dfb6b379e6fafc443acd58835a0bacb4a71695e0c8ff6d16d895081b1d03740b5c787ffd130c086192ce8832af6001cfd3260227e77b3f91fbae3ca4afb05430db80c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1267931987169836638d0acd1d959aa338d7c733d7b58856703b33073a312e1800eca08d86f5c33e5a4b0dbc8eaa66bad183652d5001ff986210f4d1c8bc08587338f95474b025cc286df3334387b9c2a909f47d8a6441b74b57ba4914c9f9f9047a8cfc1fe2fe7e4c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7de54d23910d89c56c1b3b3425308971f9e19cfc71ae7861ca7f75dcd668b6fe8a901229433b286fb2b92278ecf8fce5b8c88844ebfcbe619632ba6ac0dd55ef1ec9fa5bc0a1fa058bbf95394963f68bd69de455c9bd3727b2304212cb8ea262bc1725666445d6f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h722a2e9fcdcb02c4b7e339f236159ebe66e528e9234a15a4b76895cd59a7bc11330b9fe9a3263e314200ca67d4bbcd92579fad3f2bd6ccca606c0ded562092a60c0b62d7c392a9b1abf794b70bb02273831ac1e1dccaad020faa0c0c236f0932203f19440b9e188b0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf909e9308c6aeffc59c08a7362d1afafc27317b88b4d2ac8aa8af6657dba1bd8b3b962857eb5b796fa3bf2ca76daf54eaca50c7511698b6743812a30ad63d4b2e12e41b9cc3e295c4ad0a507d008acaef0f97522c7522448a39d46cb15a61ff8dca5006b30c143c6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ded79e5b1ee67a391c424d3efe367f4f6a92de3f71c5e6bb9c08460d8216933f7c4c9f2332351ccd7e798d72daba709ee6604d3e842c49854406ac30efce7d9966fc3e70497a9684dd03fb8a10449766c28cbc0bc80ed67ec1dbe87a1c33cfde9137b2768a4875921;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e24656a69a3e001cd0479028e5edfd8c30877b40d1c286ff2e47e80198eb19d457f22beba62437b58f160355307ec76d1f5f9550c06742f4d8fd89992df81442247b0eb6ca48041314e35305e9bd99d3598f86207e328b12a1001058d4cad6e4a409aca1e8b05b5e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd5c9538a0fb385ac36abb1dd9706ff272e4a27295cefd5f957ab989c759209b178b2343d35cc2ac28627bd453f423fa1e68df5a527f68473cef0874684c403b255f664d2ab224f39652b41be758fa155c426c3a38acb0b75057cba2f4a4fb693ac1c3ccf2c36a35af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ad4dc23f86fe709048af9c5e6993037d0cecd69e9f9127d19edeff11172af19292d04a9e8b58a065e63d53ba561a24c8ccce60518ee6f3739300123b1c169f44d1fabcacbf9f448edeaabc462fbea5a85526ba41f132e3ac3ece77941d9bd24c50881f3311e8b07e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce0730a309cc6cb7dc353e68c2da77c543589d71befee13f6035c998ea63d5d2bf9a6c53951f5dcdc5f007be06909c043b7f00a546c957838d2bc6851aca8d5610ed0c3cbb793319573230ac300dc69311e21cb1b4e562f1e8197ff6d02e080a08c2b9952f7a54d5b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ead60bf926e350604c14ed0e520f305bedb0ffbb182e29becbf1a81af47e0fa27c2a7350e50ef9874e118f59fe87e2943b7efb76c6f8bda7899dcf1db30be703086ceaa53ea87ee25c4b2f64c64afe3e281409ea8ef5aa6d3ef5fa99d927dd45695011649c455f275;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a405bf57669e8fa18d84a636048352a5363621f17057ebdfe3076646ac696ca603c29ad9ea45ec812024408cec11175466d19bac8be089e5d395708c8dc4a57d0ffc563f9d3b9e4374ff8036b703fc881785b2c6d18ea5527c83414fd4ed188c3b40f7e8b5a1b046;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c334b52f1a170c23d102cc80ceff59c058e56b49273a73c10c1b1f15f6e9b87ecb6b567755f96855ca20614a2640d67b62ce03f454bdebeb7c91c1253ce2b9dd9d40166a8ceae2840de5f96b4ee924b059a3b45ed68d545906087b46e7d5290876279b817ace6597f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f589b86db21c5816b92f3bf82131d2157c21fe3eda2bda0f6a8982e03b84c789cc72f83cf29b8c80845c8d0147c978e3caaa2719a405183781f929ab4fcc28b0d18416bfde31519d8f66c9bf317eec6c31dba4ffbc95d390a3d3678d6bf9f95d13c98ad033d44edb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he72b0ef3a3d97db1191a74327805a85918c0f2e231aded05ed74d86bc60a1b7a55bd42f5438b7e89f7368e7973444fcab5b1bc36c622cd276fde01f2e055d290456d1f6e6b6d8662bccd6ffb2982604ea920a838129a3fd8772335cb34350e33028644bce86222f252;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c50fbe8c9c73834c7f342ca4ca7e361357624074beb5140cccc3d340758f589f715336c7252d1b088e5cd87129ac27813e5c2b89023e156853be4968472a16e623406adfcf837751f0f66e1b108183abea6ee57be14bee8f65fb73db5e95d61b6ff8dabaf695320662;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e6ef897e97e8fda38fd9ad3e9f2286dc32acf1aad910da7bdba16c02392baa8e346aee02e37dcdc981e1b0b9efe867876eb603ab6fd7542dd584b9979bf1971e06a14ba1dfcaca5124a542d49f5b750f7eae58756992d3a19f181a1b502e4bad74f088ee6c3ac0e88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8c3a084bab60cb7d12a5afb3abaed5ebaae7bb9d3fbfc3a98856e28271d8bc25c8ed897e34fb18208df30387d3a8937c1ca9dae310713f65698cd2a607387b8eb4f1e3d39acdb59fc03943ee1dccd1b4c50ff75f9569347aeeabefeac9f6cceb1a02867eee409c395;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc76f7d79d97a64dbd37a54f0a4d471b60a1073237c789a2c661aa5e6047eca64af6a73b31a81397eff33c432ee29c99b83a931ab39c681f0185077a409ae74382ad452338965b35153b0c692a740d4aa1c36579566cb1c24c9067def9072f1df8ca9571f2db4b58c6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34d309249db29b2ffd664ef98d46dcc5b86edaba0468ded1903bd70c624a9362daa2d5627e601ffd33608096e613b3d76c63040c3fd72578fe4772b8a223af7521862f3d675e6d2d946f9ef1e31b8126df455245bcd5491259b92ebe362b00ef171154f63ab18f9a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76f530c9d879404876e8279c40aa4e3b2aa33b916a894618c51f71092c47c88f95907bf4c1893a0e9d2c6966339324b125893e3092337747c8f0a73b1f68cbf7a0c61d61910953ec25e5a4c4a5aaf9de43fe836b2d819b972bcaee9f14b80ebc9a088eb7eec5ed3178;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16cdb67a29874d97293feeb70dedd1954fbdf42298985547f7e8764db0386e1ac63d0d5e4f3510183a067cfeda53b4e11f827314df3ddfdfa16c642973a477220a76addd11251993a977c1c00cc655204cf47f3207172d5b3e65e98b508e0d56d971bee6f712a074704;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123caaf784e13631421c36130c66c89a31dce7f3959b38ef7b8b32bf04e8c4cfc9e5fa00e1d94b451e5764033596a81724f2145fe0e8e1ad2fb962475ab766a426be005e4c78eae475a3021bd7c0e080bbf1ce782c9eb6ff047e7348669127bba8d0a8da1cbcb3d5962;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1deb1247b6f828a47abefc2c6d536f4612ead4eb2c569eec61da1eb25e7392e398f5b950158f73bbd8f4554fc0d2fc33731754358737ff11ce7babc041ae45100dbad1ebfb56e70930c8fb8eaf16661f5aee3e756b599f347a13be14284f48d7f32227a18c25828c7cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1521a98d251813858ce537de43838f4a968524f24595d831c070c6f6b23d90536cd9ec29103f53cd6f117be2faf35f15448b6ea57a6c2db9801dcda914e2457fd5551e9fd8cc57125f0c1b8269f18c22115cb75cc3f5b621b3bfc9b9c8cd0eca481f90538bfa2735968;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b440c66cde9cec02c977cb0bdbe4ca3c0e52caf13e304a609a29776c92f25cc44c04734a7f5123ea89f4080d84fbe5bc7355bd0f2a4d20bb6bb33742f62fc0569f86ac492bb1812578a409f8ba3812031206714f542943704b42b6dbfa48d447ae5468d6c3fe9b34c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101c0d8af02a9144dfb82025cdc1e2a514cedb0f40c9c15136effafc918f0b95b561550f4b5239340eceec520b2790ef912fc25a54abe3a315a501cb6340b62e9042029a96773537b66955d9bc9217be8bd26d2816e0de0d6eecbdfa2aa65858c9b37fc604aefb1a830;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b15926a7475f58b9abf5112b685e7c1f5194d58517c9a0ee8e61d3fff01054955d8b7a4b1d46b97ddd26a782d8e3f31b0b02e689cbe9323db23d0eccb600b21ca87c961e12aeebf98c94e92bf00777744af252c5a09769cdd1a30b245f28a25098f09f84424c14bee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66114cc990522c2920848056caec8334a393f16c0f2612c16e7d729d7768a0ba184012f32ce60ba11417a0561673fcb39f6717f0a36d1578142c4e765f14129cfaf6abba9168f960b805583d70a593a037ad25ad571385f788ca33e93be3b4aa701bb1b647a9a7d8db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81a4a7a943c889d6688c40f1fe8af1c58e25e6aa9bf378d71685a32656110bcc3ca14f2a8ffd912349a3a0bb6870f77ee266d8e3997ed8b9f4d2241a92698cffee924b0e74bdbd6f828f2db711a9d05bae77e60c10ad65e22208f0fdfd5fbe361ff28cf8d0cb4de958;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b83808eef221687516d7973f772986deadbd8040ac6b34b55c4d2accfaf7149ce5db9ef0938342e1b6616cf34caa74a1f2937606683a71c43d5210c8b441734fa78330c7831c7bcfad5ae5911fc5bd3eae1d0bae8eb2a67e1ba6574855a27b3a55705484bc6f280ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ca30e6bfc318f4b912f2ce8903a216473f4ac0d606c08643b69d5ea11210ec0b1a5b4e1cabfccfc5f4320b386b209dc42f957ce38a328aafa04134edab32c599d1728076cde1710c9047f532046a4fe82ccdce87fef2484c4cb9020ca52da1ccb02db0c1a42489a0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dedd72f4cfc92eb02ecee6fe8f99241e35e3bf40f07860f4c113ce9175bb0aa18721a1a9e1bbc620c1b9f5a20b17c13003c537b1b3bcf84d8867e048b62d0978bd7c44eaafde635b54fe436ee26466ffcddb31db75adcbc24d8543859a6f7be600c8cd9b78033e2bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177b823b3aa5205d833d193f183bde75ae08d9993a8ca374e891f534e985c37fccbf5ec19eef84c0d07f4f03fcfaf848e6c7f405a218da7accb2371090ebb05461d2489bd7eb46fc705658790097449cc7b398a8dd18cbb3fead8b5ed8437012806fb518a3a2594cde5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8d8d001cefbafa502bf506e4c9ff4ac9d0e0e9130361d1083c97cfd194adee95319e5ab04290688cd8d6b04695683e64a585ee99b32310bbe5c5503a04142f0ed4426515f2cb0559dd94bd06b440315870203873c36c111a0a41e7a5d8886075b966a9c67c48bcca6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cec6f4008180bc9dce7733f0009df952f97a8b761b5341a02e23899ae4126d265047244e32d479c34c4c8dc70162d47a597f460453c7783249b3467f64d1c66e11d92e0427c5fb1f900f789b0610f69f14451896cec9e602253a6d2352d0e18ab790d7fe14416759a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1910ae6802733b60fd2438c7c974c841fff1786636baddc79a3a1c08dab7ed61720741d97e49ff98155085e4b24338739d5f158176f6e989c7fe0d3c6b456c08f1e9da0683cb65850ddc9b33a8a4f9e52440893bb556a62e486f37b13a940914071c9482c34b604dc04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h530d483708bafc111f078726711339975c44a943712136f1b4aad4e1f41b2e7fe4b9bd826708d847c9cf8406b786934ba9f7ad3666ee33270e9cae272d6824de52009c92513e8dc369508633966eb171a6e227cd63894dc41a0588113e6b641757f2558bc9e421839c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1385f4b8bbb3247652df953dad5710f2a10b9d04740da77cb4908a8cbbc211863ce580ddca8fcf2155d5bad191b4a5de79b468e3f88322c458e4297c5a53515722d4740f28dd2e0b55bde86acb446e26a39b34804d5f10e34b8d7d9cfaca2a87be90f2e0571b4519043;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183fdcd62ad9528b857f34bfbf3b56788b0d2670d019ca324e5e5b3afd6a54eb9fd3046f8e98b337877af154e9a23f46dadff1cdef9fc8f7d66a88860ce69018577e4d84010fd27ab170a6d5ab482ef76641d35f4b993f013a5038cc51a5fe0760b11bbf4545ab70be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcf14bebbcc6191dc64f24a74605ef336e14cb6e38e47c9feb539306384af083e3cad2247b6385098c9514445eeebf729993a4786cd5592fe69a06c88a3de19506f41b90a94e5252c2d722f44700a9ac65d2db6d40119637024fe81e2856dea63f5c114bbc1bc4e5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1745ec1ca21cc24358e7b49901d9b70c86f4c698947ce0e0d73c48c20b22c2e57e91afcb9862df3ce1bc9e753adca9f28c1c0bc8c0daa719e450d7e1340e5560d3361a902f2a538d8c2daff5e8e58ba2e9dc9e17561f1bd3120ff34267b8291af6a4de18a646285d8d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h699df766c6151b594d8ebc09c9b0429eb716efaa9b6406ce056fe8f0cd38ecbb01d78bea48ee4f298ce46ff40ca71c73e4cc88853b39af07c405ada21e340ffdfe02227d590b1143b1a6b90468f739c75045a9f210195648758a19c645e0e1e08e19047ee2366d7987;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122789267f9e09b27a993ddd1aba166769715fbe34c465134927df15796cf26be34a52edb6e249ea2e90117b05979b477154d0eab4ad4d27611beb52f833da107dcaf197395a07437fdb2b7466990941758e105b020eae281818cfbd6a7545717fcd5f8ff3ff74873bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde41f9a3d4bf242bd562c7dd65eb31f91f7a636fd44b19bdd06ba48aebc058bf5fa8dcf4a20a5952466c1a40093983c535d430d19f3a775fa2b8f9bb7d1fb9208b2c882b370aecdfdb79a5c97825d2ccafdb3e87875c6c5544d29592a16763871782ee1cc1919bc91b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd5fb90a5414d13a1709b946a353a2500d30552be86d94f0f22cf3fc89551ee62985901eb5c260afbff1a7ac1265d6219b0d84d0c4e8708cf4ede1e2e498a3b2e881a0f89638cd04e229e5aaf4da265fb8a1056be89665afc825fb16750efb3428eb5bc9c10dfea9d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4cf9bc48a30ffd1561724cba4fbef255a10fddf868f5513b7f5a17ebd89a03abf3f05bda580b92530366a278f76a8002ec8f9c659c5d9a6496f7eb452bd2f67f3a8deae9d3ae5240637cd24457022a66d52f532afbbc15047449b5d40206d1740f62e9de72058ca76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5a54b432697bc24499482c007883999048ebccbdfc7f8e09480224d5f6dafc781eabce30a83df9105cea7874e2c88e66e0e364d7facd5c544dce1b1e4fde0cce93039f67ad397e5b978bed11182fb2c6a928a129cf98ecbfa17443d563caf0b2a821f5d20aaa3a55f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13722a6e637c51ca7041db6291d5440f2c16c04db369ad02a0b160fbc17e460693c65aac886824ea0840d2c007a35bd69b400deb30d3581f211d95e7808eb9a0713df98c71906e42a5e7eb7b4588500edf5fa4a1bf8923c0b0c7212905b0ee0ab2df439929bcf991911;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe34c53817a905fd3d43c38743353284655282e0a19144054e9237f115818ef9ae7da447a2e9785c8ce449d7d8d8d5879df217a843534a99361ec34d2e3b641e7933122f21e8125f61ccce8595652e0fb1ffc787f80285312e6ed264c8351ea9fadd3e2fe869acd2db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1edc85663286f1014452bf6e04e04896cf8984f5597c91b5ba06c2c6dd38e74ca3eb8cad174176da1a3e7c84bc5f3d9c4cbc37a48527502f11547b7af8d75ad3485c32029333ef0ee2037085619023f7fd9c22e4e9958231a192e118039e9f1d9b1896180218de09f62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha24bf6535c282c8c60a4f2795ce6b6a6cf816f341c5af11d02565dde34266a68e62a5799093429d9bde82c5a3fa5395c9572c0ce888686d85c1e5f6d8de04cd42778312a252cfc717dc5f76a1f053ee6f50b058856aeddb249ef2bbc3a8bb7dceac41655b7e04804a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7236efee2701205924202de2455a7596329c8733abd46ede01959643f0fb321bd3ff4267bfd5e1220424ac93f7e7e67a59b909613d45e079da683ab6d0978ea0e5e97d7677ab6b119a8695d1b22cc3192a735d39c525380da1b77ddee475431aa336f2f682a9e875fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1989223439e9757470f3c8dd96c521643d0987afa7a080fb82aac6e9a25f4487a4cb3232b7bcc2ac71c78dbdd7ea3d66b5450e3ec5a3714948fc7af0e514b22168bf5c7016bcd2e8381746a2eb3ff844468763bc46c41dbf57c4fc3bef33555121393e98c9d92404cc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151b1850b224b332f0c308d53f2d7e8f0edfa64d972df4176f2c8490b8b454a6486050b5db346872027c787fdb07f2eea8e16d5e640328941832db9a512b738b963d2cc1efe34a75f9e39582d19ce13430e658f74e03168ab0218f3d2e0f39554f25f91074dd01ac81a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dfd5d14a20c0e786228df7a070edf0fdc70c23caf16a3fcdfb03a7687f19fbdc7f08da929b178e111aa12da3a8a1f185de2a7f33f33aacd7649746aa37bc43dc98f3b545de3b7c4af6b971592e5088fef351ea9424d8518cc8cd709d16ff78b9c9bca348b9b0c48fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9aabe0b950a2514bdb42b2092a51d846ce006cfd79d1be153327e9e3640e6afd799bf2033d5369538d85641cadc3c5abeb589951c133fdcb709d1c2970cf122b6108be3f110bd059b1297077f71eeb8f5003f2e89b9ee3b2a4ad6e86b0f818f65bac82c28a551341c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77d5b033340ff2b857f1fd8aebed4f5fb18194d397553a119e278a3d827965ae1fafdddabf9091d1a502499417600c29833408cfa5f176a393d40e6893f1a8300cdb1de35ef0f1f21f0f3171b36ffe5686ca88426319f8f15d9dbf1f5e52c8051c7c0e93598461fed5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d6e5ba3ee89410971b5533cfcd21af9c8b1e2820ff2d04d1d88c5d591b115c429251bff371caf4425b41d689d0f20d02e9401fae8dc166aa487a163695f5b761a3c8378ab8c99fb34be29ecffaab70ebbbcd09e319362c2d33928376d113bcfd060a6184b15a2d02c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5213091591b407a870160950f8e58d96a5884a19dc5d183642dc134d8d819c536f6ec42a6f819b9e8a951bc0895e8b62ab58b2f2143ae921a382cc3b19e26de2ebcdc5314a73f664cb319e7f298de6a6d37a1e1b259c7efaf25dc700a11c14c769fb70a9fd00dab80b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfe15280682a8be5e8b4191d9f38a5a1f5cee4bab9c3354e0b7c6b04db268e3e82c9c895b354f32002343ec39ff0b55c590061ce58ec130fe92fe8e2fc504f7dba54d99521a9c793f368e4f3346b66db7f55a0ca4164a59ad6982a32df64e02f96b0edf148b47bd3c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1398decab47b5c0c72beba8ce5f00e11a651a161e0efcc48d05e0df6f093cb9f754fdf8b3bd6f2c8bcee244dc66ac6c12db39a6a79ddbdf69002a9f936f8d07940ea22c871cd3cca3168182e108d0bbf4aa53ea4e8faddde3a50e1e88c34280af0ccdbf95c7b58c509d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1521b1d07052ec3265fc732150a48d84275ceca70aa5c98b13751b7237d6dd8d1ed64c7711f346351e1062b2fcfa735c17d5da5bfda11c8939f42b9a52f1b16bba58e86232a043aa80742939720c302edcf6756667b46bed72c5fcccdd364f012ace47085a819bc91aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18376dd05f8a59724174887db9d74a7e79f9fc437543cb0f7ce02894147a9d71f5bd45d2b9e40152657d6e7652b5197a028958ec111f4121150b896545c5efb4369d2f5b24c882e42ef2076f37126074f6f6b3cfefd4ba20f2f7c37db7848863428289d2864723137be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb508056ddbae786e7d2f9d4838a4553547c40298fff93f1d3e04b277b7940cb3854624b4c28d6c40abcd2654079655f82cbec1ea43e33b0215935e408d9a3470070454b357db48838f55a7675ac1b328b7a4a386fd165514ca9f376bab2a560e53637b35a6420d8535;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76b61e66c4cc3ef5059f743d45b8834890d99496fd923f47b2e01992837c279862db48fd4e3315912d3aaf7c2c43e1a3bac38e02e177b6a592f78ef700990c51dbf3413bdf1a05b534b5c09eb4c8d734c604d0b9e2041f4a9df5128f2b7ffc29cbde133d42e18a5f30;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b8b087a531d8cc52b52cc8b8296213d3bef3774cf91e4f6774fe20e180dca0034b0e06c2a4113e3dc3e49470b4cd148f70fc268eaf6ce13ce5ce595ce91310e91c2886084673b160e89db6394c91b632f8bda99ca0a5ed256084e2b7dbf5d6027b0a40d5494e5f09d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c134f9118f3f2c689bef03fb4a5e4ca839f4ac695deb6f13bca8fe4d7eb258f8dd83d59d21e7049a8e3c14052f92cdfe9ddf7bde23d4e8c58edf49ea8096b5aba43b97002e51da750f0c9cb810d3621cdf348d7ed441ae2ee2012c0986f1e897d30c136c9764fa027f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f67c75b81d11b76572e5b9eec3c1324ff00d73cafaa23d5fd9b392b45b2283190cb5bd71f076eea647e4f7c48e7cadb02540d8316d195e71e448f97cce78b6d27770374254ee01402f15aa788fd7c58aacd958f958ca3fc0f5c3703cdcb955c69ba77ae3a57e0893d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1193f8c1a2ac9cdc5aa48efee6056c11ac4d1cdd063c685076066ca56aed0b569de656adc1a8179858aea475a5df2a22341d0740be55a9ea7b2a7dc3160c14da299bcd6efceec137807d8051e3327a55fa90cf2b678e7a789d2428cd6d5a55b1debd311977428f9c6b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1604585e0a00904a83feca627ffc15158714c89c7da9e48017e40312504eaf7042f62d4362ac01bbbf3d143edd92eabf0941f1b2a9de852a672c45e8da1ed5aa25f27a865dff65b1276b0cd56f026a2265b1f8eb8c1b730076597c17b78bd93cdedd708729adb8e44c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18de2e246447b402a2b06c5d64ae77e31d3341484607143d32c769bccf5de71ae14a3ed0c4624da18fc45a1396fbf97b813f71a66496fea67c9adf95270c7a05e3c3feac71176b65e23f8ab11a1f669b1f974cc2ca980a92a09f203c088b7f7a0d582f6d2a511c17522;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3558e5134bbda778c4f4727c6fec5e43b18467bb13c311034c39ceb952bcdc442ca26c3137d9473d3b3674cd2e2a54a1aa23310ec5767a809a6c411b807368ca6590c3a3c202f206d5ce4a8a2426967d5d8b613ce0f47aa4fd85f8ea3d7a9837545c45eae26d60a1f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc14957a50927671d81a1685555961d5a3c597667814bfa8c3a0ae55f877aba6dec72386624f02980e2216511ec1867db3d08e4efa8376a1d83797f372d2b43396d58b75f7ae2651b22627798180b4b1467dc0c96703e00460ada05324815debdfbfadf270912ee9b09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d721d8d3b93a175b5d65a5219d934764a2c8eaab1c50030fc3b0268ac4ecab4142f15400796e99f01d9dd6e30082aeb8abbb822a3df40849433d56eb9d840c7449713869094174322d41cd04b8f0d3d095041d096716a935c2669a9e4e0d4f82ea5c1007a87bef348;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19fefab3ea881edd767be43d2838a6a97340ec6f91e024ea884bd3d3d5d2598788b6de4b1a19fecff2136e17ca2347d9329b6b43ad3fa079e35b89dca0e4bd8deb1329935c30e2c655cf0ec883a28d623d340ef900601428d4dd9efb629155b46779e592ec1ad797162;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f48318c5c189cf7c2c4604ec55bc1bd78ea2a1a7b997af04dcac766e79a179e1fbe0f0952bd6dc350adac59e2723c5872af5049ef85a383f4744bba5b8e56e95d7cf501e380f5dcd35cb14ce301adac57b94b451cde4d49bb4e85b20f678126dbab0523f7bb615a4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae09da0bb6f2cb505d262e46ada28b79a0106f2e47e3f3fcd8ac0c442348972a6bd796258b2d3b25e3871fc07f1a05fa20602060566f22a82915b2a48c1b3caf3ea298b7ccabeea25074ea65cc5775fe0f2808d364d2e6b211c38733f753f3490242a30d5cb507cd5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2e602fd9b8cd200d06f44971d00162198e689f4b4895992afad7e2db45b1eaf4d35656b46514014e8847517f00fb6476ccab80aed8fc7fc225dc5578fa0cee69c8885aaadcd7ea50f39e6ac8750a883bc158d951bf838206a52d34f49ea7ab25c355f3c412c033e9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13886b412b0eab09efcb84ccb24f9c5967f2096589707fe117ef6204ce511b7c8f7367366df512a2c9f07f9dd599decd1416ca3d41fcc8c64c542252881ecf8a8e187dad09cd6e0c59e84da6d349eaed95dd47e65d4fd91f194b57c4f8982d01d936a281e3cd89a88c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7f19d1aee4b6475e4719a8308a45534e231688fb24f487481e5b18fd5a72c0a61ee2e227463ca108ebface88d0a2964b49926e4752bfa4122fc4e373290ef20afbb3b0d367ecfb82f9f75c9994ee9dbea9660a58f2a06259b0bff8d4cf1a37f5a14cf1c3511d20176;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c71d042f1f881181a87dd8a972a1537ce116fffa475ea0a2e31550e81bfc5a079db6320312c538f4c51eb42b952abd5d377bcd9ac0a9e8c31e50747ffdf9124c847c5c655577e43f2997d6d9348a369d34392bee935740abba16b3f3c3a1adc5e194ca13b1202c3337;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fc61e2ef56c7844407fdbbc55d4a1e6adaf87e8ede5b36bdc53636572c0b93c6ec5684f48e26991d6f7f56117350f777a118f2e66ba79ea1b7a58581035778b490aa0d606a7d8da248af81b07c5ecad61991de302d3231c6a3754a2c2d320812729a20c23dedd4872;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d81add7883592d019d96685483368e53fc4f30fdc460f56ac58db2cacd8d57e0a5793e6afec02854449b5b11953d090a275fc776fde56fa6a57e6dd7cb90bdc3adf2743fbc837932d089d8506647858e513c6934173ff45241a14ae69d47650d07703593fd68a71fd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6c4bc3f60cd1bd26768403f6086ab0583f17aac9e2f9c9f67a56916d4d795a56d373a9e241394c39b7dd3a3b2598f24e76f89790129cb2bc8d592ee662bcfb17af2ccdf6d6bfc95bb9d4ebd4c3e3b61c74c1e60b60c96df159976884b51dbc97b41680262d471651;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b90bf74ee947be3c3c60aa73e1f418dee9b6c1ab98e2dbc4149ca0fe445337a6fcce8ca3f4a2dce3142f8653b5dc05748206159adf7b3df9fc6d047c1a66b9801f5ccefb2a393be75dcfacfd3f8525a8d427dbbea6a55942637048e8d211dc4598eb5ce030674c533;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6157de47e291fede15cf6731209d48b9ca7b96e8a015787e1661f68c8ad7fb06f02e3352fc030269a1cca892560fc13f09c7ef68948c66913e415d4f9c7b46c822f68605901effea641913d1ec4f09c652ebe9e107d7123cdbf570060046fbf3a50862000a32712d0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e1c556ae4b9ae4b57934d945be8be8e4f7ecda16fd1a32c58a2b0582b8125a7b0ed27eef72942eda6711a44baeca787baca99119a19b2923916ed08b66f0d1eb5487310ea6497ebf50227cc57e0225559728e477394841af33d97c553f44516b386647de476b4a8b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ec33631fdff16888a72f949051f90a838eacc0c2e605e3a529e21084ba3175382105c1cd54872f46ee91d2aa390e8d53a307f78aa10652c313f9b76fa5d4ff17b75585243dd7d8e33969ba3c26f92e59907e5193fde37e315d3541ed0150c0318d07171c3a4ee8a5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb129b16ca1620a86fa2589fa020a3b4df518dcce9f12126958507679d5a1ba4c2f94b1c762ca09a3e464db7ab96e30e9efba5a284c81c8b7c634da0fc4a8fde2c35235467e82040330376a3fa20c0aa7d6b3c56675ecaf0309d94ffff28d706b0499863141b99bc2c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8a682135231008ed4c56b83101fcde078ac4a5f0dd09f28397f00f1b38203157bf284b3ff4450593aea7d9ad270d10fa12f53d9d33a13b7cb65b404d5db2f157952740e4a706895a9275c8e65569f1fc3853860e87e9d2c9034ef117474d84d50d621d01e1d8cd5b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16275f41ab4af04e0fc0402157b9b3a15987f8eb04cd56c6f438795c282328e8b2237be292b8d015bc98a5ce1a33a86c527f29beabdc76bb056f3054ba184cb493815f321181fe20361ad04c35f96b59d8e750481bcda6170bfd6ea31f1aa1d075d083b1985a713afcf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4f8665f2c50c5a8f01b2f52bcc806de60457914d2078e5c758dd01747e798daa88af11dd946da663ba74147dba6c93fbf98ce0968c1802659962c69da2d14301c9d1ad308fc6a62d5bb1dfc3a60f9228df6bc6e3c7d24e88dfbabb535d8ad132743f060259e7a12ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bc482834da015034bf405b43b209399be87c9a37dfb5ca2216c1bb320e6e27eab9c4bbb682119689f2836975a1cb218df23065597e7f1eb83b2a80325b6e6873cc593deecbad0465118b23bd88978879fb5f8f476c53605f34399487985fe8d4f5a6c9f7fdca9d355;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e787099f1074e654afc700f68435576cf8f07848ac3885fe8f88fd8680276b726889eb4bf704478f31bdf39a7c081cac8aca6955238bf87c799a3afb611851ca5432c5153274f6e044a597aace7026052458568c2a57b1943ecb073e17dcf7c0d2aaf263179afaae0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1734942aaeee3aae611758d4ff8821fd568b5a386b1b9d56e6a7262a28d16bd48e1800f6df37aed714b8fe519a469d2164171ca751b18d4efaba72f8301d4b5764743fb35462d32eacdc7da30752d7c78f18eb206db70d75c76449833e5dabb2be513c7fb3a6b06b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd47513d1ba31df46302f128f8ba0cd5b1987b60d9cbcb35ea32f73150c4e2b05a0e3c2d4950882c2752ea7dc1ed309b0d8fe867073aeb45233823b7597fc88a2e6e20ddabf8f3720765809051fc58a73817c6496a9d08e241c99975957bd56a1a7dccf088eeb0406b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ff5c53ae58115955f17351c5761464535163b180a1ec9c5708b7244d3a55237b4d277155039e7b5ac6d53c319a8e97b6f7006f50b4120a9c5422dd5fedb712fc987664986c57b586e0313e154359387fb48ef71bfc3114e96c5c9bb3285244ea88efbf1de2a3ca632;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fee9a3dd888a589ef382f8ed58beb874026f32e536f1ae10b36a9ffea029bcceb9522a94df9754b2734e383acdc9b61aa82036e88c4de7c5d61b36164944d9adce4c8abb965a1d3b65e41a9568afd16cfcf234f168c922b9b8c34d949a42ecdaadf71bf9cc01cb0112;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192552f5403f0fc99c28cadb615726e15a4689f92ee48905e95e2b62c3adfb1e8b3f5b34d424258d89b1a42325e8308fc4f7d7546d45aeaa5c87f84575219b1acdb30338405643d317ad9e3984b517d65be28de7e15ebb3df99789f3b86a80c9ded047e4726c1e3c27a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6a0e140c182a1a6f324f34425a2fca38de93b3990a3b521d97efe3e5b78423c6ddf4eb366c09a87515b0e82576584a79593d3fa303c287845e23536f2022497bdd889451b33b2fae3645219d7b2ff8b9c6c042ed2e63512294d18feb2b32015f43f359bc54b4708e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccc3357e554fcd933ce2b8d4e135435f88a2fa6baf568db4a1b8b1c4da135b465744e7443ad3eddf1d194d54a762901b2f2f40fa2fecd652e3427d90c97294a8f07953c0ae08199e004f08ab10fc343f864ba285fc52170a84e0edd63247e8b6e264602b217c8f6ed6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f1fccd93fb0c03346da59de36fd3e568d6adcc142818bf9b9ccdc65d812365b16ad7dc960845ba008eb3f9c1ad003904667bfc66900e29272b2c1b2a2d9775842d10f50e4be7267264df25cb4268e93c6891edaef5f05fc0ae713969db141b8e2a31213ef0df7837f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b16f5338d582c6eacd9c904e3ad588965f0136a3ebd880f007eda977f79d00ac8525baa8b8b2b65cdf7e48011077155ca781f3b8c7f425629f672e17d69eb1ccf218dd8faddc6277046de25d63796e4d4c40d0b1fac38cb732491594eaaab90184282d7d57bc272b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153c477d2bdc8d195f4c21a5207ed5b939bc755ae3b093c363f65793dec35e2a9970e139fcce7248a6a71f699bb7185256aea8080d2e8c5fa3b050c8cb76ef1fde7eec91900a8df5823b66394227497f68cb5b3d96314c113995d04eb6d5c17d2ec6b3891a8ff27a1fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3afcc3b31e1b58d539cb189b1c23c4e50c8992e044a15719e4d9ba5a650951490f231e382407edbc62a39d0f8f1e42769e0ab0bf8c4376436c2bb50747b59dac2271286a14f8505876a258c5b688e632132a6fd0daedb86038a1553bc65473e545228348569f5549c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135b9090b7f2885075a16b96b21bd18e671ef9bb52ad13ef8c9ee0418cae59dbedb42e7ab78e931c0c57970a29834ed7556ebb727f4bccfd3a0354756553915e49153a31507fb7443c03efefa6f2b4fba5e76e97752129b187b2fbdf6af3e7fc4f8cd6e50c8513eb1e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha91d0e191abbe0e732c111c22df790aff9cb26b3f309c65257af2d555305441b79860b4379cddc4ec869c726aae4e2946b5137150f05a729e2add5b6612967ba3f0320ac518d9caa9c74d553073ed5e2674d053e5de971dbf57befef33310959222a00a4e7e2b52cae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96648c038a02faec2998f0538d53cef62f94d88a4936c1d17889ea6fb59904cdfcb6a5f63bfb1ba35b2e3c851810a107a2ff9016985842e8b7671ecf29ddf34a1e11e5a6587a40ac969dc49532631aceebfa9b7468570b9b4b962b254101642ae101acc127833aaa5b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a146a75dcbb7bfd584f3e613dae6b0f18141c0714a2f4a3723baf6cca5efb1204d7df91cccef957a428e4b88509d2cb675243d589f31f321525b7980d4eac72e8216fa3bdfee2b13b2c0fbffb177a28b3d0f25340eb623948d22e63f0f70217decaadb395f686267dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113b70aed81c19520f9cc7ada32d2128a7e309d7c0094a7cf835eb1a7f1196c43a656df1f9104ee038e5d9e5da715d89689043dbeec73dc2a68950de770e200668c471078ef6cb5a877225a4b0798a3490a68e80013070418e6c8041a0be39010e430247d3fd72a42be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11af744ecfb99d4517135601b9eabd26842ef60f946c41e3cc010b2b269c4de85b6ecc82651bc490edd7758c063c6a0774f45faca704ec5048b142732b297c78e108ed0cd7f3ab18523309002b98ecf26153ed99561e566ff21fe432faae44271d06a7b5afcb64ffac0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db8b01b208cef19468a5552b46b1d974e9d7e4daa554ca644cb2e2e299ddc8bbe5d0bbc2dc8feaf1af1d5434bd5c5cd495c8fede1d9d5fee85ce1fc80fd5a2b213299070bcd9c0be5b399a5b106f39238ea746ec109fe39c7aeb707bab1038734f99576df2ad8d663;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62f975e3babc2ca629f412e2ead8af4579d75182b37c3bd9636dfc45698f37b0aafc20a3b7b0f8e86aaeff195742930e9caaa4dac7a622184f7ba856962ae8cee2f4aa4559e1f3b51f3085871e896f59a74c289aa5a95c07957b2714a77d23afbaaf490607df9904e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b32d0806531f92ca855b636ba64b0c4d21b5bc705464f8e8536261108959b3affc134f7c7779245cc5703c0d23a79af30540e0237a4630bb245da793f339d25aebfedfc4298c90841b2f97eaa9e1ccadab460b03379d56e3de6eedc7d7aeefce6e040a77a6c7e7fb71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb43d5721e48d15bc314356f39d4c94069a956d6268f3892a3f1d6a5e3ef1232ff882163dbcc430f98839e917090ebf153dfaf73e5929a3955bdc31ac13e62c6b2973c84ceae7a96b4ab1fa52d15acacd665050dcbe51df1dd4294edfcba0f066afc513bf19ff6d7fbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32be9eff4ec18891a00b61e62e5474c9bb732ec1f27c8f1cb215dbb17cdaf7a9ffbd21212a3eb296e077ac351db1f0e782b5974f5a1514caaf662ddd18d416fabfcc36f42b43f0e3ee9c519044ea9cf83b0aaab7eebdeeb411c925e7a7c2a29e6d49eec75bb7684d34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba4952cff0181ecaa35ba9ef9a7c769b83b11046f203b07668b96cf22af236ec6d1730b5e64af74980e560c5f384a5ee5170c9a843030c4424fbddca8d47e77ab3014cb2d4ca428e2972c7c5be73177c3169dee82f8fb2510bae2a3be3e76c192248da5148a4039f77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec35b017b443ab42800cc3cb0c594d3e955be3a39106f12e65ced4e335279d21d7fad3513e3f5e557cc13e62ed4ad786e5a978409e32ffbf3a2ab591af79f3ad3b1294b051a7746d08f131e04d415710a420e7fae1c3e08fc859480e0c9923778fdc7d8590da9ff328;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b858823cd7a95a74668d4891b279c6622ba94e74b64684c16e758c6cbea6b372a2bcf5b8aeb40055ad084eda308e8966ec63df4963ed695121e6cc0bb0fb4cf92c391a0da44349da5dfffea18998b72fbe6e11acfd620d69312023791f754a096df66ca5f346805c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7fb76c8b50e4802502c848051a3b431ab44e4e6a400226dd9f8544194271467c60ef1d440579c61d5f325f5db80393e2625dfbf22546a3b752ea23713ac447c614718b2fe53ec796bdc7ec28e414ffd2d396d618f3d156b5457ac51e64b3a851c133756086ab3f04e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0d464c082f5cd85d963f118d4dda641793798d987903419c3fde320f97515d024b9a46d07c0f7f8d68dbc7d8f45931359d393c30021bbc6a0f739ec1c9b3e4ee64a661537e71673545b422a8dd0ec42e8e154b4b8299bc8de92a1fd5a6e3c1ba48374b4edc5482db6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27229b58ba1e2f8ab1ffbf6351e0210505756f6ac6914b1c9943eba88a25b1998ead29096a29e2562eed9eb7c1db8ec768864237a9ca509447399735fc4a3e1a3d0d7d3042f06e4159421e03bb19db37e4b394e90adfade8846eceae126c42d94066672cd52bb2a48d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a182f524bd556b2c576aff8100fb6e9992c69eb411db78c40ead0ac3e0dd6a19c056e2e756053b038a29657888a6b5d0fd35ca10203a0d8bf74d6fcf0bab0ae31a8f3d49eb41ef3d1223eaaca493bbb8dd0a34891a74d64ea45a1b5814d431c09756e372f0efef3575;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h419e22a5ab5dbe3f5fe50f0197474fd9cc3f15e931d76cc0df92f43ec3312173cc8c44d6fcfbb14bce9303a66cb7f257ce2a007bb43db1518f9bf32ede3d8b91d2132602a3e0082bf6918f0536d748c56b2989c3cabd5ab0f1e9678e6e448e68d5834fe49268bb1eba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he396aa8a3bf09143f4f491c0d634c44042b040ffcbe28fa346ca347b444bd8653579cfbb3e2c808e821d9b294a1df3fe80b96a13b0cd03c6d56ae7fe0952e6d98153e4f0e7368e5fae38d331416f1ca5b3f2b721a1c1f97e3b32abe5b68caa692870f7843cefa1b351;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h207083d6c4d90990029fe07ee9eb8233e72a8d4471fc4fa21e8aff82e4e5919541fd2b38c216c3326ea81d6e70d72ffb1b735922a789840a881de553fbdc2418a014fa14ca23e6b8aa9b9a445037ec0fa453994b137cea90d211b8ad257b380220972c1b2e09fd8d7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10dcb57cfc22e3beaaabffa43ccfbf703b0f0f51e4c96573e653e7f2214de5a1708db589a3e9fede8d791badc17aaae13f289aa863c20bca02c1084a3c54bb57d9ce41e4982c6d322d8b48aee7b9d0560aca5851c759764c18c9e1d55a97eb7d8a9d5ae262c42165199;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11490fd78ff590093f9e99f7b5361558410eecbf152df16690d804dd789b0f834f6c7cd89ca8f40cdfdf24c7fef6df940b905e79d0194a34f120a804723ac4948980339adeff940660e0d50e785108f662ab2d5f5128899dd69e05fce96b1d29c5f1dcc521b30f96bc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d890a972edc2db03ca1ca331d31940d772bb8053b20497e021375e28ff02cbb551d920c9356079e476ec7d515facbd4843380fb3514bc7b8d0c68fb7227227a4444f323ab3916faebee0a39a1336b6782e0bdb3555876c74445340b81ebd58d1d6bf8dd1c7f1d1c59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b58a73989964ede87b996b21a4f43b16b85763dca860b851f8bb2a5e8b7f815a528fec092ec67bcf901297a55d05725aaf33eea190dc7dcbd846fe6100754a5206ce11cf0f06f148718e12c7dd04ee65772bc2a029b648506f1c99a316c78db882a27544d20790624b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf159eca146b9a4a5acc6740c9bef018e988c5e74b8c41e7baeda0cc4b6e65a0e1ba7a416a5b8f8ffbc9b579c351c42fa6d6ff22f142655522286af8548b38c26b11959dcb8cecab6b03b11cd0c471dfe1f7a19d096c6b6c8390b05681c13bd0515f799084b8bf7a3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46d2109fb7bf810441bd3a5a9206b58b75be3d0ac363be0d0ca3f983d0f79e641a452d3509b190afc47bf760f0788a20497ae8399ce91282981783170be3d222d639c0fe3f45e106d16dc20b95d17d32060494642cc203be73eca2eb410d6e7776ce35d99a27f697;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h648cd36f9c3544cec8f1538c8c61ea709525b2e12c6a1aef3a442b52f388e1f4f677e72c81e47662fc7f341de056e25c25fdbacb9ed38fc2813166c08fe7835ec9509c86cd9fb0d99f9724c4bd6caa329ecc9f98c8f34a78aa3fd006d9cbf2ad6bdcad55d0071c462d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecdd605950fafd98fc77288fa5c6195569c3b91b867a674d9763a86cfdbcbca180840a296bf035e3ddb574164d0966856d5f677881f0bc7819b5cc337c68aa64dfd2497eadc1b1cd83ec69f0c18ed1f7121111c65d26988d58443c4b6839082aaab47ebb67f45820a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175c05f0f7f78ea5a0462bd7b7ae5d27fd3043ebd0428e7073f0075204f4f47bbfe796b794304730005b1d3aea89e9c79f83b4c47e2f145a04c19b0c06db42cbc4ac5d9da8516712e29aeb286e30fbe5fae31c16e112059bdf66ba22778e6a231cd35ddfac3f1fa2809;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a100ab9fda627ee979462dc7b6128d9968c0121360b99108c0509cc2fe7abe6714a20c35e59e7fac644658f32352fd019ef31111413cda2f4278cdb4b87fb84c7b6fa4f14038b5fb70aa186ef20d5d7c34a9c46609d0d7e7898682ae271dfe04c14ed8c8717f79cb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4748b67ed887c50123c19d179412702ba8df38c2699f1c4cd873859e7a7ffe936e0a2152e7e8dd81bad90cd807395594b322db56b316f86c0528fd9218488db6bfeaa1b18acc2d0b35e6973e985e1552c8b8d3196ad9f05ed6f8a54e318fe70b6401b5148bd59b61f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ccc0be3a431ff9f56c498bc263557710424f67258324296ac421af989658c3a38eb0f01302fb224e3a009f12f2b7939901b3b02f5b62423ed1e0684882d0d1e81527e7f51736d6492fbee26895f759e1f82b5aa277fd2bd24953de560d7227e1a83a8fd63c36e57f67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc18dfe33ede90f4815a647c10b71221cfdd2cd19c3bd97833fd416bbe4455f2e22cf8634c81cf1d8bf348697b4423d3b44a3d8254d55c1b8bd9cba06b92c0149d391362c9631d4df3882fa59a430ba09a25b43ce1c47ffec3150230d53560ea0f9fda0ec9cf70d8042;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a3b657dac2dab3f9580131e3c985db52345521595c7206613feb4f44f4acf7ce1d9a334ebd4454c829a7634875ae26ab9d3aae7c51cf9ec5c6ef91f03ee0b7290d7c7e05c29c0d0faba50c00edbfbdd9dd5685f4017bb0b6fc905f63303db61a9bb055a92e253b44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f13e0a28600a7c7d0200fc3d7f923e0c43f8c2eed00d1cb5aa138219abd7aa4e05246d44890a18d4398adc3cf868d3849cad75e76e1d93a747b3ac9775dfadb1709f4f48922da1b88a824b67c91e83d89f2c6368d75dbdd4c28138188ada7afd1ac410ee491e11fa3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9d1aad24908b5617c4340d66909d2e9365c2693c2512a9d2da1d96488720c385cb303e51b93ceb414aad6d815bbf20cf3fd5537c1b42587ef4a940a73f54d22f6c7ec909915b4b2e43c85403fd6b637a26378a936718529d6769a82885e7e13c0e8c7558301fb7a8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee9bd64b2ac3a64e16be9bd0fc1f013959c2b60dc194208bda0cd95e2b3feeb2f2475d226a8f1a6ed442beb7a7a4ef22dd08e76fffc5d0e6d1b69f9b74fda430a498e30ccb6cbcd4da1c4cfc3b9927d672f1154a3d7b91d5edfeb3bdf8dcb1e5d6b75c315368d8decc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha03268b691588e42a73966d2e56f3b030dae3fcbe53ead72d6c31f292dd5ff7c8e7d893fe7a2b3d2cb33991f26fd84961e5889c434e65d77383923e3f2418ebb6a184baed32845d28b4bbdbd09dd5cbaa9aad87d6874c4a8dc34eb61afb034e25491544f57a95e34c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c7542b9271f5654871ca483d8ac8abbae6e8f58f79bab6c193003411f3f9426d22a3bcae80c247c05b6679e2f4195ca55a99fc2510ce7e77810fe907d4b1ad9be7721e2c035df7135d2bb22a94ca691310d3f0d682c9e7178dc15dc70ad84407eac620466c7045f1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd77da31d74f53fd02079c719531172a67357cf9744ee5cc4fc2d393e6132159624e5de16ea943cf8337c241956e635f91f0836070f03757eece0f391236885bd64a3bce374608ab2a2e574510e7fc50283248af24dc1d3a6967624a1b01ee285f3af048df0c0798c18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b3b3db50beffa0e89c4ddf8b6e4e7e2c9e0db986cbbee5ccef55d2b192cc4ebb3bf57e721e682398ba63788560f249d57a4f402ff6489297a832c2e452ba75e7650ab8d49e9e0bcafe13965f820aa6b808983af21d3709ee021e4cfb9861ce9495a2c947464da00e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28b9a2a6804b90de06ee13ed42624242041fd2fda8f000fda1b58a2644f298a220aebeabf81604ab6ae89e805d6aa29ae3df829a77d34ef77e707b30a2d544172aa944525285ced2d22bd4a8d1033569dadf7463247e5138f82338eace88921f8310d82fa9ac421478;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10df6ce9a69305ea2d3505d9f2f5ea4c2343b081f99b20ada516e70e6a31cedf3ddf8bb71d3aa5b049709e38e88186163c0059c44a1275a2e8f985f8c5329bc637debf966aa1c98fa0306bf5930e4df117c71d0be89d654dc78132409e07f64b634abc558bb3514f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4b3c93f88c1f21d31aa33c48d578dab58ffeaa360a77d54c02a65c83282bc780d8c7ee83aadaea2448a20c4e6ec2ee77c8771c2eafbd5e47f67694daabee2d8542836b4e2dc69eab4af26e4ff95a9c51d6c56e77b88acab37cb4af2e0dfebc8a8d65746f09c1755bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14061f297e0f6db7cbd7a8c491091459698668389ee2707c2ce194711d93f1d2cddd17915722ab02cef48854e5bfd9a563ed1bf3b64a72e33d1e2ab3272e012e9bae56566b4345d2a175a36f8edba1757838c8655de5d078c281c443fbeb03e79e8d9519446cd4702e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1848e0e816e10ed4f02eb4cf0a130bab06fecf0314428a3d9b5d85abb7a0c5eda3b8236fd1572aa60b5428739b89f0ef0398db62eee0c035363452ec0c2586d3ff3a996aea39b6df9b574a1edae69c84619fa9704663366e0ef994020cefa529db11be2c81356dc3583;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13509ef0572401ceef219c5129631aadd8c2019ff54595cd2df421d35998f412bb02052f500ab5b75ad27f564227df1c20a47b969b07aedad6d8d8c2c9fefc0eac7ec31aeac7e7ac49e665b3c3582587a1de614925bb3541ddf7008662fd7c123040efcf7484bedd83a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fc839cd41015746b6e0c1ca9f08f2cb1abe6f0a507524ba1c90b0922ede841d32e57c6cf0573b4a4ea73e5e2dbe11b9bc8061efa25624825f46e0e42e86fe9c502644b4987e9cdcdc443aa160f77155983828219a604936614a95a50faa738dbc391bf2aee29a303f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166b0f4012d0910fe53be17242b26defac2bb50d9c537fbec6dcfab0a43d2b58dcb82c01acede5797534a3d2ee8dd0cb5fa34af5fff6938a20cddf3ac44cbcbf3dfd0a07d792adaec3bff46c8f981998ab7a89fb483c272d637cf5fd4cfd2e318f19cb172c751619a97;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd21fc9c03e94d113deeb3a56e7476d39f0c25e37ff541f1294e73cb3d55ed3d86f318ce1eff383afb7d62b0bba7e8ef2578173de4b7e4cfbd7d922c38d91b349f79c75362f5f3d4e095c0fe419522db6526a436e87ed71cec7d7b3489778503953b7fc79ff450721c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14da3d6cdd1853418e7d022447743c628c22cd7c58db4325ab29fed34c39ac9d78d294d32c4e23a0d40c9ebdce82bb7b7804884baefe3bad975df6a72ad5878f6e4aa2fcf08eaaf8e1d8b916bd38576194949de04f0c3e59d6b01eb9153954972489f2f1f98c2d9a487;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h24e14da8feffe9cbad8be7c218b9dc03bfb32090686c2d89419a06f29c36e0d00bca5097e0667772a58e064de70f3bb0ddee7549a112e83fc9b21bcb52efac92c90c416de9cd8bed654efbfd69d08eef56a9a3cf43a597537de19793b5621d725bc86409e2e420e66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109ce0e328a15446c5d8918a375c123b9d65909cd269f8beeddf2233ef3ae17ba9ee8c617e960ebd49bbea6c970ea94b3d43125b8eb039a1ecfaa2280c4aeac8ea52a0a36a69b0e71e638967ab5edcb6d39b5d92a3cfb34d22fd1d6df1972726cb3b462191708929bf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h314777344127eeaffee004d9fd3cad07e779a75f23306c6f93f8bbd7fb170c70f61b2fd5217421df126dcb8a7e04d0d32ded6e01c07ac7ee597a57018938e20beffe11af6b55c94597b74e22bef83d3f2bcb1c32a12bc745e912efc625b2ffafbf8ffc286521264faa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a824310db34db6c21fb58d393a42c00c64a8303ea10d8265f8a6ce4a66652afa2a16225b48d5f6220bbe891cfcb5cf075a38cad606667598132b6bcdc12ef4eea6625334df2b8b72ee459f88561d89df69ba073f495b9f09cd40f6e24ece0bb2dd01e3bd4e7afb3c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e6beba8f2dcc2aeca6dcb5a6192a8694bc7f18bd28b63247c3b62db2e6a621895458c2d9e6a2e07238098d0c998360d24e018e69523818b15b55bc7b3d26146f11df47df77f03171027dd0d9a5b701a9aabdf3d9b43a5c524121ac0e2a7a021ec33ec6d68e7339499;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce20f2097e8e71d1e487c89e3b314b8038888043838ce9cbf9de210ab47df15e05974540f7d68de110595dac1c3d3f9a0da44826574416f1396dcc8be4e0a714cdb7fa2a319ce67ef25f815879264348fdc05e939d3715b14053b74dbbe7d747f1242ef8e069599d3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ef7db21c5744b7b836a50b0e1f5d9a1b8eccae999240d26d6b1f6edc4148b74ebfc17e98efcae4c7f8906f4bd74a09eb63a3a8f373419f3ffcc344497c4a45a33b482c7a6a87fb94168cc05971e792c3b3add976d7ecb7dbda977f8923c547d643061dd0dbca7ee9d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h572cbe1959381be2565e71e4e9a02bb4cc4db0d28af25e96b089ccfb0f401eab1509abaa2a6d62351d21c10adccf6ba6d6bb36201a1ad5622c181322cdc62ca486d3735e4f1913bb39649417673cc772b79ca6e1d1ec9e39a2f97f5a70c115c45b2e74b25d6add208d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a04fd22fe86009ed07ee6c6ebfc6a93e2f50c443f90fe8f7086b6dd233d6ad7a3f700cb6268c614e2b5bfa4a8252e5431f91362017f2a0e51b934a398d41b2b7af05b890de8f5ed1b28a832ab54a47412314c5dd70a7edbb67f1293387100561750382662274bc8df5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e35293837a46b9e1500b90d26aeb00640de0ed12ecc43fab74cce0c25087e6f50437c5ac8b2173013306cd654549a672929a829ccaf5c6d0024d2b531655c6ef152b099ea89c98649c6b44323915766dc9794f6d21ca947202a1d33f365f6c2423cb5adde76e1cce8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h609e3018f70db935472e79d062f4348b17f0df54f0683029804a6421ec33321d3c7493c3bbe1220e3acb386d39f45d8f6b9db37ffab01d810d0cb0dbc5b1b5a2b41b647d8ac6f6b14d725a824f6793330534bc17d59c041be1762b60951f3ae39b93c3e4a6dac3b9fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164b82c4a871b1418a770e8422a831685c09d7d4f5b31ab41887b7634b479d1333dda52770a80933c7677ae783fa8ed7d76a078a664679fadc55bc54463190f8403f53a8df5299c6d8fcf606ef2f1e7cdef6b5af515ad739eed759f9ea2fdbb0a3de07defeb3dbf09a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1941e759cc6183e14cd2547ecae98ebe171c06b8ba5edff9e86b2c62bff348163e1aa529030b677345db83a5d0817f7f84c32d1cde6d890478e03260ddb8f2f5d865cabc0180f66fead756bb1438a01f0bfe792c7f9d4f50b3f701ee6791793b94d84541049770ea158;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6a5f364c73a5bb5279ed6b3093e057a8c6579f8b09b6fcedb84d3d8750df0e8b3c11c110e9be2ad4c51c70f799094807e8db91dfe227f333d4894f9a8e68d315aa32870d59d390c68f0550b6b5766840f1edeadde04a48a49fe3f77b383693c21a520e44251b87db6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a250e694f18496f0ad5f6bfc186b91eca289064cf009d217bfb1133b7d58861f0f8c1b8a4670c5304dbe9e72a90bd1548d24e37e955a48ee5db38b54ffd1c4b872278833ce2c54811f0e4992f110e3cd40ab64bedfd7a414bc0397f6947c5ea22cfa85b68edc7a95e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1994020abee6cfd2c9a5d54bbc63a1d1687d479b4cd0984955e7a5b255fccda9cba9d90992488e9e672f12ea82447be8fa717485652ebf7b56531edf6f7131e6c4d5704675b3e3f566af947c52458a929624f323d2bd09f553e4ab03e564cd022b6daf8ac11616ab4f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8ec183bd0c431d36cf4070c01e6f24d9d2024c67e66967fd3ebfb51d735f588aa93998bd1117c52962b6006c83523d03595518f1fb0cb2eb9744719eb2c04a740c39376253d5c9a80713a434d01b0e36abc1a3dec01166b39f168970aebff361bf15b0238af808078;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf772b2f0a16fa46f1bb53f827de211ef1845d58f5dbb3b4ce7f83a74edb75b326bda38dacd912ce8ae8361d0aaa124298ecc87c6271bf79a1dd98e49f958b48cbf2235369d0cf9a29110f419a087730c9f71a9b93e607ccfd38ce21a4baac716712da4d5923152fb01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9a559fbfe09da5add5abd41d502e658b7cb0d0f04a14b806e6a15337cda8770569a13b05799f75785d6d22fb783eb0fc2db30a80663439a27721dcda589886d5391bca5d8daf55a19cc0ade9ed7a0ce065df878728a6541b1d595e65a9dcc35403281a2fc45d8302f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23502c698a8e5bae2e9ce1aead06c0ba02fdbe5c88da6c67da0ecce1d050f203ac2dda81e3c4b2b4994f2630c0c428e786b5f32dc6a66df96f74778eee93d88624762d336e35bb73964d77365a83f7f763b1ab2995c3ccad55b38d9fa91b7388fc6c2ab4c158fe9e43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143bf71635f5a0d41d66a1c1fe354f52e2db5e2716b9665dba85c9af20533f2f8de076004dba1a6cf87397d95b80a3c88fec8f66e8b808ed58e972f623e22fde578db19b23d3ef89c776c17c9b7ac1a5f70df9aeced5525803d4effeec5734b22e882634c6bf55a019d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aef3808c842e06a110dea417486821e20159af3a3cd25733a19a497b645fd99080ae87ab52fe6997577c7beedc40cf73e6f48ab4a2a617edf620abe91e9361aeaed6cfe6430dd0916c49714216fa44b63f5072d4dd776824a9eb990926c352fcddaf6808f5d32f2994;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fec9de83a5ea6734ac659040e777727a2fcc8cc858c4863be38db2e8391f8edf771c9e1d3dc102861b5a26306736d79ee768b575c23ad5ec0b1b2d87786f286bf151a1d5b68fb4462dfaf7d1fad409a5f5991a67d6e89100a57268c62f92752286c459125f912c3997;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141f5086836e17b74f0f6759b94a0387c595f6c8c77476662632ad2a18f47a0b70af880706f74f5631442d9f4acf992a3ca09f22fbcdb1500d090f238a5fced7498fbe28aa087398776c48c42f20377c3e3e6219f8ba77cccb44e52303719227f18163fe73e6b55605;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9b55b2988d4de88db7da1b76135dc0721426e1f63189efcdc9dfdc7271bc83c6a002f389d3e2912c90e6f0c886705153c3433d1dba17a572e37663151e9ca7666e63908ec99bd5a8ca4442e6496e1cae830a7dfba8d443d1c1d3654181415fff670fedd716f9a632b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0d113487c566f0011f4902373a9b0aeec2e4602877314673d4ea8c0297b980704e9566112b067737d7b04ddf7ef25a51dbae0936f0af67f7dbb5f4e5ee9be0164429859a81395d4c60189fe2f00b8bfa61231389f81115b3d7d6ea1d1aec6614ff90fc6debba155b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1461f515eb5fbc2e7996ab706cadb7e9d4aa1bb8ae16872cb630e2cd14fb428a99cd77926c24b5e7c4dbc5f77cb8831482f42de415da3bcd5bf6ab173886828dcb56a39ed13e1e80bd9da91419248f6ea71bbc0a82dc285054a67b52bd9281069a26082b10f7b85c2f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c508e79cba55da3499e751eb01b8d877779f7505845cec934961b64cb9a92df76c77634fd9d898d2ed4c3548ba99829d3a7354530e9ac4b5321dde6bd279f14e1278fd2bec53184f18159e70bf4a379c4f45482e3d6ae1fd4d0b29f49f8434b237070f873c58764fd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1adbe2ec4782a6fdc20cd20a9563a6d55fcbcc887c090428172093f1420423396f27b920b4fded2cb29ac4e8a7687e293b3ef9eb6e05be485ae61d651ab510090cda098573b8fd831b283b39e0b573a9d96400ccfcc5cbfe0d95c38ee19f3c9419afbbc270043225760;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h909c8ac70322e21d502b1a6973574ad9f5b7bbaf53db278d5def33a51525f121fd067dc9ee4e88ab769a5f161b4ec2aabd45a14873c230fb91e87c64370d950710013dae3f46a0fa82eabe311b77148decf8ecb3e981a699785d53079432b2dcceb2268ed33bc25aed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h346cb225b67d50951df10567387b64e760846a6dcde2cc9639a75e64ab8c696bec4642f6c70ea337c25cab61526b13e39e7adb43b93a0703debf0b381534824d51eafa94ca60823aaf16a1f34e3d584403e148cf5e01b41ce3651627138cfe9947c197bedfeab2d7b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d271cdaac3704e65bf49cc10a900078c51556d300e371860b92f6cbda4173ddcecd8b349067d8d74b2f330559229ae64d96caca0d74cd7588428f8c92001dbc28d5089da800d224dfdcb6c3b6ac9186fbff520e2f99e90e6e5d4455ff2db2b30b01c0643dfd844c49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe66676c73d5c62acec03273df37e5390a94036817393e64cb7cf6a249192d20829e37f1bf5401b3fe4c933c9608523bffd5c3e30603f99b80b1e15e854936c56b8463de90acd697bf350a5ee6c2e367a1fe96983e990728181c1050f453d6867fcd1988e10860f28c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1239aeeb2b9731310528777e5e3e9cf831be24004659e97dfa20617558041d0a2c5f2a355200d300f6150d2c0c14251dfbfd6ada3a77ea1f45981e4eecd93f2793908d113082d9609d0d290f7b435445b081329b52e4b3d8596868590c98243c5003de5a47d53333b18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63bfe7fa5573ee0c394524f74d3588d12215ef97b4244dc111c5323a29638fd65116703ff5c5aa293c6761413ec756d0d66fee5d64b66324c8059254340a3ed0b4783c04b9acaa28184a69ea8e4080f76813ef783f5bee2a919779c2ce5ee854e3f9757bb8721d6939;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153544b339d2247a69910b52766e369c762f2ef2f7f2c0d5d2660255ee7a324653b7750c7940b5e36579a18746328dbfe5b95ee5c872a768b1b43d1a14109374426af35909fe4c01da6da54d05a8e580b7fc51f904d788ed14c06fa6e08715d224927b60ece93536a91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d495e0ef39d8806adfb51c5185eb666024f5cc8dc0224c89314610d7ce863d8ba72fc626fb7397dedc084d51987919ec53db70c8b062b2c29f62edc8306c435f11c3898677a9d353fd2e1ca5cc561920e0c06143be61b47dcc102cf50c5e59772426ef40d532b4383;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16914aa8b29616c3327a2b565d9fe12543c03d47577ad0df5ba96111302ca63643316ba933d7196ede3fa83bb20814f7dba99c0b6454dbeed761782b9a1f9acbd5f1562c30eae42be37b2e621d344859e53c09cbba33bb3205a7918955d1f2157e7f4b556dfc31be711;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140881ff891e61bb5135e70e7c3f73c4ca3cc3c1834a75a93ca3f01b40abc9d1fa3669f4955598692538eed78358e783aae3ecac5f440e0075e42cbe6597019645a42cc9cf630586719c4b1cc2058247e7e41a5e4565258c814fbc71a3b1acfbfe0c80208141240018;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fab207387b8aa2709b1434a9e3b489c4511e783c4c3b8b0b54630cdbfae1591d1c20aff8bfa0d9bb67f33b5553341e70eab9448fecc098c1247a362d0e12635316c5ca007e3a3e4652c9d81c5c544f18adf031174370784115d2a2930f09c5d37ee2fe8b4998e6402;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab0dbea054684a8985ed70e4b0b72e56d59c38ba5f42ddfce502660e3f3faf833a30f97394ae1f3071093cf73f67eaced194acf96d68c3eac4e98518d17e1cfb2010af7fd3e74f4391ea9d0f7a7b375d0edbb20f097f6442bd960b479da92f47ec84ae23c1bca519b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a9c6ad34c2a01f6fcacab10a5d07cc2a831788b25bd2cb566a0b1521e27ed73e1d69b0b09613f3949b40b28087a1c0414fc53e147c734223769903349806fb4fa8bedabc41975e85e3ed6e37459a3d4ab51e74dc3691fbb98733155f2345eb2ffe2b2df8e146f8203;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2722caf08dce8a26ac6730628734acd342eec43cf3faf069e39cc7cfa410e20566aac5a1bb07a453dc6ba7ec04307d74a90e79d4b6a83d37783dadc70ecf7e569786f5dd4e7302828eb35ea862cb2cf2c96f1be63bed7b49ed3488f7fa60614224ba605c762a1362ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf29183d371a44c15f51bc74e362c53f0f620f02fa01a1ca057078fcc124b9900904d8b32edc4b9553d0e6624ed28f9529c68014a10a22e4b2faef3444fd46b9724d7f5334a53dadbf031b1aa0ee8fccfb6054b27dd0eb939c83bbcf653cf3935a0cfd1fb9788d7938d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbec824f545dc1fc6304654fa76843f82482d61740dff5d539b546d0fc1a214e5b5092ada22cd86d7514fda667ed64588cf20a6c78a0db2dbeb7a941513c7736e0e6b6360eb3f2cc792e19859bb82267beb28a0ad84d10493aebe39757d7439c59c7b668afcaed1aa9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6858c9a081e29ce768e3a1d1c9035b7fb98d3fd6aa32ed0e031f01296ab28e6d2010d199ad7dbe2e72b9fc154d6b61c8c5484da52cbf7a1b9fb2227aaf32aa3448c12b1b640067ec3cac111739abf3463f1a04b5c38d0d79de70fffc56c4a9a0b6c90d663fa94c7d4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0cc4321b1b3bb673c449e31d94299c0ff1ba9d8332507b60f6383c8bde35e377be64e485abb445ec70760a281689e7cd45e5b27cae5e7cf892c3d278e37ce9c6f021cfe0ad0a5efa51296cbdb9067130f21f4df479dd91392555dd42adacf6b67efa0c2e10e45a141;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bc749433e5f704df2499991f50bc765e164d80643ecd49db0b7a0753326f873f71e855398b51e045bad8ee8ef98f3de986ef7965eaa112fce968adad1a5277577d2fadbc5f0b3490d7d7cf1d23b71b0462813d7357ec179dfc958e5706d79aeefa78502273d78ef85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148210c693dece79a46011394c3644fc960faccf78c26dbb91e032f4e795442df516c631557e44a600558e05ee70cc91c080e8b17e96943cc3724018ac04f88f09b32a60b07ed8a9a76d4e1e7aa0095b1a7245eaccfa7d85507a1864d8a0f81287bc8798e6e3d37235;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182ab25659a7ce65b2586500c82e29eae7cf9f64708afa96c747fcb2d3c3c5027ad1c55c43876e0b663954fb3e62fffbd6c264530ddda8b05d306da0eeaff7f2a185fae8fba6d8f163fd5a8c765039a012cf64d92d74c3548708de670826fd6a478f25ce501d61fd3bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2235674d50bf3fed39705bc7df60aff04eaffc97b6ed44922e31ba90953a728ead9b3917daf0297c3d706b565ea8aaf82e24a0b182e0fcd7f1a3d0fafa0883a8ef3843e6665c188ecf585911b1d07e86326d2db28bfe57d6b04a426d23a0fbac91855364573f211e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed289e0647c1d686c9e9e84cb6d8c46089307cea965aa2695b73fb843de0648e03c8841b0e0e3f49a446bcad49609884005bdcfe3619968691782a25354ac9c3547affb1b4203da01498fa3cd2635b913842f902ec15a4ee65f5ba1c95bbe6ffe85753cecd38105d69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cf28668f66f1c50f25b9acdd71835dcce68977b0c5cbf4adfb7fc58c322010dce3e03fe94756f8526d3c33ae25263e7b961832e8260a2bfe27f4780706094b87464edaa6841c199359a3422daeefe6c766f91433e21a678880d1fd45f1d8cf7f91d0be43804fcaba7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149649d42f24a11ea57dd1ecef355767814fe37a870a6e247b9a06f8feb57ee776e064d2cff689b402c765994a5911c641d8e0ce5246b3c7c40b091967516f0145e5a54f9bb7860dec3e3fab322bede2dd13fe8dac254d81a10b9768a84a294550dbbee104324170fa2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5301815294b34d8cdac720c5bbdd6930163f024fe571e62e183e4dbf711659a72ad827701ed9c292ecc1d463acdfac0a0454dc33b2c80a6ef09148f1c6f0fe0434a2456e55b06dc78825eeaf6f41f264d1f1d416dac9450aab82a4f8d1e783eb487a3844e4b2e0e6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a957050c45098ce3d25b6d04ce9aef20ab18a43069600c817003e86354d867ff41e0ce1e1a27780bccbc80c95dce0a662a798b3a61f17d36a60bb7ed931465b2ee5ecdf10902918f2015771326ac62f5fba45b7a97d1083f3ad9d0caa6ed3ad785ac1ad843ab2c4f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec72b267133ffa7942ff03c6301975461df425ed88f820b3506c18bf4fe37f6ce407f569fcef70c9e857a25d78ac8273cbe3e03fc7976a3b43ece429b434075fbc34b8b4aacd14f2c618b36b80e5d7b5c049f4fc46738da9ea5bf9a114fa89b8ba1c4a35497fe76389;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13eb17892a3bf3e3ba041b49eab7c79418e3b93ce9c6f27a9e53779c1b8ea478d458bcf438f75271c4a317707538eacc16d74064c06671dd09a11ed40bbb25af4146d9a9f4d6dc295a4578a7fd2c13836dbb27596b2886726bea23523471efbe9ab7e04c68ba84df9a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195044ca523ccb01d262e1f48d3bc48459b7a822742bbe26f992f9ae438e4c73812bd3426b03aaa360835e0c758a808e7f965249ae7eb487b5d67c42277b4eddec1796cee05307bce7000797a663fcd8902d6403c73aad23a176f5fe68ac1aeb9befb1e8edc76314ca9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2565ff64708d49941f12d030226f86646fed757549dd3e5b49d7302ace70303f29217486ec2a540f00979e0a5397d3840b859f323ea26d370650f7f8444370cbfb5f884a33df6bd65ec1d93fe81981a90561ab599f1f46260c8d43bf1daf61a37f0255c8cd1fcb935;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bcde06286d7d3b6f7a6004aefb6e7ce4bb512d1c793e23a889ef33836d2735d7354a829c22c6588183bd25ea8300babb538696281f55539f3036625700c0fe43a76276e72602c2f875175fd74e1a3083bb234ed690f4465eb2e6e7ab6393e25440ee2310d47804353;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5e3425ca7578dc822ae5e128731b9ffec602ffe84ad24120d3da0c6713f0f6614a7b85ce6b3d856140ff601cab78279b57a999bd7fd693dddfe803a94c4d2ab0255406857fd0f204a1db45523a91c0eb9c36cf27d76be2d6cd1e0ab74850a3827118ed9eee160486;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145c30ec7597593b6842f30929591bb92ee98a2214ae44e153b315cb237ee72e28c5d1cd2fcbf6580df47b93e93022e5ea7c524d1b9d50331c77a135602a26293dbbf1ca14a16f990851179faba8b247a35ddb8b9ecea7494f28d6cf2ea559c4100466771aa4889990b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10abb79a8b869866783b927e6c807281da92666f2a81baaed7bf33b13b9891e9fb21452cc8927a76526b2d1cecd9cdbf1a213b0614f4097dbfed14c1681167eb759641c33ba36522f760f26d5d17ac7643d5f4e02d48701a68b58cb6b9a982f343128063f771f0a8f93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114c1fdf3eb02781f71c1b2df1bbdb8b23b56a377679b425143a41a7942eff1dc6555a29cb9e283411051bc7dbb029e619254e5a349d82cad33172987eb13f8add51fd8ea283cec81674806a9eaba6fe0b54bc6feb3204259bc74e7fa45cc6d824642ebd3f6dd19ef7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c13836a99f3eb5c9b2d1e14a2497e55225125b94d7864f92827fa57d6bb9da05abbb3929e676717d003b7c3c06b58718ce05c089b5394fb67d669c54f7f2d291279c2e37a578dacfd789bd10ec66f77fe50ef178ed3c9fd8de0a867ff393e7b0d021778b165f54eef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6a82c75df8d368166c0cc62da91e40d042edd6f01388da9473a951cf0d43c11f53442409ad31bc666df6ff286435fd2509181c04d737458625a281647c99b17710898b50d4b93ce440d4058f61393323615ff2f9b4d7db1668238038f051d1a770e36e6a164949f05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1378631b00dae5ef6ab3b9070be7dc674beab3f33dc186773df541570e2861ca43f6b9e45ba8f5413e445ca9a6c44c0b4bf38fcad24f62b471cc45d9cff021e3888d1d37692cd84d4ab753892dfdd137420c47000a504e39c0e377e166bd030999fef6e6bbc73f7ffa5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22015f39278875d90b69467dba032df37938735222a6c447dc023c599144e79e04d3b876965da5bca10495d0fdf2d9bceb6d59abcf38e3d917e5f9b081d83c8c98cd7e95a9cfd5ac75e80103d9b36524ec92ecf4d16a451913b9881304eefec73936a7d52b02d8813b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62b58edb07caeb8f4fb8586a5c401ef3ea6c3117d9a60039bdebe3a5925b91780ca88c8421f22fa125138b7f109d73d35a2cbaf1b1c42b03ab3c12bdabb387091a78fa94370ce26577093e218348d165b5ab1519dc6c0719d7d759a4c10e4dc193b195381018f7c5db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e674adbb3564609f593b1dc251e9e50c9c2f7acb494cf3486c3278a3c6ef8fe52ca6db108c4afb401a37425ac42db017319af9c9dddf047bf1c7b4b1ff40bc86edf66d66d6c5bdce2deabc0794a9107b65b7babc4f107723fa5034ea457300f5d9741a0ead135d8fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2b99a04923e979247e1087c341cefe44f20c92d0ebee11d5d8e1080ae80356fd74ed1b54f3ba58f4aeabac3285c88531dcaeb0074022a312ffdd314f5066c82d9c65f25fa23569ed3a080c2dd174b4877f0c677f39dbbd76ee6f84526ca4b53ce3da4520723264b29;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he899396cc902135586ec103d2b85e288027233e535b38004c9c1906026517125a7fe7207f7d22769d87ff7f21c14d6e8615cfacd9b641cdee1f004ab8202ffe2dcc6dac8ed20b1147a01b49118a7bd79fd7d5dfe60e4daabbe902a2bd89ffe9b0c6e79c6b5b15fa21c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c49e2b68a541971271f87554f255c513c0c211575a0f4c4c90415fd635b64b7f93844d067035889f1feb1a6bcadfbb4d9e92da94a271b2d8767872cff8a7a8ed1c218666d391e22b5e41d441a9a5da187ce66efc8c75ae82972464431c83228a193b2a58691e3adcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138112d6c429c99ebd96067610c854a29e7a9d9d4b56d063ea91555458f21ec1add1a7f6faad920768e89fa93896c30cf2f537ad0db8f69cfeb683f503c9f1083f6aec257ea65a40942bd9fb4f7aa68b03abb854479546f8d951f8a21498444572bd2cd6a70ea4b223c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h516c476bf60662e5ceeabcc7dbe40a7773c4f243c3c50363f2fa426633999bb2d0ea31a27824502068b388a732438ad386b6d466cd1e26e3f1a32fb4316f3144ecea7281f82adc6d53358aac66183118abf3514f89ababdc48d48ea4fd2d1b00d54906eff57d6de655;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1986a7dba603d4b65d4538e517981f5d16252b14fe58be182be7cda29061f0eeb7c229358690d24eb21c40c56025b6ae22ff37e83a837296ce19c05d9fdfad1063f13870c742982fc761bca9752490afccef7a66038885b31f29162ecc3f4c43f358677af577723db09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfebc90ebd89b93b6ce2fe9db53379489ec6cd6d10c069dbf8bbea64dcd2276f15a7fa7ffd4ab003a135941d4f6bf989eb07ada393293348ba919435058ec9612e231cc9b7d4a37d17238624e550a2f52db8be9cb737e75b3264f663088e4b3ce3ac65c9c4dd6cb5fe6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb2f80cf4b8ecf132d300eaa6061ad7dbefaf6e9a918789946d526c64f8b5ee16266df0d1bd246dd70400ffc23a10892d612f86bbeb623f2a19f653cf7379752507911285ef03cd2896bb00d4b7a8dd81ba41cca3cb2c1ca18b002e79e5bc7b2162e2bb7ede31922ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f239c35d07664117d1fc547a893d9082361086fb09048041609093a19975d1c371e07169325a831c7d2fa0fede057e8acc5152d64aec2cf4af2c54cc40ddfa89253f66dda295802a212960760f8de90a1db9418b010506fed72df26193c12f6b07863cea42c54b2ff9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf4c995c9475c25ed3a0756f30e291a5cfe5edfb8ffe495309447f880ea0d45c205c2547563e5720521a779f6bbb94957fdd10bbef4e8883bfe4cbcb951a094b7e1f7071e2295b9862e00dfc4c706b6e1e5726fb13e2285f8cc4ac16e8badeb2ed8443b5bfd210f852;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1492f3ead4ff1dc38d229a49c7b5a6e43133cd031bbdead53b3178880fa02f6ea7773b68689745578219e38913958ad9d899122b6f1d8ff20791f57f74384d1e1dc0629d8936ca9f713527061c9a7ce4cbbe9ce6230d3b6004ba33f866afa8413a92e696b3f1e109fd7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148559e207fb67c22e510a59210cac61c0abc1d551f02198c5dd3e334c47cc5c12e8c6f175f041389d70c99c9ee75e4bb2f461e7e7455f210f33fb330c45df04dee0e054c1570cd000f25cedfd7b6403235637c925f0ec1996592a7856a8cd2a674ce19dafe9c076231;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee1e25af840f1209bc69a8524f6d7a5cf84d11cc9b00bbbf0008164fbd1391bc4f50dd3002e91842d63cd2e0fa1826a308d5279b6cc1f2cb5913846d771710bcf5095150d44ddedcf18db56ca96ca7474855b263664e28bc5da23193086ce1c2e66516db178287c3e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7bbcd7d44fbfcbd02c753d9963e05581e472a33f4ecab83db6652f7ec44cc383470692c8d5d34227e8cc03897f42df07165977c8c8873ac9eeb0cce705ecb69f8969033dd6782223fa2d9a4c7ccc9e18d5d881fa419803e86627da6b48056d2acf76c164d2e2ebf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hced45db6ee636605eebe75cbb90e3008717a145443bb6413358ad99c70290f97f1edbe5266d347db01e6c92fe172152af3e8efcdd5e397273471271bbf37a68e78617887291104b2fad039dde94a93bdd37f67cd73ac1670aa75abc519ba579fce1672455fee50f062;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9e03df998404b943bdf053340bc460be74353f1b2ae9c7a35ffc9c375c04eb3a8d7bfcd55d2bb42fa6d1465455f489dcb9a53b9b79c5f9c6c5f0abe7f08cc91eb0ac95575346fcacfc3b538dee6d39e8d2dce3d927c04e698716d02920b97e63a460da7f7e94b8ac3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd91c78494bbd7ef5da1dc2ab96f762d3672f7e1489c5cb11b0c313b72fbe09a19b087c36591c1f485916eac94194c10b806124e2203173ba9fcb2d8501bc07f9369392d8d94fd55290c85be6cccd094e2e3b61716bd0b8e8ff76395f5a0184f8d0c6be213644836ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7d76341e42335924971ef6fe8888deee1be49d7dbb76ae5b7fdd522f0c3e59f446aa7d15105127aadee506b2042e7712635ce2b7a6ef6b2e9e1047d36c8599dcc59e9b97bf548d27831b6d61b116cf074940e949e3578237cabb6e0e0191650fc5c04a4dd312d0bf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1100051f3dce5659716e6685f22c551904fb11e442f66009bcd62987621ef86155f96a967ce92422803e1f8de22b92df8a193d47eba23405306b27b5a1b1c2f1fe8263f74c177494bb678a6071a811c44f0ebced5655488a06571b18141d107a218440e7578412504b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a69ff521d58548942141d60f17aeee9da4c1a9c60d98d8d1abcbaae2a32242373cdb27bcd71cf2582f7c6491cd7cae503df6c4df8f931a4d6eb6cb20da345238926eb937efb0abebf2fd869d8f1ba72bcc38fb9cf83366ca2009e04339ccb653d2fa7e280ffe8cd377;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6649ebd2ffc164dccf6c8cf5046fdd4c915b7db1df07f7ac183b0b4903361eaddeee49a50de213d29c5e62358bea0c8ccc321e4f21ae6759836ec2d4f4e2cc4f8e0bd0da4da853a1f134d0f75e066a4a7b0e7f719a133ebb007c690e2753815b77c472eb9af1deabf5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16505b940a57e3334bf15130d5f3e8734cee0ab8b59b3ee2a32455424aa78522c2dd346a0cbba92fabeeb52e569c71698c962e5d5d7abb3b37a92100d969ad7c38d90143fbe2b6fa79aa1ba760d152f90d962d9e9b069e76836d53ea1f36dc549e6adeaa14e7c1b45c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ca348b8b49febd956a7bcc354826cca8940a58082a57f42d08251cf3e0cd4ccf1da397b6c0c9b9300ffa07f017b65401e246c5d93e8ed42b559565b4f1d1e350068694991076c6db048430b675de5aff61c039448f84cf0eeaf203d8831598be6d5a0d6fb4e83721e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1992065fdf90c1fe64943af5ba14365b6095482eefa805ce60a32bbe4eab7ad51b7f139e5735c65f0a3184a4bdae368a967a9a102796e610dbdac4e7a8472e6c32159dcb535707b8d0a46b7c6266c14ba0558da34efd12e1a5726abb69974ce532992d0e32933ed1b46;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e40209596d92a64cdb36f9f51e5c3f43673dbe4fd9e4054e167e44b3d7679922ec13cb6190d1e6d6f8d03fb46044f25a0a7c81cb0e429c5308a2aee819d33a7e0b0e305078b0e0e3ea479a474619e453cea5c57300a7f098163c8b296ec7c5c8b753a7412086a379c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d21215c530dabe2ab7a61d6b4d6e8e14842571a923c7cb73da696568a9af6281fc909fe5606022ac27b5b47b7a8bab896e70141b844372d661b55c802be48fcc3a28336878854f6b986186949c5917c495b7f9d68e46cbd11ad918d4a56513258704cfada37514478;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb016a8e32ffb7ab974bfb0a8fda152b74ab43fcebb7e32949b6080341a4c1267b48276e3943add52e0b2fa1bedda1fedd1bba3a1b4b48a7f62cd29e144713d8e49aa0246dce89f75614cff7dee00fd02866481432a240e902e3c8e1b79071fd8ca567a134e1b35ef44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38dab26539a630375758a501c10d7f0d1b38bb76b5437c4288701fcf3633e90dc54dd078d5c337440c586c26b458edc1e056fcc3443116df0e1c03effeff99e876a4db08e2c61ecfdf0affd8c701cb3a28d6b987ad4dc6cc89e7a5d796482dc187a56ce24bf7ec5ea9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40762dbfd4eac594354bd38d25ffc56e698088a78523e489a79a3381cbae7a4322c6e52933632655828086ea78b30e9b1299bd2f1d66716e6db3a5ae645831f6996151322cd91742a98dc50e8fc8cf7ed36c4ecb07253409398a79e09e6a32cf23af74831ed85dfd34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bceba2e2bbfd5f31eee6f26539be5126b34b5d88eeae303fe937df14c96e79f22ffb66fcfb07919f0cb863a6fb8a9eb02bcd69cdf325411b310594c6b63287e57cc2db5d7b48995130c0f431015f8644aa8d46e57a0928916eadccd398c62351e7d728ac7a46e171b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1325dc063a40312d6bda60b90a5c2dfe14307ad599af691011bb9caabc8bdfc81a5bbe70cbef859aa9bebfacd947a957bcd5d8790ade36fad56012b8fb195d035d1e47177563447d705b98b109de32ba6341303737c10decd7f02b2fcbf55ad26c8c64965dbe454e573;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ff40bcc408d20724aa6d31218bd319b818042af84b33c4252844660740ce814cd417057a3814e29ba0aea81f16346866c34b9044fe91418583604aeec0da2a1743d3abae06919cfc2a859d98d8df7fa02c01505b57eece727db61d9855d9de23a6598b14155df712e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81deb65e517196de06424ecd203d15b33fe6d515340cd34643b0ff4a7f48ab93aaa51870464f15e904668cb2d5fd5e8057831f54cc8cb34b1d5bb514a1491812eb02e2d79cd01eb03d30b2dee5c79911e9346c4bbf98477f0bb0c6cf826468cf20a606dde65e785bc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43ba8cbe15a8500387277e622659091c7f7bccd14a1ac949ecc751ce02f79f9af89ab3eedbb873d76fc5271c44dfacde991d29b15b1eb44734287bb7f2b2dbb5360b39b44ea0f7e456f931f3e1846ad2cfce16557f955a3f9dd39f12b3d1ab9d26375844284523a05c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4a19bcab882e8b58f6949ba30902d3c0bfba16316ce58da5b83b35fdbd3215acca7e07c7cab6431e1d869a3864999db370a080d3bd11d310e29342e0c340640ad17ac333a5efbf9eff0acde87ef2760ca7aad334bc18d9991ed31436e0ec3cc3bd749c6ed46987e5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e26ceb08e98d36610be711a4fe21ba121b155ad8dbe6360a3013f607e6eed4eed1676e715e9ddb38cee50d163701f89fc2df8a9f246735e8ab1b363f7d5c943c2faa28beb013d11d5b2d733a60dc1e713f1e0c85657c80c179ad63188f6ee0adfd8256f339558b73e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146f2720c216a894242ea5e399deb242ecfd502df886761f4baa2e059d16cbbf68812353c21169bd203ceedf1f4124d68cc36452abad995a857e654cae0dde88819140ef6ac0f0b314058c0de19f00857b1c6022a9ecf064eca2a0df9994376d77b4397a7f9e6d9ac39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b97e3728e1fff9cf27ba4d3fbb33fece965617afc0f082be5185bf6a0ee546cc68eee29f109a6e300258981c3f467269f65264f332d83c7a060c154ab36c1632e1af0002cb3d3f76eb226c3fa152d04223b852f8aa843f91002dc1b145bb6ec5eb341f3749c2f9a6f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h436dbe11e4a92236ca662de3a46e614247b70577ba384b53016c3f9e811f2a78392c41f44f062795090f3ec9dc51f4d108fee6062bb22647adfa1759ca531540b05fadfadd9ec008e65049d2388219c913d5fb0e7f47bb8cd07a3e9d4b72eb4b5c8464a32c8a156ded;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b97cdbc1348ce86026cdacdcc27ddecbdee2461980b57a7da5f7266adb5c6b883c6e98820fc08be871c7baee6ced72e2c160e96c32bb6d726809778e981f5783bc9690fe6ca89991f43b4949b564f8aac821c5708c16f992ee968355e8f5281ed45d6fbe2264eed4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58a3bdc2e12f8421f8788306e5b185e293d7cee4b21c791e2af7a778e54aa18515735190a64e340732a73268a6673aa4f912c77346d901d1f99443355d463a6c5dffdad15b8501b6046c812b5acbf28848e4d1b1dd34f3137a43b1e5371678d7db451c0a77b535f861;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175f2e284b317d88eb14fe4ef46e339c3b2485270ee13b707b538806965cbbab31bdf16d3184194909a2b7ce5436b79af1ea8908bdb073cf9df9112d463e1dcab6fe774c323f2077c42d32fb31c3948137ac2d9920319ce3a0d442262443cea9a250030868cb9d3124;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89cb15d15569385cfe782e692f88374e35a0ef8f3605d56cc67e21483b445f28cae2b71b7953a69641c73c5442c8116d70b93361cc6a16055713425d34c62790fc823949f8575f05515012fc76c694b650adc5a8b92f5b3bb02c46150cfcd20910e67a7017abdf545e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75de421eeba01c5473730abe1f84819f5cb24211b7204479efd120165a015d92bfa6e543ead22feac45189f1711382e7eb427fc6206205f18995e3c0436610eba05516bb8b98244283ec50b69c871a6856c658217814d45bd5a51d753f4282e8592c980a61fd7e78b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1131206b37791102619212cd7bedf0dc95c36042555bdae24ae579ebe1967510c902a24dc2552839c10ba88830c8767a57b155075b79a36f8ec8edce2248c71bc161a998ae6d40ff162002a75f3f268e44ea7e7639b3f4a0c6f92eac9341d868d6386fcd0e74637c565;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0f95576b330c538bdfb74f842e3755f6bdb2632e4899e20b5de077cec3aff8deb03356021b8401b7de6f75d91292a22c4750668c72be193d531edf82c483380c067976ad40315820454b053fe9fbbfaef69f2eb842e9726a3f424656cfdb39072650aa5f85807b0dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1f84c7ab76e37bffb2d4de02cdd82144960a901db83ea6f594db379b1c39cb369efc132f8b2acf04024cb5324a7e884c1e3d1050af344149694be4a9368b2c17034982be8b5040b11bd0c74dfea858cdb0797f6d83c9c763d59867e877a672a6cdfc5182a9950b91e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136be05b5263b16ebd16b4e76dffa794225f615f3648f568e5035670493ac91227cb1f6b972612bff941f54e93f9f796f54d1687918483e608c3c296be5dd73d47543ec5f52fd0e60b88ec1780ff1880dff4c39a533471934809a01ba0bdb123a1be90025d9fe4d20bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9cf9fd77313fc3505b03a329036b38d67753926475c204e7cf8ca2b561efb5fccfdbabbfd51fdd595d0116653a16ba421bf2d7bfb29dbd9d03f19d7862064e803d1f1b9a4d8f86632b57ef8dc2bfaf85cb3992c6a3579c5c8144b1ce96c96b8f26e8a674ce572e324;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfbf9c5219df1f75a4007adba8c0e94784b3115f753845456810c6dac2fa7bad7354517786383ea960d1084f05bfde16b0c41ff080535f059c872590e1e1180cbbbeb9c7e3755f681cc85b97e4739a9eca31b3623aa7bb5f772ba2d19d5a7db0bebb5b01e549294a36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17646651ad6263b0ace099dee42c7e1f6dea901b864c4114754d7346cf4a66071de21c6831d11046a2ac1009db67a86038d126420c1601bd88ef6631fad51ebc6af7691df5b139f4f120c9c7e084c474c409fc3944cf474986eb035eb518958c6c41da3015d924844e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb306119eeca1f0ddfa5df5fc9abc4676a30af55f5ea37853a37f1420c4338de97fae52a2695d0ce9ebfba2e5170a8d169206913b2c363f08fe8a6e7c553c89138d738025fe7937c6c29ec91b5b19933e706c4fdf53ae16eaead312901fcf3bb279e09e7856fd4ec8b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h233c16cb152fa184212f94c0a3802a39d02b26095507ac0aadf83eb4ba4401c31c47b39b7ba9f319abb570d6b8d5d79312792e04fa50fed7b1860485ef65054b4c8f093dd86bef5afc1724b5f13bc3ece8b6914d688c4bd6f5cd78ae4586328b422a0f2c93fbb9c350;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff21d5ef0c9eeb0869d1a365561add5c681010a1c8ec5a72696eba572cf0907df8e4ecfcd058759d255c58cfbcae6a8f020f6bba776d01d6d3be0d51093fbe5b219bd4171311378e562cacd1b6ce671297dde42bc117a9c1444b560d4cb4c6f0067e0d41a1e1c7d855;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18276d010cf4996019d64525b7c6c7b0f41fb7e8d824823866b45dc530c4518cbede5c182efad8fc9fb998426dca7e6fdf037e002e4def9f981db2263a37618e36e69683f26ad4cf4b470634af32a8fff9ed6a3d0700865a3fc5fa98a26eb879e700eeb8b23d60c252b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e05f0fc9e085ca8979664fe32b3847a3ff8fc29cdb1a0e4fe52da005d8dc9d8ea04d1a9c03374a4ab81b3e5b14ed88ae1f06fb84a6b1bd2aee6cdc59985644946d7118ad4379aff7b1e344bafc62d918c41ed6ca93d325c0920a6ee53d4fc2b6699ad5310ef13e36b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b55a1ae6957baabfed879374d4038d70653050fc08b836c8de5c09aac714141e7bd4d96e66d7ccf52d961be1d4d3f79fcf41db2184aaea9c3c461e45d5e17983ea5c469aaaaf978ecf30901dd665ca74ceaec53a7f1f0dbe52b50b5af787b718e3679655b14ec13f39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbde1c5b083bff6b63c85061780ec85e7edb93f07679096035949345441b51050c67178843f20aa60c0cf26b51dd1bc8f06067148937a7fd4479458a56a924775e74d7bfc197d4f170cebff4cc340f2dd94051effb907900d956fba7c6495ae7661dd231648bd4d9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f7ddffd3e87de2c31ca935330604bf90307d9467281b7cf03044415b663d8762951f4b5657c27bbc9433ed6feffdfc321e12f0cd8053e574d04e19a61bb8c0221febee80668dc1c5eb9afb667f051bc5be08c608473f1b8bb00ee732e4bdf80316a5aeed3490b8f9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1952c7c487455258322243ce5f660e6e758e7a64558a8e215357eb302a8507b26db6f7805875d8fe10ab7ee1cad9aef6e52bc6b036dca57e3b2193ee502c1f55c5f1db7a5c1b70d2e2976bd6b5882b5a0a0a60fe811371a9648a3e35ba81105d16013f2752f4c9b9dc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff2bf6f5c903e4b976b688ad88d206dc82f1b831e6b6cb74044a11e5f1d5d84732ee4dbbdd90eb7423322c0360d4d3fc07bace741eef720de8bf2341e036177b4dc41ba688d519298f1d2cb844a2fbdad2aed8cfaf731be3899f44d06e9d49e091afdc9a099c345f07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d520e4044388629363b873a4a157d088769677924b4afc931ecd321f9f91322cba4cd750935a755b8dcc567a8e1d9fafc2eb0b6ef82c42ff7c390d649af81c8fcc2c73c4c7b7e9b0c2a32f6e5fe9642c4c5d6fb1746282cb856b872a47ff9e23624bf7f1a17b81301b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131e4ee7d0b5dca772f49ea543707c3ad8a6d1349a6ec0578b03b9ed7999bf4d8c0eda8003d073783faf56eba6641d5dd62cdcd86ff54e92d982473d694ba201040fc598a3a3b7263e1119d9c5b2c0bf09892d43eb431a1968d5a5ec1513f0beb7f0f746c37c8325e1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5973bb4fa0097a04981fc86b16804f7b212e9df90e1eecaed336c031a58557216cd9ab8c960d90c7cb38534b5f34b23a65cbc8915c10caae670cc24267a97fc19cfe23ca37497edf377f13cc332e968be929b0487b9b8cc966da7a15ba81b40448bcfc17d2612d880;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d7daec005667a8b2934ef3cd7c00242556bfe1ff7240ab2d621bea24bfa12d3f6219ad27568f44cc574d0012c74e14f1d19df228b37ffdbf47e3e537fdf4aee978b0190a35ea9b3b085a658f2e4391dd027c72c18447652700ebdee700e98b138877115ed00677243;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b266df785e65fdfc0dcb51c0fa3c6918eea90454b7cd7fc607e16fa91fd72070163cdad4c2b81c032af1e1d6e7311a6b12d702aa995db9bf79d47a8914213629f6875d2358853813e8593e9b4235d3d7d82fa45220955eeec99163f208eccf23823765bfaa80cf153;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad3bb3bf145a0e8186d1b168d9133e1bf280e2aac83d121af60e1d05662d3a5719feff38cbaefdebb2b3f94450d7921416bca03601f45330aec36ef603a228bbbcfced134821faac5c92a775721806f52cd6e4a51fa7f50d79e0a74530dd907f3ce7bc670d2d66791b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5073c7a2a9b437b61ebcf5d5d8e848515af3e0f840154007efc4060d14e57a40c03cde26f7f6945208e9893b815d39e507205e3db5be7f5cdafd49d7ff8e8db8b9213315142c5e1199e87d57efbb643e68b26840703a7258c9be54867b2ffbb77b7b3aaebc5c7f564a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce9cf52783370266b95202a9c6960bb60d3a3204d7d08ed0c58e3ea8925b216b87f2044d55311b5b424fa0eaffe96a9f41e2e5b112fc0b7cdcd67b68396ea424f4b861c9e17527b53114c9993eea1fd5b1600572cde7cf05a7a758b3e25690654b8343a4d83780ef62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e24262aa6ef5f9884364166546d0f8c080fbc79a3089e6c8fe601a7ae95087ebd82bf1a54715457e6f26267bb98e5111700a1dbfa968c26ff671c3e4b438cd84ae7134420b0a195d63d312faf7229c6c40d2ba65067d9b31651d938f1e398c0cd043efa9afbd70d061;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12711f2eda73422d6a34f77e60820d913142caf8c4435c0cb2c7e14da9488ae8dadc49e84f7a6b6c4635f8ec64b8cea7649bbc512c2df67cd5af9ba748f7fea21cbdd62da03d598803f0ebb039c97379b1ee54d997180b3f8d8bdd76287764b3af81c131ea7cdd06e43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f772dab0a0923dadfbd3221ef1c5bc3232befe2f28bcc0fef13b4516e6b167b0f25d44fca1e2d3f3bbfe44dbe7ddd7d98c90fe4c67eba77dc0a19075c6ba9c2018bbbb639efa4cd9eda07ede6f45586838968d9855368a691258b57eaca4dc5a3cefa8526e26464a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168eb419ff6e6d997a263670eb78e5f37418fef1c81fb942ebb538fad67c72750c961ba055de941daf88b0b399d34a5d848288fea90b61fa9c586d767014071cb15a3bacf5e428215726d04e32bddaa28a2b4a51f15e6d036ba2ecd679cd1072ec1d8605f789898ed9d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ca1d1b0fa732f97406aa0c7e86977c2be86f867520d24c88aef296a78bdcfdb1d23b2c5684d10f15f646ac84cc3f1bc4290dd8fc131648a1cc735e13a2a1c27714c6bfb7058488242097aede7dd537836be1838151d7f94176e0d63a1be47df9b5f795db0373f3a39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfd560f86cb897fdcc563c03f17c5d0d15dba4f7ffd32a4ade15b7c12fa06048964d118f693f85896ba9fb978622944a1e5959e9f3498f1b193886c276a59d93d851610ffe2a2468bde98f06e2f43a97adfebfdd63587a839309ef58f5607f24fde0a2ee8c46528c3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13da8fa59bd9be56b8072b46cee9df3c1a4f039454ae515a2f12a4d7ca1052cc92ad0ee40422272c61650bf257f87003d958848581984db39546c436e50e27a3b6c9d56a06a53264e13d96930a678c3d8b9401eaed5535200159250319fba750f19bee217c299c2b5de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16998be6c116b62ff263fc1f36d4a90af5f3d7e921efbe9f94b7156986088885e1bc547194315cf9e5ef49c8a81d9aab517fe87abe1c743cfd38f321952644da0e1b3143797cba476f12f25b2a88ecc1f2bc4cd6097f8608c03f40c06223c1daaa99c45bccf0468d6f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h442f68dd0f87b528792e452aae3a83a739ada8eae1380241a8e2f96b0b3ba16c696dcb0153495a149a63e5d35409b0558823b10285fda52e1b14229cb9a3961ecc995745849006244d883a5529df07994bcc8724e15294ac6057a8cef9225d639ddd50c668ad6c9e32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h859a6dd71fc68244e5a582c8830103b3b3030035fa8f1e0ea16fab2cc2ef248f4c3d12d980af1dbea9ce96576ccfc4678c77e76351dedab1283799dba4fe645518392f11411f78319ee38f694e1f631d6d5e49ec0bad3abd39aa23071180b6cc3d3eb79aeaf16308a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadd513da66d3bae772ecb454d222b5705a7316596152543e1040afb04fe10c2143e9b16c9b00074bbb07be1c424b182e1a8db0e6c0f02a053ba8056fdd432ae53eabf226dc0c4e202618f9057fa120a381ac2d30afbffab1b829124f25613493bf3c7d1b9f1c21da97;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1633d4aedb02a27377465ad8f276a699bea3d593ce9f21a2f44da632ec969729cb6338c35c2c8ca1a004924efd5dfdfc7b77f9525793ee33744a9b42788dcca892f0b2cc7f583deeb416cf9f1653506c162ed6c2d4e1ecb685524ce1b5c6047d4d400ad04de3c8d9cb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19995bb903486254038fb3922bd9bcf9685aeed2c966452d4a18fc55b87ee4118caa21874c6aa9664a0ba50364fcbed49c25ce398b26b5a33209ab7fe27ce37e0d02d1d61c4b7d5c980bc4b84e6521cc8d237d8a073daf427d38d6ccff62544c1cb0681050ff34aab7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194e15d59cd2ce0ba2573fc45f4490a2bdd0c79ff475913488a92bc342cc67c0743cad7fad45d489a3ad94269b2e5334714408d8ffc82884678ddf337d19dc8a05ca16bc9cb46177857c7a032bf420c026f807206ac28e2bcaa5fbb58ebaac137d06454275320c20d37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68cff13f6f8d0d3bd6f225b3fafba02a230e4483efc7d784d01d8818d99e408d129667118b6e0455be937e2c4c12903c195260d9c74f99af085e5d9cd2a3c181faf8cd2c9a971ba5de46e15ea54ef4191e26217cff7ee00825cdfa2e90e764e25bfbff25028f9ccb2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78e6bb1535cdebb8ab1b4dd5b6487c6ea9d14e2824ec1fd219bc1f2d751b4fcae94dd8be8447abf652e0e9bd874029b4163f2283d288b74ba0126a50016688469f916133352e0423c79089e5d991753d2c1375f9097015f9c8b2ff4cb80c662d9ce77d94840b8862c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1185a83307e0d60cd6b0052ce69b94d3ef4d52b1cdcd19c7011f0af44f3d301a638d1793b8a2ad7f9be4611ea3763f9b62aaeeabd684ec0468b469b6c61cc319e390ad77d2288f41278fc149927b328cab431c4fe898bf83e9976ca24a19919dfb20f2c7a7eb155cbd5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10cf5be9e9f5df84fcdf51863771d66a72e7f2dfa35bbd793146aec7515b8ccbfe8cdd7ed310eed1e619e13599a861cfa3344e733b03b9d4dd8da9c1dff0620da27b63a26aa114b53aec9e845e082595f89d495584d14593961c2724857877122d1a996f40b3f5670af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109842b78c9498cef404028bd627bd9292fb882e7b53cc93f99e880258c50f991406c0932895291d7d9e43bc8e81a68f3d8c0d3506d6e7f506de6dffa03f424f7bae1622e3c51780cb55fc727b2a4a1460891fb62abe3ffa089f1cc8fcc2759253297a2fd7d4f5a32f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1cec74aec3c28d5ed2ff831ae87257c26fbea65f1128875ec13cc5be79fc9526f6a0f77b3449d0c33f895703262f03806b540d27c48558fa6086b8ee3f8027645d459b0627630ea48f3096333b5b4a7c20db91b043df442b92827813d0f8ba2e09c7b93bccbc0781;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193b6506be34636d0cf1a76394e9346758eabe52eb422c17b3c7535f69a8b2856dbf8fcd66cd8d234783afa8b280dc8a801deea3a2b546da29bb7f2370c2b8ee68c25d7cdeb089b5743779b8ec5e4638bd3ff12ae8a6d2f34dca84f8629d1663aea105b2d7d8b62f5ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha43fac6e70c62bc7cef23021e26a0a7a6bf4cac86166ad3b4c27c5852593c9dc54188228d93399dd871761c67651650f08cb8ce69895ebafd82a4db53f6d7479183d68d2e70abb8ea78c6eccf7352cce007734a49e8803da469bbf849b3e26f46cc2046924246e76a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1192d2e39f32638fa7f26bbbbd32b1d1ca2ca8e7659ecdff5975c825cfaa33b33f0e5ac02758bdb602f6652da6f55ee52b0e7baf8e909f77e8e371997eb5886abfaff326631f10942e935d0f57f194d14c03be10033b89b803e0d8cad88330e376a3f578aec79d3a8cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab880f134d0b8c0bd3716513eafcab7cebc1643a450b45102b4f6c000ae1c41612eb6e9125b5bd559551d497e65622851fad0a0218d58e098cbb90a3353f57464d2e8889d711cf793076d24ec3ea6409e4bb201cc159ecac161a3a593fe92ccf546fa964450076440e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76618d873195d8989889f82e6daaaac8a7be3f5d1a6ec0f8f50b6320ec66585ba2969aadb576a8ee048d57636baa64d18fb693baef8308680d8fd6a228b48b85ab9ffb7bb8b6c101fc841ad842647d3f13f38a87991dd7a175bc22e2195c35c75e1d9bbd676dbfd22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142225131041fd13b2f911e72349092490df2ffc0833c33890c719815bcacd00ddb1d58828c35793e52902e6a414f17afe97f854b2497e5c015733d8f08294a313d3ed55d664a579d063fd51e6cadd09418e7530d6ece79b7302a467e7c19ad0a7ed625231dd6e0d529;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c437d7cd9dd470f23998e417f960e5e0b516a94b03e57f03119381a8a56c21e8c2ea926bd3c44b865680e63f3c0e7140bbdce63e747b166da16bce748248be0268e2f73a82723fc2827e76f44cbd62478e5ac4062a21c6a664221d8f4d0b845db08b07ac9db5526dfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a786bb419601c75a131e9eb5eddf559295a49cc2d040308ddebd3d7ad282a0718dbee461dcb9501ae1e8bb7b892b8bfcf41ae1f6bc59bca295ea9d13d0847ebd9fa3fc86afcedf4b4554b4edb0c17e1811f0ae899753a3051cf95f77b35db87e5ab024f88841d8a2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0f06434ff36be7b82e409b8ed0029df7480e613bb92b9219c7ff8c1010a472765640cf7eac8d760f8c2bd930bfb1a18e1cdc425c25faf36defce31cc0c8ab5a0ee4c77cc985d347e216c7a48fa6f2895c481314e9f5cac3777927e8c8263687cab6bda48ff40410b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8141aea0a5d1392a05c58b92458d4bb17bb5e89a817f42852e71cc2367db0296c4c66bc1572bfc6077cc52176ef438876627654da5cc97ce4928edf55b444102ffd1021cbca3ce2f392d3b7d19c0f7308c90f1ef3772b99e0c4fef6ed4ebc068e7db2a709f9c5a6ff7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187ab5f21b32fb8b83efcae43fa01714f5d23d7e29f1826e762db5ecdedc291a2303ac99f20113db026b6fe02ce577054b05baf16d5f14a676d3d64b98316e982e7d67e1610914911346073689d778175f1735a5c959cb9ae2e04c442b4e1d037337811814140537da3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h676322bbda89dd16d9efecc7a4f1567040d90c3ed29ca20e32e8d869a141f277d3861f5965207c875ca8d2471ee211fb3c37b25f13067567315b92d2d0131ad7bf43068c68093849891459600bc5120f3daeb69e8e5f42c401e02cd71a54bf32ddbc70dae01e9442f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13eba40697b66144876160589d77c8ae9a78091b2967668bc207c708c8ee8644f937c1f67d1c55dfafd800bcab973c488bf4b8fca685f9a22ead5931aa90c12d02a75dcf0fde6c48810c6b19a1a253534cc8a6e350d050266150707930e377e6f19040b8f3b88b53f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef9863b14a59ee40d545b2707f5f258f4c48cc6a6cda1e032c70afdadb76d611c88b9922bbd28fe10b456e40699b31d362fa126be12d3030c6e3766f34eb68d302b336df926822c7764f84fddd1a5ebf37e0fb93286dafa7bbfbc23f91ed4792f972446a4dca5e4ddb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hafff445ec917720c3ecb2d6ddef9872535cec15eff62fe09fe238090aaffcc2d26162d028db0f68a258c6d1f5b91a2633e68b1f250b5cb2e3af84e259b90f6156c77b531b8d473398eace1d59789c17fb241d00e3d4df51d3155e25e6db0d227df620f3a55a6b1fff0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e670015457dbbd3e4cabe3fda054112eb48a0ac3850577088c9a05ce20b5b5a1114b2ea8abc63daeccb2828e76d62afdd095a5246c5eafedb5f74659280999a29e12f325f8ee0d80b3b07f3976e9e1bca29edb93ec2c269eebd013df318c3db2061373ca5f29baf054;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56cd88fcb906a3e8cdd2bf8d6e38958c7c6b715d5db1219519c9f580fca85784b2bf4ed9d9f720b077b19eef32b8c47e22269513711ef5a43d41f6d7d41e3e1a10c706ab12f17f944b2aceeec35d8ce50ac62c9620f665f6331f208ee2724d3ed497ecfe499ed9eedd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168517aeaba1f828ff3936e70cd220b4d29c20ba993e17a9946660835919473603cf31d8b80217643dcb7185f67164705409d7c1b69dad028ddec59296702819d27cf1a656fc5ce40a16703d25172a60da69e468a8b4dfe9f1c7fbdfc9848f9ebd0d8ceffabdcbeb3bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25b073b152effc66959cc166e78002fb4e2b9b145c5cf1b84f5d394a026797a832122106a3c182532580d03c4b37d86c25a4b15eb5e555a3232bf8d96de587de2e1d63c26708ce9ef63cf604d29691625f1dd879137695dc4bd298633ac6ac958fc7d7af14d66c992d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39e05cd6feda6b4e51ddf3422c9ef26450690677c482e73391d7b7b01e4f2fd6511f04d2b842e7f07145dcd17ff283c1c3ca39b37f389094da800e9eb7862a02d106a4594bba00d129a66569cdcfa768a693267ebaff60bd0ca392e1bb1f5c2f85ccc3dda525e9ca0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146bc925b58e8230e1ea0285b7032bdf3bd29cc9a4ad2a85c7de83cedd5581705f77c141a3d03728051f63c093485d5eb84a448c18e844a97771b679d367f907efd84bd390bfe46f308cf3b9e6f8c5506f403f7309a432cdc39c68e0638a7d75d55762e81150a896085;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h726ca7a14282430fc8b5166fc1bcb5efbad309ade4c37ea8ebe2e47ea523667c0c29a0db3e641d46f2d4c6d8b961d0362495eda4afd73c971cdddb18e0eb11b9fa1d2be325786ab67e0370c64ea7c0b12cf6932ee1011498493e21e5f22f462152fcec29d04dc654d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b3781c4c4e46144bab176f69c6ae61309fd955045e7984ccff8f42c54ae8ba2bdbb54b12749ef5a4aad7c322521fda9c6a980e5db54bda6c6d4162292e582b1cf7d101f45ce5c53441443487e1dc0b7cbb90934451a977997dfe686817289ea0296fbab9721c9a5cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15fe2e455720c69de789ff7ebe0e7b08e2b0460c6156a321d27c9f57fc017400e4cbfd4e50e18ef3b5c68c6fc2552da853efebd61f1ed10f7a2e08095ccea9a8e52b74fb9aa5deba74e403af9c32b0eb402ddda72e9c08c85b9067a703c3bc89c65d2140e93fbfe5bfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17753095f4f97826952156d531c57d157c2ac2c90d72bae628148fc72e73b481bf133aefd3a3bcbbea1f9d0c89e932d5f7a5e5dcaf9a330aba496ef2665147a70774be6573da49af338bfd5dcc3e99e74c1b0eaff050bdd1ac87956add64c3a2a96b82b2b1bef48eb1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118918211c18d46db60408e43de2dc84d673c53245e4cfbcee5584f613062cfe1e3c375ee1b81c8ed7b4362c40a06667a88fc286ff08061fb206a99f0a0bbad526ed2aa6d94fb526c6ed43c54b2477febf5070ff0ff5ace904eb46885de16df2a4f8fe40a19ba3d8e4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c37c6c7caa3be7dc6b0ffb1f0be9c6dfc23f3b657616942d05d990384a083fb26271d09c7f1819dcee2d77534fe6695020f424c6481cafe800e64835d11caf3967a49eb737733357f804092dfc480fa482be7e556e2a8b66b2d5e8a3c67fcc0e5d508ffd81c079285;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12852ae74c78f21a00f1aa70924a2ddf3a3b967124b58e0dc01ba996e7331f6ba8393868a4025b7855849752a14f78b9515c8d73239dee42c1d2bba480fe71635c8769ece9a90c0851e6fdff25f1ad53620508fe99a07b2804854b78c9e0681e69413142d4568179306;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1498f840d24851a7fd6f7c536f5a61e8799c5fcfb6d35cc0a304cbafc324af3b538e3543e496cd1a0cc42004ba1a31a9f308981d44ee3d992ab522240cdc4868be5ecc7a06d0974d417db9a10d6984907f3b7897f6cd8b16cb2d79809f9dd2dc2f972517d9992ad53ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c72d3fd071533fe6e67f5e791dd5360580852996c4daab75f2a6ae7d0734b203b439a3e684c933fb4adf632093d48830116af5a562f21cbc2766c20384b6ebf328458aa87360a625712783e21c05c2b3f0f781bc037dd6e9fc447caf0e56c0330cf70be99b75241b91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1585d2ce439e3a357797ad5f68e73c234dcc4a7ca84a4a1025a5af390c3b10040d95b7d1c1476c1fed6addd1ddc8f3413668b080505176751059ddd3e13d8b3604aa397c7c3268aa3001d2b7f7b77805b571473041b8b5d354ebe8cb3db82712629be3db7008a2bdb93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115037e52ea782af413dc5784795834952999441895a4a0c5ccf6a0e3ac8fd6afdd8b69235faa97967d114b966ddf524c5a68b148601f80742a8c22891fca25976e994698abc6abd88d04328ece7a06f76295d7c2ec4dc919c63eefcedc259769e38ecb843ac18477ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c241225818c31fe082c0a476cc98ef07096b6ed7ef1edd7230d9ce3c05233cbedea0f3fedefeb9d4a7b52fdecb93ee2f3f30023396bee26e38b9a474a82d8fb1d23363496a91d56bde9dfe6c14d498478c99195f1b297bd8e51f8839b2e0013ec419423f96416060b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe56801ab024664036d2aaa6abd565416d9e95b6c9edcae2460d3ad9b67ef2f537810500760769a0c16d3b5f1ca0867bd1c63dff1cea99d545d07b9149b0fc52b9ec83abb53a1a5888896f231e8a8212e69c4c249aec88ad1ef8268e1792c43acec831042bea9fe05a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d7bb9a92fb7a9be93cf6b24d82c4fc7d56c0a81c6d372a4075e9275a9f3743b3232fec58ca96b654be0b6798373d7b1ae2b96ac0555a366ba88e4adc8cd6ad9b274fd2d100c7a9e789c9db786142cbbb1a7bf21f42ca57a985738a7b3c4841826284a4305e44dea90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169fd5024aebca39cc36dd1acacdc98898229ec518f661214d6622b1502278a9c103bcb76aaff78af8e2f046234f4cf30d832a5ed43403ad4665358e9ca1450d358cf13c14bc7d2ea37d9e44348e1d0752418c15b059551720c52afc0072395fbe7663ffe4416f6f1cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h804c3fe95960c1248a63528084d836351a049a34993071fb7f73e5749a533f0e46e3491f803cd0b5580b433285446028ae27dfeec8deec022bed75bd75edede08e2caa399523250e6f55ab396703cdde96449fe483c0aec0abdf08f2156f55ff74b23efae74b4b47d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb98b4a68fe506bae383fbe07a056e31021a37980e79c905d7ec42c42e7024c73b57a3ce1834ee529a2863e63732174cce74cda29323d59014d1dee4f3b37fb34e9bd44f4ebbf212d72634832b763aa373444b0fe78550f433ae98cdd19b923d20b55823da3f9d6fd92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e90ffa28b89edceb720ec53a29cc96f6aa2c7f111ca227a3d50e2a248e9b021919e85c010cbc253f64b627794e0701df1bf87e66bbbab1fd37b9c0aa30cd80111f69ab081dd16fdb67b6a1f37dd2a8ae9ff602240afa6da1c699faeeea37c644669624ed629d86b92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0ef6faca9664250c5cc19bd6c35c5db47d481ac61a1630a0f8985522163866d115e806236078bf159f53159e7636a9de35fc3c7a4bce1757da1536a07c850b8f6cad040253bb34b7a9cab0ba8a6ec40763e737a2a370345ad543654510a89b050b8e0d370e632de95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1173b414421bbd50f0b3820a443dfe46ffdf5a2d0dcd6dff30e4efbb0ad5183cdfd3f3f5d9331cab0fe1a1d2875d30cd3243b47c89e4e888df376b1b7b59095ec50bdbb8ead2598aa5d8542a8564ec21ddcb237cccf4c94b640a695feb28c88ec322b8faeb7313cb78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe97096306bb3228294087ed0ca32654f46fd9c850016b5276bb3f2f32d1408a6a43a2f072e3038afde5d1892fb414d56d00df2a8fb678e9e49ab5d6d5e4b3fbef47e05ec7c1d8adb54f2d92e8c1b0ecf2c96f14f51a51ef41b5486e1516d01abb0e47760b7a8f72b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb079a60b053eca63f8c6891c045370131eb6ff79bdf39ca1d29f361dec2694b4c3a2bececb636b1ad0bc037bf8b970cf980f2fb1149027bc0f1ed8152c7d0817f689772d5e6773330b52b020b81b3a47be1779cf5dac3044984fa5962f7bea9c07d87508f9d2a9f4ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12923e05f7c71884088a03e69c6f8e5492127142dc2526eb8949aab134514220d4a48927249deeacf215bdca21e8ced1a48954301d1f1c9e68796dfb1258bd280bfec6c5c84ddae2dbd2521252989a1ed5dd6fbe6dc81d1a7d6ea747c32b826d0842d399004358198ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83091b032dc47e09020e209cc985c996b6a4581faeccbc6ab02404cbb7362b4312437e48c8e79f2f9e213a26d32a8844b273f7d842dd5115acaeaa27b0b2b5c0dd917a861121c7322fdbd374f824d2cd849f10cdc74743a5338a13692f66f31bc7f7cdacf9970106da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a841f9cae0844be579892d3a0c5b2db6253a2b860bdf406ff02a98363a6bebdf29085f64697e2f667bdd133873ba6cefba06059c3f0585bd55bd6d0b3cb1c1980efb95273fd81a9896b75d5909d1c1f623d6a98f4d39b6c9a0d2cc61b198a71b89196c74491864c36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7856819b6a6c7f9fe9c53f7d8335bba83d60c836e009b77c23aebff86bee6781c394c52616eb5c1d400d2b2a813d82f89e3714372726e2ef1463a509334f031438d36b611ec668097bd54caef1e4aadcb8819715e4f1cfcc6d8f503da314ab6b3f0048dca098cb739;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110d76f94d0213d5d79bc121451bfe1285e577614f5314f3bd9ea9789294adaa6176ccee67dd5607aad0e154d1de0f9a76e0179547ca6adc86b0843f904334dc22a037b1d25a33dc9e919d595a40a91c8c1644fd432e7e21e7815daf94bd6a61068b221a8f69dc96fd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19eb651725b5323bcc7b489d5ffda69e0165e766ceef5aaf3c8cbe7df7754387721689470ab36381244e8625a691b4c3f9f68fb3b0510f24978fbb8b25144148cd3ac7b1ddddd0a668220cb34107f74dd02bef65aff58ffe7eb6e6a8659f2d6aa6acd90bfa90bb3e565;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a35e65338cf53913610610beb1945a660e046ff145e6509788716bf01b58215aee910b7f7f93befe043e51651f51dfcb227b21e7d3d5cc212679696129b44f1fcefd117ab08250bb14741d771c4d6c04a466e9ff344737dd27812c0f3adf26f3260ad2c9b34532771f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1b4b232f1f25286c3307027f8506aac0ce4da26e50c5802918a15fce2d81bd64559721be698f1e47d7a233d2072d9f1c43c7d234426cfd0aaee96b1d02c68a77e3de2c3a62d35806a00455ab1563dd1dda3e6a0c4130fc8d0b26c4cff80128e7cf1d3840600ddc00b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf5a4c460626125c56248d4c50b6eb0113fcaa0feba6f96bc7a7e6f1a71312503c35ba38acc6d3cfd2cf8d1f3eec887cbd3cd994326fe8607a04c67c14e78e0844082891b898f004f52535965b7b10ebd9c471363343787b2db5117e3f52c1f9688cd250b86b14b624;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ef82ce44878c727b9f41276ae168dd4c3c8da5037bd1c3902afbd63e8379385d8a5720eb417a725be46ed09f00fb3b18e1dd7e93d193171977ea33d3f57406c09ad818dbd7656cfcbd2b070c4bd80947861f8a4c6ec1e47d5b5de17b2302ef6177f224502e0c83887;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7c17bf6412d3b591474ca2fbe6249b7f7031da841e1c5dcc8d9ec0d89f82156e69046a5fb5247603189ad1f109e05a2887ac6a5a3202bad9dc14de5d2719ca31ec8d85f804dfc54d9da9fc17d7548e1a47ba7e1200364445485cb49aea147218d997bfda2b16fba9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha899978c37ca453f2d00090106aaff384551eab43b1ea7183673be1c0bdd09a19c6efa2630391bc2de56d4d47c89e767f355c9f4e9cf31ac13ecdd421cb7f92241075c7140d576a973174e83634f368c793764d094fc7c66148a38cd640f1064663ff5c0be706f8c32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ecffb476e18c8f5b27233f768d7a03f3556ea42f42aadcbed78e2cdd413b75a4a476abfc16d16e4ff0f56b817b9ff337239266fb66c3f5d6cf20376a901b85b53c4a1c28a28f4823d9e1515cfd267797030806ab734fc48eee122f434d1646561c7db6bb1d2c8959;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d858db188caa8f6bfdda0b2fa88e370abfdd8fcbc771c82ce3a38d45a73646007ea2ddd41d9f9c29ad818f457d0e9b564b2eecf56ac030aa049217c13769e23c5390bb82c408e1f5705125f4cfa1cbf875663ffce6ae2182740cd657862cc9ac07aeecd23ec447a80f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45e61bda076cfdafb1f16ca930978a9fe48eb2edc6831dc0ca16c4a31436a335e42cf5ee3ea2a99c48bf235209ecc39d0deaf1db9874af5439f8fc601adcad05be5d77d79d60e0dd6feeb9ffbc6516a965c324b31bcd805656f661a0fd63951baa86dca9a6486cdc22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162b5f3d1b0efa54acd97fd6e0df20b0e17dad5b16eeb059714c07cd55bdbb728c44f5afb54549ad93b71354bb90a75b29ad2f1698a1fda8d8775fd28e7fa3353dceba9b381d37c0903bec1e6b49166f96c05b607f908405e638abdb2396b754e915d499720e5bea324;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb876f254c096cc3649ac21f3aba22607893dd96c86f01f8b7d3381e2da92d258beccf3b11911ac31e4d7df496f5da71de2c5d582e2aca84d14ba4d0ce2c7cf126a2fcec5d42bfed5bb2dba5d7ba30ce72a193b88ca18f4d16522f7f9331d6a0c42e785edaa7ae021a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17572ecd9250013af76579522b125bd5964ef1298b1abbbf3d9903b0c0377942860c607c3ae64e3c2c8c8058ef2d428a2c1a7fa112873d71fc954131abd1c3c5dbb9053fda1e484416ab7111fbae7638937d4f6f7753e2242c227bfb2af7e75ff82dc45147cb08d1df3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd8f58cd864c1bb0ea062e22e411909e1268215bdc8155df5d36c81c10d16d0c6142e4047e232bb95185b13033646b06b757034b1f1f6858f4a4c873e3501d2f7b357dc8cf1fc316941e8c715048b778770e1dd3c9a6fe93d25098a6fde51a95a510beb5d657ad8a53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8373c91334fab55dd16571ff36b51e16787ec861faf91c077dd4fd8cdbc78de5bcb91d5e30c1c067ee4c3ac5296d8c59f71b9e0ca22e5dded57afd4a034f32dc7e84e787d13ed9e820b7231cd7d917f29f3608de7e6a8e93d14ed1b347f4562cd655fc1fc95db0cccd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101c63e57abcb4467b19e1dc1cc56d1258280b1edaac07307b98a33c840ae5479dff101abf19829e2a2e5eaa7f8b0d7e503c2303c5ec4c491d76843455d41b1b330d28d05c01e9c6c6acc8920e5d75851bb64da77d6b441c2c17422b0ae91ced62ebc5773a7e2abc7b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e10f338fb3ae42365cf7a5ecc025b8ac219a21867e849ca9945b9abfa51afb8c4665b4cd521e2627a36e0075a95f60b5e4be27a22d696d79c99460f31d57f6a6afec9199687c010d0a62f3b8747c5a7fd1c8f6ba6636021babe8683b37c55834b4b5b334c611e2670;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8ff3784a62100acb7c727fc63b348de32970c5543f9b7e17b36d274e1c9ac4f0b0c5e11a0135c0ff10cb889fd567657b4dc7f17b8fdf45571632aad5cd52e0ce2b337a73a23f0500427dae74bde28041ae711a17515b03fe0700ee481044fba0bfeb3386865949bfc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca94b85572e0c6915c9ec0e740c61a801febda8c04d47ae686d8eafc839e41fe95989c2e5e4ccd75dcb46e7b4c0010cdc6c4ad59284fc0883ed2af6652bb8ba8cd8173dcc8544178df4598f5c33eaa790954d4e0c095c4eba492f06985b8bee299f9bad523e2d92652;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha77b091f969452b6edfdeb97fa7290ed34dbd5aac49b8088fd74cc26f5ea43b91b8f87645341446517d953a6fa799502128a094ab54578752d574a60499705a110706bb96b08837e9f35c328f3a891a0efe31298fe51b07d5de54f44879194780e9f074d164ac9a814;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6cd1be30fd60c8cc78ab39c8783cf686bfc0073305e1741e2dfa05acf68bfd651f44f0f4a601a9ee75970bb051b81c231ee01df6adf370a47a31155b0d869ee37b924c9471c38abebaa063c53ef9a112ced63a82122948c65e8bcd8ea1f5d72be524080a071bb3e9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a920c961f432431f2221200b2204935dc7e435437050bd97f2966bb6bdd9a2a97ff387de05b1218e4c78d7092de7f5ed61bfce4223a29488b4077d9c72f9dc06a80edae4020d0b2bfd81f2c267de601aaf76ae52ebc227fd480cbf27cae5530caabdacfc0e8abd91a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h885c522b90424e37231ce5855c636d1dfea4cc3e7b35a7724379216bf7f13cb25ee6ea6d5b084f86637cb11b33f5d100d5e8b1266a7bf99ab4351b0eb983c014cfa9c3cfc23596e614b0c25d03b5b1c8b35448afda9d6d94b0820c253e68050343ed6e91b7946eead6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118b352fe097208293968db87f6b378d81ed58304f7b480d3d349fe6b5e02ab6198a44ab4297046a70e7b2d8b5896b641ae35a44fd7153e6fc2717f076313977914887dd6fca8299799829c443a9b4634246638f795a12d2e1c00d1227b4fa4f34de471fa3b5844f915;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h266faf993c78639b14154e6a2c8c4b9782456a0cd03e3a49ab326e72fc3244f384e57a5e624c21d7ffbe0c3a6139b88c9e7f6bcef3a32f5ad3127eb156f38fc33533a72ba5afdafed1b2e03992ed5fcc2dfc7582c6107881af25a0721b4f76a994280cd593188252aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57af6692598cfc046868102ee2a9af7611f56fab94dc0c325c23fc50d1ebd6c722cbf9da1df7d7c3b1f4bf31df61188085e02ed51cdd8ebb5b5d7442728611c93aecd93bb8071f2353367503111448410aea10aacaaf71913c0792e17b1c7878330f8cbfc97ded6005;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac257f394a85140485f55027edb68e3f184ff05d3674fdfa6d60f66697ed26173ea9d386e035382dca6d98513059aadb59ca028ca1d6f6850d328a5465134a3f30831e77c72468ad342388267d9a5c3f05a678a8d2e20a5b1a1165f1d62ad53e45accaebc49d73f91f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c1479591e4522e1d093769c1321a0b408a2ae1ff00beb96118a359951b9c08fc94cae8c41efab54a97176984c3405206db947b6ee953e6f2bf42667e67e7a04a01f55841ef8b3cb49d39ecb8b31a73d02efba4dee4c92047c1404b49d655c40248712db7685bf1fbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c00f65d15549d2d2c265a23cd08e4fec38abc7f1aa5e3e18e210c871ac1f4aed602c0a4e3bedf9e4d0a4e3041f1e8a787a01fd282829fd200f341289a7ccc6a4cf8efed51d4a5db541c7d2b94d17027428d9a38f3d4cdc9649e6be928f3b8fefae473e7ed0c69da3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1effa25df80080678b025b33a5c7feef694e5d9c038ff2f74985eac94e4f3b9552b45826f2ebdb21fb1d520bbd8dc306aae9c8f48046c4edfcb89adf36b53deafe7417ae99badc69decf2a6a125d8b6f097d683b7bfe4a234d638107485328c908d1f459a748c803c9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h288018ba7b1dd9d4637bedbe69a6d69552a67755f550698df064b67384601a3642a6096ca3770fa59a15d6e170f1090a4d3f58e2bd9ab5f1969bb210dd5424fe9f6a45be714649820c17cdbd7860ca153a12c21d3eacf9fc77699300ab730772f53b8bc06ae256137b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14078798612f2efcbc5b8131c7e6baac07f8ccd49120ea5096a8b65674c2db0d4e1667024e026937df9865b809bd427fdb67620ca4d4b20f8feace71a61303a6956b516d62bdf314814c27136b2562e8830a9f3e68f8fb2ba401c890ea03626188a80e7ae857fa2aea2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h488a5191f90e1884a97abf9760a8ec2853c5cf2e722a9f8ae4076d580d8a40c1d364212121fcfd81bcb2e0de886f92a99c64f284f4e4e580abf2840e9dbc36589ece5f4371f5add844f13e5de24817e9538afd81dc3561c82e11f404d97fd4bfe04a5af9d4ee1159ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e4d73b68c5c2093fd38bf441a543be65240335c03fddaa5fbfe946e4157b283111f24b3f5414144df61265f5de413446917e445e885f08b06a0a5a9cecd7dad2cb65b24e769108560f6fbafc89e8d8f2579970c4e4534d0d3e8bf0c497050b4194d38c995c15875f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c5ba5fd5695c412492477c051d6268c7094ee67f4f0e2bfb77125f3c45b05b1a50aab45ea2a550a91002351c301de0f62ff04643b5b7db5c8296eab838e04f94af47410cd06f659f5fca209cf851590df7dcd5893e0a01c482d862b9141a239ca12ea739aa22ea259;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7792719ad29e8e202e58116c04ce9f5206b82bdb34ebaa38fb18459b564d865239d0d1b01a773bacd3425103e7bd229265ff1dc4632c0bc90aae562866671817d318f6220ca6d4dceea5cb2a90f843e7a9a459776ea009106cf16d6e457f7e2310210039a2a1a8c4f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha012554ce3a5a8d116430908a2415b9982a9123b7b0e4dae03a88bfe8814a8db44c3954b0b9fcd98ee771d3530412b73aea1b77824b3e0962e310f859a25e73fdfbe0774e4dc33468faf4b019de11b31a469775830b7dce83e6d8de7ee63f122940f05d90f50d7fcf5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h583efd8468a0720ff9891187d0586135d9dbd08d10f7671f839dbe54facba34ebcba643c67eecea0708dccf1a63b41a7e33ea3e4f2427f139b7445f972f9930740f29aa195c234b1e0d38afc25b98bab77538862451eee6700f55bf919c574b22c2460f11b2a163633;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hefd099963112b14bb173c3dfa4abc2c19fa1c52463776146a870d97f241703caae3b541f6459ed518884990808f257eb316672b9a1a0c354df0f65cab5f1d7e99abb829716b04f38e5d17e2ebbd996d2ae94cc512b89af409be3298911c467dabb6619efa7c2ff8db9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h247d50115df4af634c9a7047270cfbd0865d020f17023006a7231f768cc698e34ad011607c22f645044c134034096156f06b8bdbaac62af6925639f4dc0098fbde333e4ec62ec528b89fa4540fb2dbcb4532572a604be9e2122c3e659253cae4fd34d322d22c29d710;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd93c8ea43280ccd57f65409f052732bec29f6cb1450ad4d27d4d356852ad576f1f49ff624be7c4fce8a620e7f5fa8ae0ca51da724bb68338be315c3203075eb04abe22227db7197d338e534be85fd2df1a099e5b72749f73793f1823518cc542f980a4c11bd2e5b85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db5c2b8fd986c00888353ba9a3cc7c2ae4ebe0632b248939da0f929bcc57eee154cfae0f24a20924f10cef7a4d6720dfa3bbd09303bcee1bb43bf822ab8823177add092fea0967d9efd58971f823c2679e08c177d4f2aeed9923203cdd8ae595340699b3807ae594ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h954046599892b648bd37fd79241bff09be9aa01b51b9464df5f1c0afc2da709103fe98cbf674a253ee460a00a77ffbbd73a3095be13f2379558db8ab8ea8c205f42637b43b5508e2c4944c530703d3c71c102408642da5e9e3d4c5eecd762aa591a2e9516ae331c29c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf9768821c134b83a257f1eae72564425de57e41d1a776d1392beaec2e4371e6c189d6c8da20d2cbf05501ace032eaa2a5617876d5c44d45701f1c51e3d065268d8b1a7a408869f380e32480a00391ad0118e1914cb18a209b3e4362c79b93d699411aa2f12d2d33d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d948aec8c09e9d7996f0000474061bbd32cfb8f585fdcbe7eede5b93300e11465b655009405c619652586eee73b9f2a60cf83b9d2c476650fde108b7fa201039fa44877bd42a7288038aac2de59e051aaa7d6b0fc93be6f077587fb2a78e340e4af52d9eda460d388;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a142f533d031d2ebfa3662d743b39c84b7f6a90018f29b563b6dd4101ae947c8d91ad4b13c5b860d770cfebaf36288fb6db9b527dea24ccef9f0c56b47527c99afb8597944a69d48c6981c3b9de73d81ea0b6df0d168e4573042f9a46fa3e4ed937d81cadc87734333;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha82e9641c27dc8d0e4fdc4025ba05a82c23551e3a6a36ef7b5cdd9b6dcb13a435f4e619df6476a483e0a8a869400ab172175a502ce561d233a76f495a0c515ab3ce9da47d49c56c73bf195f2aaaaa70242d8ea84508c560bd5d5e85117d8efc613bacbb2058ae1a207;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa2e2236e2b170fc271323def6b832dfbfb697cc49c8c20d05b6a0bfd44126276f0a25f0beaa8613f983b589340aea4260ec79ff4e620498e5abbfa2f386098c0765e710794155830ae2e94949a487c30b0865be693c30212dd094cb6586e59d5ead4d623ace6df33c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114b3df5bb63737869b2e113b15eb57296219d95e3d593bcbc5de75a6e425b31a445a4e858f40d56b75cb19b69acb7638e2611b4221b188eaada3e00a99a68e643d369bc2cfbb7aacfcccf0fc191fe7474fdbeef15d0d2ff443d248cd7cd2c9f13cd154b51990f6288;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd49f630c64bbf2ca9ec9e7fa63b978781d1faedececedfc8dcd31f94b877c1497833f5c9b9304fe4003ee947ce5726a3492a29e9cd4469c8ac8fec8078a715ef119494e29c3a3a93b31710c1b21bfd7282936b507e3cafb59679526b3caf5def0a0c8d9b17c0cfe92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1d08512b5bbfcaa94c5d109317e287c0fd62d1a736fad05e5d50859522a041790cdc4337018a45ebfc082376163a051417cfe4754b4e6f83a1e0fd366faa42d07a3ad593cda88f8decc6fb46f2319d7751136913c0f7e5e5f09718b60d2866fefcb2b477fa0e35b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha227ff47e81bf46716fe6b26e3b637f0e08a23ddd048970ce22c2c5cde4fa376e2bb8da2524cb5808336acc9308df7ccb76ee979638cb62304e4c862a810f6b14ef76e0672447b2bb0c3ec07fa114f5a4be0d1f1c878b46415991feec92d1a055062e2013ea1945ea5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83bca626f391bcfd6a92db1ccc0b9153433372db997dd1347cff166f90868172d542881c5b431ddd06e41ebf5a9f1419f992bacd13521fde403a8f9e9abe42140b15cb49b63807220b6d11590c23531e8a77ddd6542938b04ffa617003035826d930b4d9e471d5eb8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f657028b7202da6d6662a41aa1f16ad19ef133b23d39002fc90e489152adc17d142db66927377ce8774faaaf10fb4297077bf3b530b15f39de0b7fbe5f5ef71f553b4537321941a53555c18cdf1a9b08590d16a57ce1587a5ba2aea150da711800a6c221df578ef51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16218e9aff4a4364d572c184fbd5d373c9febe7ec26ace865187ebc1574080ba8e926a44dcac48bce21ce8256dc22360b929648e40f98f0ac9b0b8edddd35cf74757d0f40730f1dc8f7e51b4bf3bd0009ce92b8a8c5e6039f32efe14ab3316dfd7223549988e7175d56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a7bd48856b45b59ece502d79135a085426135c1cde353b0e25bca5549e7c7d544752dccfff5f3137c559a0814ef933e7010649bdeec76a556849c4f2c38416ad4f5eeefefa4ee3a5ef1a652d1728827fd3c44e6247c7bf89ebdef69672f4ab07615f6ee0675c0d5bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103e2345d2d4f4f05edda3fca59fc80990dbf32d701e55cfae8f033b0a63a028c8750e62e11f9a4a9db61a51a682d301521cdc4f949f8e36a584bcc05152f6f03b05efe4257b23a4d5d427efb846cd389c5a893d4b3d60196ce5d0eef8236551b126d06303cd49fd368;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1335a902a6947a82d460fb440ee30c89d053aae4946bedf5dca3d2bbe95be1ae2d0bb12849edc5764cfa43cb73383a58b1813474da61bb595f09402af72dba6f77a219d64b738ed8a1467fc5dff58ac37911f1ad843d1a26cce2cb129f88830c5b5bd9d5f266bdef5d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3f1c88fa573cdbf6a7f1ee065605bcf5a65ea51180ad1fa44f83b0fb14330145cb43466e892fff95f56adbd5b235a3789ce7eb682353bdd87f527c9d14c0c9f652f74597d43209ea4481dd3f02fec07a8a7cee81a67907dcbe7133ccd7328c3be41d8d35c579c4b51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf0e4c5b26bc5606c138f1d5d1fcf963e962055c86ea3b57096ab8de35f74dfbc80a6d41a7ad6ab1830d1985773efda527f62a4f7b301fd6caa03f1c93e6d91fefd7e7bfd958182ba06d1acb016139c2b5841afcafb4b846516216d1c5b2a19e9592ee617b226b2f1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8f0cd08d32045c93d9c36dcaf9b9381ee1dcc191abb807258aace5bb8965716544fb0767f82a5a7e638521a09a2365833508b103603b98af64cebd9c76b98970ff22aef30b3696323e42ca5b4b9c6fcf5619dc55c65c2f0c3501b7b0858750a0ec8706da0f89cfd76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heeb65aa4675ab017207a1150999139206728550f45a8b4d910d57acf1252fbe8f7a20597f17ea464d1a9cbf787e954088c61f18ed9863103f2d7ab977ca26f384962ddccf4e773b18117d1234e06225bf9d628d225bf9afe76229069462d18bdc98e73e5ec2b0733c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4b72c77f7dfc8fd122ff0f2eaa28b5ec0ece37b6f7c34e6d29e69ec795c5ac560a3312add71a84a6ee5c7f05eabccf85db1504a80d5f69774fe2026fb2943357a57903c9291c0e7fb3b6005d8320e0b4b619ed11779c0f34817bb01ff478c6d96b39c0cedcad7a9bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e3261ded541beaca27fb72dd0c58894bf1f14f35efe258604c931b271899d15ea0563005955fe93374a3da79883933bf6858e072517f9ccd6d2f745b73d077e4c1b1a967eaa47199278a130e2288f89ffd534dcc35958f7d801ec081256ad141dca1e4badc2d5fb3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8eed8b598da45ec9591cfca946c6afcfe5e8d4af0399830ee400379704da76f7e37b39be83e11eff089017efb310558e0bb6acebc6690642b051ac47e60c9d98a313d6f1d03e75eac152be0e68a978a0348848b02d1a5729ed141176ff1c74d3c9db304f1a83ab45f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159374cce53b9edd8b02f59b01bf3678143d13e3b0bcdf8b00e7610f282dc01395e23018ddf744a3ffa2067b29ed726f8874f5ce1f5d9f0a2821e2fad85e1b156a5818aa386fe4df441a183997ab5b95874050478a725fbc4f2a08968ea698261660594f46f6308efe0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba7641599d4d6c0dba77075ecb5731a34574f37e329683451c1f38ff844fa6f04a68423541862a787c91c8e554f22c23eb735e68b52cac7305d5692f949884000f406fea41d328a8ac14712c1ec4a39b56eb74894beb2d795a894ab7e6218b79febdfe48b1d7e3dbfc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70813af7763a3a772016945b276b9a53f9981ef39346666bbcb4351401fdabe3c951b21ea6ad7c1b83f21f065d6ba976bcfa92599c21fcacfefafbc2fedeb5c33e5db02f1c6a670ab5bfa38e1dc38251309d8d96eb3735d4c1ced9aa71aa21df76c41cec106d5f33a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bad0634171c5cebcc21efa1426f794a77f1d43e34707ef187288f5c2fd8ecec7491fe1633b5c4685f1fa6500cf3df204bb2cb38a1df25f44eb3ecb88e0094b9eb8789d29c6017811aa58789912b7b66f56e517f39585d6d10464f81bef48f9b3f5d4cf8954d7cb2562;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce0a970b50555cddd120a85f8722b35f025a00c5206e44bf11089c9d0bb3a9d89b968871b369ce0b14491d84a1cadcf3687a45105284c9e7ccb0cff5c353d235465c965d0f9c3ffd7ab6c6ec9426036e434a0ff6b91b4c67911717044b0b96695c186fbeea216bbaab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c426bca85685787d822dfa0f836d6b28ae44982c40cb173c9f4f35f15e8e9c8994cf98e5c9ce9e1fa7271f6de778ca50fa1025843d56e4aaba59adf149583b7c030c64109840d23a4a14155575c17c6e25b8764a60fc4360bcd9f4fb7fa86c32c9ec215091e7bc79d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196ea180b3a736d8587493f6da243ad379766a16e55e17bf183f0f0854e2dc0c395fc91f23ca157fb5090f543f2f97f6b6ff99f12434b1cb849ffeba6a5000ff60f7ce77a0ec42ff8889215d1ade5779f71566d1481a4b3967d4da6399b3b8d19515658fff4d9de0a91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16280dde8d9a6cbb5debaa1e29ab29f1666e7d62688e8a756195938918a1728e57efb773606b6e3e77b38ccaab2c721ed7377c9e58af3658c1c725532c092a1e9a4dadf0d4cea4f65adb52a71178abbca9750ada1b4514774c60756f4a7533391787d76b243c0d794b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ee1dd22ef692707fd512eb380a318472cc2cb751cdc545229f1fff0227bdbe2966b4951613157e4233989d0cc08cda1a3c4f37a5cec68336946752ce72435aef2480ba42a0dc3da8ee6e55403e565b77657bf5b776589e765798eab3e373ff07363deb806969096b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8490b93a5669fca15edd2d16f84482b0627e52668e881d6eaed1e49e1c9846564f388b51b58202498054132c03bd403616ec89646f6a9d806aa6376e9465fd7e9ede7a4150a28ac7abeb7be5bd8790986462d815ee79b0c8a3bd746bb9c1b4da0bbc2da3c239b6dde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61678ab4c9053888071d539eeead049abc0e9143d23bd75d379cd05b4f20e3aa379c1777b77a848cb1c61b09084dfbf3d25bb2fc1c434e357838ec8ba7eded3feb8af427cf7227cd947eaf4051ff65011753e84e8c90ffb27e26dda055baccb6cf7475845728f739aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc8bc627874dd8aafcdef57cdc34f2fca6921c1a5f5e5e2c952d5827b127416acc5cd720ce5e65ba10b17156ab3af48cc29c12de243e0bf59cc464f04646e091511c2733f2bb129dcc0ac09cf458c7979e7b77313f6968f21d2dd6cfbcc8ca0027b1882be990ac8215;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151ffa159f59625c816059cb70a66e92e213d7ad75d22adbd8faf84ce1598d907f80fbdb3b7a06cb323f6b0644e6427b96f188ff5d15606b0e1de7196146109fd7fced6211f19ddd4d99400b10d2e310a3f899884b68e3eb4d45fcb645403bb948cfe9981b4c162bc1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e7f6a30ecae010fe4d0e3bfa0a432dc8758d1528196d3d47a05a9aa9259785290bf9d7d4bbb48822477c0472f5e2bd5280d54ff2729a3d8f414535bb8386ea00295286dc97fe47c324d4372e0b5c0a453cb8e0e393b0ff14a29299c33ae8ebeb90e98474d115b2d72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a999eefae58b4127bcb82b628646aa3a506bae33939a4b938083a6c4e6b90a8b9d5c72b3380ed0e1d6d8a6c99a9006e731aff22b7d8ed68240ee1b902dbfe157047be3ee1a4e461ef82f5ce655e7382b45e25127bbd86d9b5dfb507884ed6fe930fda8c85ed94488;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbb8fe9cfabbb480401f93b72b6bd05244ec32b0c599c3e46fd015ec2ab75ccea4d0602d19316bdd0933fa663050b9e915a11505332683e5a6eb5c70f8b2656a34d784fc15b0d08fd071d57f9b240c313dc02cb7efbc31a2ca429be78989df58ae08a4005138185ee9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fcf647762f8632d77ffa5cb534afab71bc9f6b9282f53fb61c28a8ff8c8293ce9ecc16322cd1a77b9db1b1d06260f684b8d0265e801aab957747b4e5a09f5d2fe92c7d61c35a6da40f9a9a48ff34f0a4cd94a54287215cd278baf90ee0f49bb1e47375f699e20589f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17288346d9a00d13301e7263d74e6bf104cdb1dcefbc2cc021ec86bd1dd111fae077d43766f95036346b23925a00401443b07af40c0ac6eb9d131bf62e2978f700b41bd4e6a4cdd4a987a73cf3ae1ff87f19503732b37c1999d1d5672b540ce220497afec840ad206cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e70dcd33b73257a30a0b51da00e4742405c4a64c2879bbc1210b5342cf4bd17d799d04915bdcf8272dd8af063c4569291dd7d37d810689bc188bc8ba3400c87f767eed5f975746e521c450a0e1044f4c68922b7a8eca162f386c803f75c8056bf2e15eb0028176684;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146010de34a7702c97ba3b043dede911bfa721750ee4e2a0f80292b74bbc361437e7976ff8affd15c95742fd9b08a3f7fc5d2d4ad38d6fb95382156ed86f8d7537631510d1510864f9f2ffcbbf1b831850d250ce27598af09d8e5972d0bbda5613077fb667bf2c3735a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87bee5379a0127562b65e9431265a3a1a84487b49839f5f25bacd65687c4b58302a3015b9940c0f977ae56b0d263b51a8c899157ec5487540522d9649490e53582c0c1e9f360fa72edf8a8679e6e3f3446f8709d48fcf94eac30c8660c4a8818f86f5ee840a907305;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136b5d08a570151c75eac809b406069ad3c85d9c279318cef2b34d235390b81e2759fa946a718ad308b019bb66c7e511300e24f904703805a7800cd9efc5135988c37241dfd0599ef68af2a5101d3bacbbcd4690d208a64d6c9e081943f720b51b88f0cf21a5109dfb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163ec18011560865c3c9a45c7b81976b8a0281c1fd1cb402205a0a5660602ae7b5d7fdfb61715eaa3ab46c0b45d337fabe3079cd2871a5feaed041b33abf18d03036a23026c71227393660771f6c42d49e5cf60e3052bc92f3e12bd0ecfc21ee2f9720f48e67849106a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10575264e7a440d1090d3089bea226f84c5d698e809ade889eaa22a7f904603e8e59f0f46311897db6f7e4703601fd07cc1ae7ecf1e961509b3c70330cc27111da94340f564b82fb1449b628a9152bf7fd5f6f350ada31011a65f6146f188e5544dc3fa531a39806b0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf0ba3c6fd93b67cafdb98c8a1db62819693049a6717992e5200d9ab5a9767c7ccb7cc14aaab7344137480b9e4a3f46422e48a1e02946f594e1fa6dd627521dc8ea6603aa809d569879faf604029f85044e66acefa836c2afdad2fc0f7079730cf5578496f5de3d2e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127efce5429bb2a97e55b3f033e7f7ca70264ea66e096d6848cfe6437185c35c0b25b785e44ca07f159ea6ba47025ccabb5213b4b5edaf7c1600a7b0a368ffaa6fc965b7ad5b715700c4f2cf78b90836fcaf365a4469a59ccf4e76597e7c7ee035d3155ae35feac2bdd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heaab77444619c508006e5b37010f17f5a74ce4e98e96e13025d497e377905ed009f5a494291f5a4556e59302daa298000c0c6408f907932ade3f8c186113fe3dfc6c5e8d74d79a8beb0aef183f401c6eecbf00b5f19336d37db2d6b3627bdec26f1260c0316fbcd76a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cb54318ade5fb7582080cdb501a66c186a605e2daf89439d58b2c19a94818434669efe5a853dc1f844402f29605dc41caf82708a8540b345cca21546c0d36f3af491b8959aa05683bdee54a0b26aa08de4b532afdd63411a53b37911b72291492283d6039f68b0618;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb450c99bfac3e1808938a1bfb7c13357e86177e2ad0a79c6a22575ff3fb0cba1b3378e9bcb3cce8e68ff0a48d8341b5da29cd521bf3c22b2790a21938c6f836b078d573439b1cac9e769de4adc24fab91c3c905c4e12473713ce0a851f30c38590f1c2dc7bf0c694d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac51ade411d1b4fa44fd563dbdede0c4294ad4ef44a48781635c77c4ab7fd2d030e054698662c7030ff14dd86242ba354021781f032a80d3c56fd48ff1a5e5ec2e33a4db8535ed4a81cf34bbf85f0d79bed797723c4b96d671eb39b9e47a46758ab4c4609f16d72dde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5a68ea4920bfff7deec8b7d1f9f52ef405e8bac5f77d07b4bef757cb1a73aa2f0d570bed24eca8c78068f1700829aefa47b65678cdaebd47bdf0467f649a450dde67134b6e7f322106a6608168f64b12cd9148bc829dd94697ca0e6f0a5b0ca82375ade04a0951862;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4837dd036136a3185e783677255733c6a8644eea608b82adf042ecbd1096cc0803a8488f65f5378ebe9030c3e806c15e4d5e06d647976b9492da1cd211064f3e73beab6771a694c4278dfe306a1b44afef6906375096459d49c697664bea7bd2b72452b5e6e0c19b88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18cc6902baff1927bf80431ffba564931bb5cd3c340f5a15b6190d2a844be5af04de2bfb6b6d650a72a8a78305c42cbadcfee447a34d912c8b24de88560d6ec10db3f4c8e088d3d2a89ca1d673748182bd71a30a1a0fc6820bc49a8739e5cd59617b9695fac4a3695d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142e33f64db7d84aee2033fbed46d5d93a7fdc948c22219973ae68bfdde65bac93b0852a6138751fc6ff2b50b2d63db9b4d4bcba8fd5b2e69af9a9247be10ebca6591857b78e3f2e3b36c5c2df63156780463da11b8df153669132200bf1115da7c392c68217adffe95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f6ac9a2032e0af9ec0b07b3227897bb19d5bd8e43f20786ad8fdb761111706b9acdd63d28a94e9d9d3109d1cb39b952af96bef28e1e685f6cca4a540a6c517f85aeebef56a113e0e875f1ef0fa6d70f8e3b0ecfdfeced000637cb4d838f55117bb2c07723390879;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113768c337b65ac82e5bc24f19958a91a27ae278ae7790fb04f0ee5a28675bcf27565b9c243a876e54c5cbdad96e2fc35bc95398b44f1a5ca57d0607229cfa572a145933032fa34e4a91d2b0384aa87e700da0837a838390376605db8198d6417316b950dcf194397aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192e303ad9be8b0b8a4ea55f5d2d5712f391db863d641738ee37afb7dc55a138f3311e4b47f597770b7bdfffae838ed0344cdc77ab0dfc7820459a389292aeae56d70493629993c4aa5973f1f833abb7b843454d2e45c5c2dd91e863c19e8c7074bdc559d547fd04ad3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99ff7b4017d2c86b34e19ac5892b6484425f9044861ed0225fb81d0913c347c31b39a0b31ea37fcdd607f550b267b209c195df9a2b78ea240cfdeb1d4c0996775a1f7c751a20e398014b7de30b65ddf63b1f2334e0a5979df3fd32285a3b98f22f8ea779c8c0b06518;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1637884c68d297224503a7b240d8290aa6877d7fc55de60b5d7978e0fa25974ca90a5f1debc6ff2e0fa78370302d650058a97452b7a6244a7e83fa521dee67b6cd71d7ce5108906a508cc967657ce13f005bb8d04cc501a5cc9aaca1ae1c68547b578344a9d4a4a8369;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118f62f1fca7cb63a8819d548d4343a8aa942585d675a69738f30f0250f652257839f202c957764c226a7b9373f82bdb7829d53d02420b8e40cca0d57d02b9e9895d25d04494d49bbce1d22cb9b1dfeb2aa0cf473b3e519afe74deb60b678c673b80fb4db7b76a8eac9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5efabe432a3053c9febe6eeb4cd2f33779e623ce8e46023634ed52add355e6d4663c3ecb0754d6ace82b5910ecf13d131826b8e36cb7cba0c543e4591fcc6b90c91d7f59cea9bad750a3224abc1a01c5721b32b24e067723b015e3539e520aec40539b03b49af215e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60a3c197a294bf5c6d06f70e8ee201060e660a157de049cd3f6f56062fe836667e997e4463bf76533fdd6dff3c50ed0618057e3b33d4afa6752c7271c9d791daadae10c0fa80aa7fa5e56c71440b6822c35198d2a0ba85335662106516ff00811dafde2ddadd539cdb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd864ac08a231e68ddb529a86f150b20df5781f7adb694a058c18763bd7f4290aacdcb2f8ee46f5061fc7da35fbceff93a02a8d887792f938956e5f397d46925b2ecf740103ac418ec3e07a7cc6de31f048440bf8cad2ea1568f115537ca1c3d42d564d438052adbc70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58dc48368cf9fdcea1a67cbfdd8f9cbfcfcbbc6cdad9fc38b6f146c8196c42ba47cd37da8a331a72d6c1609040f3497838fe750d7f7197f04b78e30bcb2925fec9604dc221d642ebf88e2e1346c01bcef9656535a70efa62e6e226f194d62cd22e894fc36966ed894a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b57c74e60719ef05059854124ceea8648895973746cb29942288ffc8e9eaa1ef2663b840c6088625b27f8d05431154926e8993ee380800b12b5d549a1af29ee5ea98e2f6c6e4cae811d5937d74277b13bca0386bbd9edd89625d8fb7be469f89f1396845dc448e4c36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a483cf8ec0927f664562481e4a154734a3568de66f148b1cb12af6c0632cb3fae36c5246f4c914730173638d979dbb6b9fe09a4e709f7e86fd1b89044b48dc7a673f5e863800f1cb6e24ff53f666e1f41a823c52e9557678b76a976efc107e8349e7e725dc24295d21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a3e8f61acecdb24f81f099be1d4067916bc62153fdaf20ad67f0616ef10b3754ac2ddf1c7f35edd620c1fd30b7b635407e06bb485255b6be53732405c80e867c574dcb0d16c4e35323c09ae1cf2d6c498e56c44651a9bffdde69c481b4745577d922c935679f1359a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2267ab6bd0348cd61963e1cb303d59ed68e75badaf685e5cc7575c4f5daab574492c2312a15ac13aada4942a932c0f43bbe3227185e3fd2a9e11ecbdca0bb9b8ae76f02ce8e082650d7f78458089e998a3baae0ddab7003689633ab67b28a0dcf03630d9622ac932a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h682f1590f862e4ba151d01bf866c6518525aa5ed7d25b27b81ea2d5c37a994a4c29507ee840d7bd4f78bd83fb46b2d1cf492ec252e6ad4fc5366c76a6089c0da37eb0f7d24ef26c27c4ce8147f8ab664e40a01643a1ac1396cb36c67b65282de0f74cd4219bcf6f090;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8db355b3b0fbce2828ec04743bc470080da6610ea4a054a5c3c12ade4e06dd2169f86130a4c8e08c4995ca10cb8143d23700af059076d4dfbf942a889339cba9497d1f213a4d2d782295ac9336cb8bb99706fa89c0258cd037988c19fe242b41f379a36935ab76274;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae9709954424218a347bc477fd2985392b6f6da4c21c25eab79417d882cb95e706af3d3aa7b57a9845b576af0646c05abb97dd0811183a0e924b4d5344b03d0758a9f978dad6aae9e3cd3dd8d1c08299dda06f1c2959d90bf8b6776cbed586343f294df1dd5196c96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1387f8dd0a27d486e78436aaa913642cb594eded31a1d060f4dc11786ef36d0f9444ac69528ca8f156082cda8b16262f31466b4f591f29de5c48602d38a2743d0a12c9b5f94bd1944e539c894de19fed3c3779fe2400d2588e3c3f7986673701bbcc47d9df52887321b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145acc7a99e29519269030ed433cb0bd4fc3ac19da3a07880df4422645ef150c332b778622ebc9d53660a9040a4850b080a75c72b25ad27cad8d26800a4c8977b0d348ae82661751b7149941674b00ccfa65d1cc07adfedfb1ced8c86de1fe2482b76f491e8827c1892;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c1938b6a446a6708bc622b95310fb1280f12b218ffbb07e16b4df79fd87c4909ae5ec7cd6d08327bdba148e306e0fe3b1a51df6a16eabd91e226b555d890fcdfb5c275b9b6ac5295db6edba8f6071d2b9fa0f5f0c9adc8fe321771b369f6c5316a1863ba9fd4ffc2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1509b976be08ca3b7bda608df164edd4756ea5e60f4ddda99f1302697942ca01ebdc773ba86768d018af11df6f6e927209a8dc0350a32e94046f27b9ae0dd3b002f352c12d290d98e39dab31bee98c5cd571bd557ab7e5cf8042d28266844dd2e3896d31e5d5c5ccf36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ae62d65e1bef459147e8686dbb9b2ed7a2264d18d392fdf2362f8079d3d33e0a32975e729ef061aeff748c24ac999b46ef73c797a6149fdb00893bb8083aabc1b7778d1720b433a05afbdbe6870ed8f984cb3e3b1afd6daa53771b09ba6c144c9b10837392cead6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac0ee0762232bc3d8a45d8b8d292fd3844014d1c0a1c476bd60fcc99bbcb888d439ba8371b8aff922e7125592efd43979425a8ed30c5d8ecf39b826f9d513c30b63067985ecf212258cc1f58a31c9e6ec83e12e6ba162196865377a4b488d6ff934927bafdddce25ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143bdd163204b4f2caa05bdb0433708d71e645551332a26860a5792a7eaff7217634005408de312a995329900dcfc91a00f964348e331bf034316b8d1881e132c4ae36875f021506c6df6dc31268852a46a76bac0cdbfff3066f33380bf436a28ff9d8b818d159aafce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha225460f627943dc327b8fdc3796f0fc3259f9649f37071fcdef6bfd91c8df46667f685958cf938c1a9f27a056326620ce49bc148ea6896b856c0e222bd70abf73669d7d5e75e54eb8d19df291b0ee9fca0dbeba6202bd7ecb92c865cae879dad5dd5e7c3585b56f15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6afae8542a736b736875766d503650563498b7ec563c5f4022f08504e38cd5ce8c8e05d72b861c1d87b1ec2df414da702f03ee0c5ca12aaa5c0875669e06a174a385f1edbed04b5dff3fb1b1278ec0c5188cc23992ae440258b7595f4f8bfd603989c3972f47e9b4cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bf0cfe15551f292dc9bae6a91b0f7ef69996f8cf0851c2af5a84699e8ad7ac5ac4d6b01357ff08009c0eaf9b2328dbbf337cfdd28cbab468642282ddc59b515991fdfeca426af1c6f41dcd4771722fdbb60b26eb1b07c4a92c458715435424593c6c16d0625c1f51b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb664784d9391ca71b4616a6c8c7d60033e141f2248bbde1e82dfb9b3e82cdd98edaf0340756f28637f789e810757244dc30d26a3091d40cb44eb1c6e2f833e87c6c03b582100631bd0f75eefea044cc0eb8c80a3dbf6e67e2e7e1c5bd77fb4e74a8b70b5b63fee349;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e924aa5cfc0890e357117c2cc7b6d450cd03f2b4cfda7cfc1d780ad809d364af6a4e8c5cbf3d8e02aa9b3d0aa6b8b5a48a66f5dc1071d136d8d489701f1711891d28fd2a104591f304fcd0c4f968d8f20a20df9e0264bd7c68573c962ed315388d41f0e59a0c160f05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c3344f2cbc5275a9724504bbaed53095491a28ca4e384bba9c914ca8547ed09644ac7c848de2061cacd7fd862ca950e0b5bba4fde3b598d3010ce3fc7d66aa68f7d2c42631803bb4f65f57463cdda06f9f79fd7f70c3000524e72cfe22c3add1e514c136de5576a46;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d2a06c4da92018d4a71041ea52681c0b4bc749690045687f0f61194ebf66f0b5b740b358430d6ba98ffb042cd53371a204f78a2500e808f787ea203264f4a699d7b2bc6f6b78da705bd1e65c7edb6654e652cf49363065f5f4548368b52b31cb004b27ca7ff5cc415;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ac16b87d7e8d6bb689910f05c79d21b8b4c627e5ec0e4b0b01f8af0e1547e822eb43ff4f4b1cd68c8e1c29609c8de544feeee7ae603641c43fb0359fb0fde96ffbe632e2c84d11fea82c7809d98866d72a46c63c4cf2bea6294426fb38520e3f49b14348ca1956dba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff4cb6d218299b5390473e558c837e33cb9ee3e76ec5a83dca229e74bf9cae79cb6ead3d543cc35d802e26fb170aec11dd8f4b1000f362c92064d09a0e10bfd795c108dcc3e267012ed1f8b68bf4d82c1885a93836e2a28fe5dfe28648e96bff0b63a9721e4ca325e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff9f6469d5ec231bbcb3e17429e2a4cb4efba30a157659164673b486f66868b529f1a0ab8219cc833b40b312f3ecf701b3c10f7402461b99b194293bdb44eb4b1f00b9549cafd75b5d2d3bb9eedbef238ef0bc97caabcd8e7061e39db3b71ecacdc015f028ae0a07c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f51377db39820a619345011e9e018fd00b2173730fa807a1e3fb6670f7524e0466cedcd735ecbb13945515a51df556bc2949f4c0e791c0c44b94a93a3446f5ac24093303ee56563edae6f75dbd5a4f885ed818de87c74e514ad09364b473e0f4115b807c31b04cbc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8c6527da0efb92416dde3d8b10b156f24200d33d549b133dde7971441ffb6ce579a8c74daf8f6a49e89b77665d6f6939f467301c49b4c7f94e4474295b55441d81d96e62e93d3c386c8fe13abd6fad923d45de47faee23d9c4314e6bf5719c7821d98b338a727dca1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h732ea802e6ea9df7c2161a50075ce222dec013d71b39cda7bc6f8e6ad5dbb14ffdd322e602c24cd41acc30a33d3971d8bcccbbe06f13986f6d3b2e3dbd07442f9ca7b88327f00495a974cd0bdb9401dd26342619ca72a6589a5f432433c748571d19cc87abb47f8895;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3c575e88d52054706acd999cf805a33ac3e83382e0538ef886b78c96416b37060727f03430b744e0d5bdf4d5c7c73f30a0898eda44c83ce4454563fd2dee0884289c29ff83bdbab558389fe6eab5c48c1b08ef5bdfddb81d62902bee380da6ecad3fc80d6feb6ccfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8009cc4578c6134bcde8bc100007217bc8b334b16a764098dcff34bfb588c6d45bb4d178fe9bbd5372b3e36280d8e78f3ed43c0cd70b5a98ec5ef39bf94b23292673fd6161869339f2ede69e28f02e00ca7ded039501ea63d787648237d85690245f8d067a98f7b9d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbc061e5620c5626b7c766647be0d14fbc0cdb89e6bb55e4d796b3e5f3b9cc8e69b78fe91bcede17fa5469987d53af3216cfda4a9eef6dd2457b94668ed79020c4ad8acc38daeee3ddfd97e52f74a72b576b0def262b0186abacb1b27f95dfef25e82b08ec1901e76a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a123f664ba1b2fee6741af883e97acdfeddec1cc1533029dab183e2a0c216d5b09b9a4e74560f48ebdd8e0e436c715d1048b616d59cde9959a50523b795bc9d31ac670137a826ff745776532e302b618bebc5b2e88b09da1dc4e20b651068339bd0b3b0f6b7becce12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc666f53e7c6cce50463c0996a0787eb87d9db773ca30bf078f0ac42314ea374ef22eb08e19fdba8bdd86e1df43642fc97c02e57bf241c85fbbb7c7729981ca637bfff3faf027e93902c4bac62d71e8535dd6f4075adf26a0d5d214ee10caa5869324cad42c28d82ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd335dbd53814e9eede5ce4680304c6d9a3a540c0381aa75c31ee133aaa2ea2e81296e194c7f5fd8e88194b7357072dd096083602e273b57afdc97f1965fbee4e32263cf756970efd8f61d1589f54f3c66847f88e6e8a8e529d09bf3f74c690bfabec1fadfbeec59e45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a9cccf4074fbfd892b2cf7dbf858050f61f63a665047ae57bd6694dd1c1b9e5f137c8d91785be758e0b6c22a5b4d83fd2dabc2e9209870cbcf9e9cc5849a0c71c898d80ce9679ec42e35379bf52d074cd4174d41e2459990a8cb0c7a2fc1d488f09f0c9bd84d53d5a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6078ab68c24477dc5f86b888bcc7c5a0526efd7307d1efb45cc6c16b5ba36fc7853d2289d67d1ddcdd9d6e96ec06a622b82bcb30feb5af34446af4687b43b036db4e092da4a623112e8828087c3ae1b2cdb12dda406f2bd07aca0a1dd34c6e533dc4137f2ccb67f4dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c2395a03ee789c9e3da7bb3358b15f02f454691f8e175ae3250ba33edf1e1661dc7a6faba7606eaafafd57cf7c7a7e00efbe5434f94c09531bc3fd0e87873f5eb64503216b45017c88614d483754d07bc4140c827496d93e6a0fd8c0170ef6559364570d1fa6248e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17cd0a6101b33e8e7fded744046361848c48a42cbbe1ec0260f62e1f6998f11bd4bf0fb5789a2aae5ad70face4a01a6e3111c65d7a7f0a9d468b7fca0af0dc217c8b7f53671ff4af88c2e63cadf6eed0fafc47264de3ae83c742641cd859ba2d8551e0c0436fd13f2a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d01959ed810e2406737083862a7ef1ec90a89f3e891e6ae24ef3c71b34ca76fb13b40e8c4224ba01d3bf9deb9b5f7b07f40848d5da4294c20734f9c8db98ea5bb7d52ff06f4488bba339ca0f19c95b7d734bea259458ef8a07e83da8fef99afd548afa8f5f9c4b3c3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bcd456534ffc9dc11f604576cb211ea0666a8272cad05ef8e5c892cd7796e4f0e12b3d796905209ab8401e7e76ff6bacaea79cc7a4065fd1973f4899f9a273446b1fe0175208672e5e1444a17f58480e6e8345417e741b6445fa91991cda448ed4c4a02753ca143a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a6812a1633565139cf1b3cf6b03927a24b269b276b48edee92c9ebd5703bd52a4ebf6910385f02a7b6907d755fddc3b058cbd1e761a6b88f5c523d75abe53a50a19144d68130b260b2ce40e7f5634af8d4fb3944db24663f22100126ac0c6cb4bbce9404a86438587;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eaec51c819bdb49a8e2e8eccefb223e73bc93223a9259a0c45175ded2ecb6034be70f8ed3f71b4ba24d5ee10f44324b627b56ad744adbddeee6dff3d175c8cfebfe65a5f0b41e501baa1fba49a00fdf0cc4d0fc17b81287912677c4c48c5c8b235c9bd1e0ef5c64ab0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f70a5f6c6f03b3faa98c9a66e5d133fca71729413dfdbfcddaec3d4884f01723e1b346f149b1248fb1daed5b7ab77f657e1a0a98aba40bd6735adef29f58baebb86e103fa40d3bff062cb162c89f158c43f3656f3bb82c2f4fa4024b82ef924f4cbf2589f4e58977a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46901c2da1523f29bf10c7648ee632bcee49f9e216b2b44d04f021dc3b0a032f559b7e52aae21c5f89d262ccf1967ef2a6ee04187d8e2497ac8b977df3aea5b1eba71c0adbfb8dd0bcdb392d1a159145fb749e8a90529e739e64083dc14a5845699f2ee6c121118471;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ed367af13db1bfcc24de2d4b3a1bf29efdc8e24daa8cf0354607f8e17fa312f2eea34f9969a456e36822f893339bc403e07e91df854cd4beb5347ba8fe2fd5afcdcada3b4ebf7bb9e9ab35afaf92b02561c13bd846ba885bd9f3edd8a6e6e9a417233ffb0381c00d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b066bf44402733f49a55278f13985b662f81bccaa63826beaf6594d07a5800cf500cc9c8ceb731decab5e143cb5efcab7e311e5bc3877a8060767040d33deaad08fad21cf2dd0dded480fae9140cfbb49bed9f75e6099ddbea6d3520be2321e14f7ac55022c9b99bd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3524ef5abbf44ef28699f7532bbdf3a83ff86aff9d21a693ef3e5266b0f1f41b2f54ff6555c3af6df03cf764d97ef5220da6a85b62f099d73c1acea36f6b12e78f11dc15272469613439e1277161c5b810c4caf714924337929655cf4889f5fca65840fb3e4259fcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd72588b689675c14bb4ac40dbb1a476d35b54c3de756c83d4d10170b08486deffe401acf5bc9d5a2a63ebdc3f447e144c23ea5bc261989d0f03304bd5bdd4ec2fd9acd382cff4e73a612e27c30e86bf88ff86f2782cdb6122906425a064904e9d399cd89239cc7a34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127758801e08830b8460bbae4c774c74f002fc4005257e94fe5e77cb48aa0f454980f543a88fa63516979b63517ba33d866c01cf445640d0beac5d2f83643b9996c9ed7e8f3c46a05c3f75c4fd6e4104d784e374a9425a7dde1020070bd311bb57bf38d2e8b637e29ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf501f997c7d72398b49bf04e4cddf7936fa0928121c2a698db13827d9fea59074461b7bde4abcbb8693fb8900989ab818ea4bd9a481acd94bb48e387d4c32dfdeb3bbfb6da6013fce4ef78e32ee6bcb28c35e42d0c1b7543d7fcfac6ab1138605f8dc24b9c3a9aaaed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7bb971e20544a30b76ca08781aee2fea1f92f9620918e1debda8f272fe24cf6fa86a4377f5df87443d1ea2828f88c343800f9fb113f9867290fe793c1ad89b4dc16eed5642755e3363c07711c2616dd7a68c50044535d69163a2cab71542672e80a32c19611bf5d01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14618f93785c2ca341b86c58fffd45146ba7bbfda864df38f8e7227eafd86ea33b1dd7062722f993a2e2c4e91409bad025f4f080d253763f4ba3bfa4bb2ae1b097424939ff7c0d1ec8784f3ae0b62d1c61e5f89d5b1f78f0405658b07639b3ea946bf827954894b86d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h859c99a245b102f94642776bc78f043d3157c58cee85ecb8a423fec92a22fe0ccd3af2f4e2d723556a413254fd07313acbe76661c33e60a267ee033c785dd22f7a1804b8fab396c91f2056414038c7b88fe10dd5dfeb6f8de987cd9c43ad63f03212c885d13f24a10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he07e3978a5a18f801043b5188c639c7369b62f2ede97b0ccb08c96d3f531e260a33738dc7e96b9a151d39a7d46998cb1c52a3cadd03a12b365be16af66c15920158058b26d4c66fbfdc935570fc08573e1e35986aa1e7ca6c6ffaf2651b752d85a2d7d6b0ffd7f5787;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c46fcd268c29b7c29792473bbb64e0b0872b2b9eb2f633b5fc97310b8bf28a0a0d8ea1b6b14c721b7e4fcdf00a43b0b96484781d6c77863408a42dc096d25ef4180d06a45e485513517dda4bd043edd50bc68ef76b19830b53bc097ad161ba9eb65d3b7b1c50c29cec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h375ab1692bf348b8ffe3ac11b9dee7d12c374018d0bc24bc3e2940a144f17cfcc1b04cd85829a68af9877f94cdd83a670936a27046405097d995eebecf16171dfca9143a0bf23071c962122a781c2a2232a2ac3cb286e260613267d501f3b985ea5ed6d1a733e31aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc7104f2afa2d696b27775acea08f34bfc94c6af295cb6e3b40aa81b7ca244416bde1fca676ad9f133fe35906b17a3d7c3295599cdeeab66c0851bc9db57c9ad0be42ca3e3d39f26e49eeb4a0339b9d6678199fb1990745f3f1a1e606af928b5240f968b2620591d01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9d1720ce182a9a7d527a03095c76d1efb71396bcc53880bc73701ffe37a72d6ac1c9755946199bdad0317058bc1e22f028cce1aaf8973f088c5b88b47cc54d1ef6200a502789e82ab69c397dc19e20f8fdece24f41e3b9f9ff74eeadc1d95845eb9e5d388be319964;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d92078ce5db6e088ddde22a27a0475ff3439d83e4ba5ed8d4067d2efb9872057095eb13097b7e91bb731766dbeabf50955fd4c5accee02440e8d813efb8f3fe47f9b85e0641c8744fe8c9ad8dcb4f1ff32dfa732ee671f69ceee444184c16f0c0fcf9ddc6e04209d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9fcce6aa2e2a258d5f20f85e749aaca0f9bbbdc6b25389c53bd8bb6b82414a9255cc08afbb11d628e7501bd67bbdf52d4619e868ca6beb2f26efa4f42fd2b1ab0ad82d729b1139cae42176fba274e2bdf5fc11711490549ae5b17cba680cb50d5ded9c40ac03aa9f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3db6574b91ba6fb287e502becddb1e2ac262eafde6e89b44a6a4b20d62f85cf3923ef06013318ecbb17b000b3fe998c13ef694dbd74a2787721b399102c91fb3970d40a00d96922578fa76b2ea471b4f575926e8e537fc9ec031fa9a0e8a6113dea6868d12ac4e31d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90a7f6629aee46170ac011f66e8a57a7e51e4733efa9114c04e86951df2799080c3e0ff85d00e3e1020054dda1dd06b8274c98be84f8d6530f49e6eeb174270a075e2c291fbf632fcbc997d49b04ad6c67c8cef7d063edd5c59776ba43b853e18d2abdf33c8466f029;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b4e49cd5da2fc377b17f0e8fb7a465296d6648c2f4b8565e8956b7aeefb02eb7afe375c1daeedbee4d7cdd15af276672fd6c434f17d100f77736edc2638829eb3d12413a4ed5fd8ce34d081e8c6a4130f3d172a6589960b1c8d80b2586a138adff49a29476e33cb12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha95497b72f4a1b4287389909a52d051fb3d03d3dccb4b14a848c77f2f306fe8784f158169a028bde90deaa583102f12bdf343cf8a7dd4d3ce495fa979e294a490f9a8234626ff7c8d636c959ef0107a6dfac211ca1def26189a1116c3fda7655035f110921cceafac1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1286effb36fa129b860f58f669765737259fbe89201db2d1f905d94d75b2648ba85d6458e6e2e6e49afce723943a96c92e2f7e786524103db1ba2e382b015f542fb39996d73926bd4a396da7d9868e455c6a10df652527cc379b72fefc0e2b1697952bfad343edd4bfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1058a88aa385a60c6e5a78ed13f564b77f23a53bb87ccaff6e0ad80eae6badf432ce5a0ea4550fa45e6239c7aa76b38f70d3016c7322cf0537e84450eead1898e4e81f7e13685f78c9ef964013e8192057999fe08ffe517873f8646eb8451922ba4ccdeb3f6487055c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bedf412eed64e98e939fb212b10782ac6e378c71071c45a2aadbdb4010837973ce0b87d07857bacc6534b2adb5b93b99fe667e8ea44cad5f2b6ef66d4a997983fc5986cb7995ae67f671ae1b48e431c88da36a8e59b03399692b84081cccca464ba631b8e127e727d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5797b4ab432df86e125ccd2548cf8474497423bb49952dd04610989db52f313ee9b3daa7ce141cf8cb60de7ace41b29acbc11e407955766bb89b223584c0197b56fb3d743e56dc813414049ccbda717975b1c960d4fb4d0ccff4a18c7737ceebc16c7c1f7e1bed9764;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78c011ac5799610e98f1bf6185cdf81a043b6a74a4b40b7d2d1be58758852e96903386be49f16f407022c5bb2eaa98ba8f0c68921b60fb6be0250323bb90235d523a0ed08f6e7dc73e0e4772ddfc7c0188014358e669150765069a2e82c103417f096ad8ed62190d75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fd18a2df447bd45a532843ca9b231119a6a447181d8a976cdcf8fd68734ba14bffefaa3f9377cc78817fdedf667c86cf3988813f771a459f90e23059d2bd73fdcf71ef2185c8be4b58b13f161a366057f6ce55ff83b58ce2867a0d88cbd7ca9e7fceeb80ee50bd19c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e7b954ff38c7fd90e09b0737c0252d66943a1aa20e74a1a902c66ab139276fdeb8d347c05b5bacad43667c0b98f62f46f22eae7a8412b535127e4d7f65c5426308185eb031350563280e5581d74ec91cbe2edd22eb44efc5289bac056a53dbf2b68f860e2228dc953;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93f0ed2c1a33600e28716f193e8bfa7480955b3f6b4e290e91a8d8041751d01e0ae7af197015683e9a157060d80c46fbcc8b723cff115441912f07880eae5eefc68600107745cea7a9f794c4644fe84cae7c1b7d71fbf0db589589caca887bd51c1e6bbf3d522b47d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfeb8a39ef38558bacb0264f7350ffa17a3050eabc4d620778f05803ec9082237e5b9e8051e17390c43e006230769ec57578ecfa78229bfed3890cf45f825fad614fcc22c49aeb142823ccbd8832b9a6cdfc18bb96b7602c08d3bca86daa587604c70f207536e2d1ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11075a0b89339253a170e160ca8c6e3d7c091687cecde47c40554ee6693e12e12bd0eb83ea73155188869694fb1bdc77f78f4a76e95877564abbb55c7881a8901aa49a7abad906476e6331f9a651f8f3ceacc8a5dd0e96e97deb7e3e11d504130ad7e30ed65bf1a3425;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cd70427b9cb5ba802b878fd62fc1a4dd2568f94ba3871196eaf0dc8dc6d570f703310af354591b2bfa0abba3e64f43787a81eb9ba06f29e76d95e42721e19bb6045f34ebdfbf8f54f8f45cdb66e71f0f6b2c8b731f888fabfd0f7a8c8f5caf64f2efdd652dab68647;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8ba78ece6935732ca31cd290856456165cbe1c29a672cc07dabffa5aad96218156cf5bcad77b6095f3ef75a2315d14f69a7de8010e650aad7a577f5fff49adf596d24ae8493b032bd10c7e338a6110502f73330957d06a2d978b81d604e5719dc8425b0f38506867a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb21ee98c80e78d83080c5851b81ff25679b69be6dbffdf8419749d0557c81639631ad0fbc1936eb7447d2b73ba1e11355afb8784fed86f69ad0e4860eb285f4d1cf04dc7aad85a491d8154d861806f3896f3c7a8309c013b922b06a654e486fc0a39b2f29de13c8c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6415c6d1519faa91b805566f0e473e1e693d9ed557058b53b30c163cbe32f3daba2a8b64d17d78281a979427119882a761a5b1076cff40c52b65786b9478112728ee87d01edfd11aa4bfc7f5b07213ad5b53b55afb771c9edd64c31af0aa058e67036df1ebec168920;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf176a33e81e17865bd32bab0dd70c117b4a0fb5bfcd8684460359c283d3153f275624dec1670d827ba73a1428b43d9e1beb15323050ae8f7a136d4159086d154c1252a6d6a34dd42c935bc79dd535ce34892c28dd536fcfd60451733c63f94b65f55b8022334a01d12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3dc187b99a501b8a6c3039ff173bee668a28d22e9f99d7a59097abe96e76803db9fcca8dcfb7cb0ea5f28fc022ee7e68cb36d58029204277b666e962dc63cc7f3c243afb1fc90390229b8ae57ce221e9f1bcf095f943b47e58ec2d52cc8b3a92e49de3dec35efd734;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e94410aa2bd39d5efb7e120a700530e860ced4f3b0fe569434bbb28e496c4eec89d288eec71ba2294ced0842095218faab981357b14979e365b0b801b5cc6c4e5114474e3230079df8ec2bb9ea367e0ead28bccb8cabeae351e71566a870b6f4917166787c99aebb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd6749864ced010e6429ac2be2e472bdf356063120074a4d095f9326de9fac193e660fc9600aa9238b9095c56d556f1daabf86c2fc3bfcda3626e0b46089e9c95fa385ef9cb4d125cfef64b1bab4e8bcc8072f4d41916f22574683e8585de4b9da5523f2a1bf97535d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60a5e70458ca140f6bcca5262b00e1998e11d7d7749bae5d73ba5e27ed3614caf4a18db468fac25e6c5f763a9743e4b19ec2c35170cf9c8f3f0dc4d52da231b2ade74e6ef6744321c37b25bcf94eef8e320079d96e1f409e79e117333b647496a0b989da82d3c5ddda;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha550c163e2005da2de2b12359a3c3261648c10d6316c53a0b98fa707c0fcdd6bffb6f5339c9d46aab23b96c364ea4f674b4fb1aab9fe24a2d5faa854a56aca8bc87d79376483ac836ee4192ee3e7ae658f5b34081cb4e61e6fa9c1394468a3deefb49a5d7d03b9b54a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h495bcc0d1376d0505186c5c93b4b83da851aca9f5606bfb73c2b39598bff7ad0f3bd8512b80f7f9b83b52f3debbf3907e340c37536afd5d8c39d939f27446c6a9f5391bb5d01b73cc4422d42f44b40c1c7c9f0561d93d0e66e30c1f30bf77e21cff484e76a1542e9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166ae95f5f0ece2b8764b1a725eee913b544e9b7ed74292e813365a8e941b4e135b5c806fe15d49be71f022784deb75a2987e30b8ca3fbfe8d9db9c27097b7318367f97387e71f56bf3b2fb5623dfb13c73963c986f372159c859a64db253e17a9ace813fea1a1ea9ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e33991c0d986a4e7606bc52b561e6f946415dd2d9ad95eeb0df5e2f4a869221e5639928fa693b348b7aa0b5d2b3376a3b721427c09b40b6663a3f8e14933a74050ba33d609678e43d19979339f97805cad0d53a250297c8695483c749337529211fe92a2f8fb6da8a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bc7a3ada5b1eebd1712e7507c10a6c716f90ba37cbe55533b4d3c4d6c2fdec202db25096eefe9a7239cb9d94616549ac1d4fd3c613ac005c51746a59c19005f127550ffe1d7e4caf8b5a1eeeff5ae9073808441e6e9bccc46e06a16b11c0825c096067ac62a9ce0b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0edf8c2ebd96c057f739a34666e0f36284a147e99f30ac21c745ffe274b80ba3a8f46d9973d834771febe4d93f540d791f30cd899775557f46f4454fee89a492a12621a03cc4e7241e81529fb342f84c1c16d51c67a6bbe34ea3cf85c9ae8c5d0f21afb32ec14217b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h741ed1d1fe632a3114631cccc8742515ec2d02d67dd9aaac9b3ceb06d30a7f77a04f1131db161c95ccaf3d6d329855053f99d29078053fe91917797064ed8ae267167a82b0fcf09057d13c54d2e42c4a4bca54335b4110886eb3226012b391f0affebc76c72ea1feb0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c9ab3e7431b6e5ea7c1a8e64203a88a7afe352da83d465bb0fe5e0ba0575f08dfbf4cd2b0d26c53fe6c340e023a6446f84bda0c572c3969c31d94b1959de6da1a714ce6c05a12580d2e4bed11bb3109908b648a18b4c86da1225ad15a54def8d71aecc7ac435f8a4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f550971559fce521ab92ccd45662e6a544882abac6e85ce6ed935e30215c57953816c1b3e24046871747c45f2ad4f15e638442ad0af3bda1517a6b0556ec5d5414f4024e06d3db97729d67565fc61428d0d89dc04580d6613225d281c4c9979491c0468900bfc3d9aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7f4880aba08e75d14f08f3c2642a564157e856267753996e4f8a11aaa64c06d4f56d6b5337fb029b472b304faf83f8cec3612d1d12cd0ccd29101bfabcf60e1637880d3cea0be9ed2cbfb7c4f5f3f9b1a1594d68463f53ac57f4637eba1ad1b3a1db40d11e028e003;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197e9c081889d9ac61ea543e1860229b801524cc6a33d46ab5f6adc81469321864e48288949f0579ac5c9aa9b72be03907173122d7ab1cef0b3a7cbeea9857a6a3a103b351dbb8c8abf3b8974d2fab95da8dc8c85f773af5693a75331873bc76061dc5c6dcdfd694eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146ae78e7790e44914bf331d0ed4f47106a7b1a25060eb9d1803f8173e18436110ebf5298d49ca7ab4542f5595e04896ab828e1367ea5fcf221ffd2315367deffbd6802ba055a6b9bf880b2c74222cc8d9503d15e5301c8df8d244a506355a6f4f1d9cdbd5e82befac9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178e7e250c20df6b059ae8687ef340a0371b6c806f01a8a6d8315e6bc47388ce45ff3f44ad7d362c854eca3a3168984068a6838b5fe76d40eef0a16b02a26209ea2faaf6f86af4c2c8eb7e783bc4aae684f0fdbef1653b2b5a3395646d19be51c7fa1f4209a20426e11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a9f3a8a15699b0c34db434ed50e011eecd35a5281515c4c718996fe4c06300fd59c635ceab0fd69030b184d116022a9fed45841841bebef4ef2c2cdd3bb3714fb19731a73eaafcf0fea87e4358d0e5e5a9e56c77ddd1ee60f0ace9e5d7e4fbd647af18b8e029b012c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187c33282d4859024f530332638f1b45a413eddff30846691f3c44b773ee25464260a3d79c54c17c3f841594b320dcb40260686beff7e7cb37554d784b0c99f478f2fa4d98daa229af0347cca03fe763c43400850834e5fac29ccd71ac322ccf3b236111f2d3fe993ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1c54d42c884bc5f072036739149f22dda0427b2e8bd200dd241545b8d55836f068da112374dd289db6353633d8c9fb8476cf1284555c93aa62d681354874b3a1dd9136c38221a6214bd69babfe5eea4cc8b09411ae502122c0b23379d45eb956371a64f2040925cd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h765b32f3227dd3d9b5a617f0275a1700f8f17a7f3c57b82e077ca1e11c5ea6d0f410a1b8e79ec5e37a88cb815e1974f0c272c5820953bda7fde565885557349def2dba7f87ed6cbcc7ca3df85e42cfb90840a8878e641b6499ae141468da44ccce8e39520206a347d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c67fffa50217f1ced1def4d8ffb73b4a0c74d475e93ee91339e8953cea3c994b439c198f1a7d8f9701f073ac85ed09c5dcc995a499552d678bfd845a2707428258e5ca7ab0660993a4f4ee3d469ff47345bce941d945e29ba4aad76f5e9362756c54575e859792841;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16334a8ca0864d16c46ef59dd48c46e40773c3f022a4f3b96091e6cd66ef2eb7296344ed4d30d450a64e04326b48880871f0be48b035702f4633991f02fa708297f1a19a6066b887f72573afd92ea7c92c414c78e82c3dd34a6c5725cc36572c445a7a78a262890f896;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b2e2ace0b8fd8071469964e57abf7009e4f6fefd745bb13d6c118a9e9e1cadb49f6d2a52cee37ccc8a5c713fc385f64d53ea141c1511d3aa156041b6daa53b0263698cec43cbc4dc72abe92aa30b4447f0e3d9d2ef9a4a276cc2c573e36d080aa3e0ef5387435c00f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36460c79922c6bddd9f7938d28aaa11fd5e1eb6cec4040b3a67f2ef9d1f3dc5b8adb64215c8c5db8ef09c4f0a102e30bb7ac940727cd574f1bc2e0a99c9c3ef07647a997735f55beb9bb2ebfbdb43a3b81bd55446879879d78c5636f69983ed26f88a3b056ac34d896;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165e5d3de256914e16a39ccc4a19e47f5abb7c7ec84970cd6f8f305cd1d9d38ccc21aa4e87360d5ebe51168358b798222be092005aaa09556338b66f7c2e9ea4664d3548920e674b765f0cb2e649bfa3b239fa0498b841f7fc39c611d3ad14117f40e8139e474e1fa52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e153194278e566e035c2215209390e2503cfc84e1d32138ae1cdd75c652d7b9169f754933b87fe1ff29283235d3a389b585cc4bfce0f51ed21a55ff15aec39e27e6b1eefcbb22d4ea3bf31e249ab803254a3da00c91de2aae74e67702d0c2c97f9450897118de77f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbcea3a41e1f23cad211b358a8e6db405b1e3c2a60d6d4d565b301ea75e2c55e936317c58357eed454584e6aacb38f35b8c1d78d4d4ec2f2e28eabf6c1697f160d09457ec8d7fe7d5118d7ccf3887c099b38271d3a0a92e5e06bdc32283c2f22d00c6e3128d68fb8ca7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90d468cd362b727f4cf933558b22c35b8c9b47ad7c077e7fcaf38198d4e7132bcebe957321d89fa2333aa6b94ef195d034ef12e64d0c76fab34174d9c0f74e8fabc57fc556872d50cb83a9dd4df2d9b9f48ea0fe86b625c1c484fded79ae4a76feb987b29ac322464e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11638438538178cd2c5b7809e10822ae0dafecad80f593da65a7ea3d59eaddb77ebda972351d3b369a2c3d02a345c19a1de5b1c85bff21a660e856ffa70651ac3dce2416d3bd6ae9d81f3dcbb4f696fcff405080378efff67f2f0f5a5819fa6148d52357b51f510b21c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cbca765dba77dc4b99ca9290a831ad93c7727b3cd4d52cd296d1e1541d86feed85ebeb8df99d98d3022ae6bb713b4f63c79715280201504216ea981bf1f1481fa8290bb72b9a58cc5d5a7a5a51ec655da19e06edc03936bdbb1064b4fbf0e82b64b1de7d80596b943;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e080fff52bfe19284bffbd6c7184b96d108983f1ef58a2821d5d0f7707de4a1761f95338874ee97c171a9602dcadb2b770c0d28093631e29cba4f90e5fd3956a27ae8acb23faf3b8ae3c00fb87b488efbc023ee1e4ee641ad812e919f57d14a3822dababa86268edd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e6b54768f6c59df883c91327b349377e1f7051c36adae33fb4b6286199084a54af545bfe47c31bac6189db5c5853c9f631f1b410fe1815c2cbd8c3a29e8024468d47139bf66ed3a046ae797f30e7ea163f65c8eb8d2c5e6b2498993df79977123625d335b9dcaffc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10336e6d8935f1682ba5bdc7b50ad644f8cd72e5decdd202aff07186ca7753a76ef10f56521b22e427f5a38e47b4f7d15d3d49e72f9450a12fbc50fccfbfe5a0f2110e0dc5f2381fe5fb3b1d7003def264683b844efca9898f739b268b186724c2cb6c6ded42850403e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1d7f71772c2862479b734b4b5c21f7fb4f8457c76184e0a146c0269bd196313414ec772d2c7d97f799d1cedc24da47bc31c3340189359d657e3fa868e7e390ab5742d1b1cf199f62a5597a3a128114174f70b280390d2cf4116d685dde1ca1626879992b2e61b4416;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104c0ffe4921bd8c0aae995168008b1a857b8834dc34e1213478a9a239a3eb5338a7d7fe98595d09ddd2aad9ccca402343fd7797a3d69f4d31b3bf4fbe11d4a6f9ca91e8f345291e2ea02295d0fd94a71ad2f2c430ac20ca7f464a2ebd461bf13a13aaf7f9f06c9d1ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h372ff3f8e3ba0db074a489222154e32a963457d04b50f6d73d069a3c50294acedbaa6776a13736a35640c20f4494064163676456b53afce626f2567e78e9b4d62f8ec80d6acc6349869caabc035552ad5e4afc1eecaea3316adea16b7909e130648f4d85e33e75d3be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2aa9e534b947eb580bee79b1472fa9e385b51e1e9dd3bcd225186369d38105445b28a9183d5594ea5806a608ccfd5ef4e2f2218b32012d153c1a22514fcc841c46ee1c385768e6c99923490cb4861deb56f4349284126d75cec702ffa701f1dfc237982a50d80cbf4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bc49a0cd94c80dd406266ae4118e345262555e16e0d3a498fdd16ac05701f2e151187d42ad11f59f75b1958740e26c8e22e53da116c4114f4247924f2109a84c8fac4522492b666d466b8c8c9a95c2bb5a55805b1fe577cfddaff91d8e5fb6932ef8b813fa2548cf1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd287de88036c52f7b794aa76f41691b8aca6230779726112dc12c1c246f5042b81f22320e83bc32161f7f3a015c4512b75ac623ea6e737038c5fd01aac1d7dc02dfa0f9d3d31fd6fa0a807e68ca4a267bc360d9017b4dee21b2cf1a95eef59680793a9e8df9fd84156;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43b793c1eeef7b4c1e251f663cae8f55c7d9217bd494b237fdfb8db74250f92f12bc1efd965f3d29e1d4a57064e45cd6bd4095303c7dbb97b56db66547c448344caed9b77e3c44c1c00346628727c8f345c454cca35bb9f38bb9cc1a7912ad117634c0addb11a0ca3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fa1292be41fb7f6fbfb8c1e9b110b1ff4fe501c446573ec8b4316ad3527b044df255f85e20a81dd82b822f82bd77c6f942fde1abc9850e185c3611d3be04e9f7a23b3c7a569ffd38b1148e7f72880b425191863b081629ffc17d1ddaae9989bf1919b2312d79cfc80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3783bfc0ed89d3076a569b178daae973d500a746bc46a82ddf18b1fef011380acd85906a915d289b5222675bd167c2af11b364ab946bade157169072cc221227791864978b421422120286e1492cf0ed5b6e48a6748fb425df0abe1a9eeffdae170af13426123a0a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6ce3519d740cf39261b7c8db61416f6fd45794e4473ab1d065ef7817b4eb2e25c1c5b278b059e95473ad2c0e44728323481f4869a750fa9e70eb29ebdd73828c8d7b95c4bd400125f341b67d22e6aea1b035807b1e9af4ffc9976e771a42cf7c79c132bf0f56401d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e5687ed61bf2203ec35f59797984d8fe9f9f2d48cfcc900ff963a69591a3f7cbd0e231e63e89ccc90114b7379cdc59533150b17e3e9565f445dbc67d2dee739f4df6825f97071a42223aeb3aed0082d1344af8d87e76033ab57234c665e26e37e4ae23d91751005e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110b1906c5cc921278b6e9022ae0949883d13ae10530ae25da70293bd8a17804d4e09603842fac3ce0c28de833cc067c820db3a8d55a6c15e13e7c7673afee0e6179e5d66d89337162c21bc4a9ca734997b7aaf5ea61f7e3dd5e9ede60596ffba081e74948b1ecab62a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf56998b0597ae733486f6614d7853cf04dd40e851635c73a370d08bbac0c78cdfc0e5776c18c930232c862d73163754a165f6dc0bdaa7f47820b6b40c352733dc63ba139f186c6ad46dbdb5aea4ae856f16bbeccbd193503a6609a539f2a2fcba8f3b11695e9768c35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdeb364a7b4c68feb2fbca7950fdcf0f611cdb4338fc6173481b61d73cc5922664592a86467b714e9fa7bd6d5f1e7ddd9d093f52bd61389686c4934637f8fcf5972f71ed47feaa939c81be5b4a081fca96043544af83b9158cc18539c6b71efd0c33dd69c892994bea3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115686bde1bbc531a0b4c5d1197f1000f7ed78fa8750923826df5114b3e15f7144f174e5b8d45c635f08cc6c07691725af91c71bc67aaabd7bec8710466e46d0e0629b09fe7de15aaedbedb3f99bb09fcb56d91b52a17f4c340af94a7ba0304d8660f028051fc996a00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8faa89a2300ddd43ba660bb5ee72675d5211656ac387589bab7545c041bce00f1cbde040498642278d3f3bc07c1d3b424424fc2ab63c8aa6a4234f2fd57871957b4744d8985bf6f8e0771e87818e327696e8e290ee7f48954bd342f2b8406cac99f6227d76f5dba936;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be8a4c1f5f0cf373fe55a2fa38c3ac9caa875ccc66e770965f9794df75d42bd17e913625b0571f491fe3f2e47cc6cec18476a4c126faab9ea8db1ef4dd7fdf0fed554ad2b928ab0afff6d07dfe0f14778c52ae73261da33a8fb7dbed8b829c805d64337cdbe9883b89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3ac940143b5cf3fbcd9d1926654ffd25046c7523ff48769e1734aff6375375dd3e0d0e6f7941b92a52467ff4b70cef1e0c8fcb4021d29eb0a168ea2e96e65da92614775dd0da2cb78afb1a278d7b1aa5690a1493bd694900e421fbc55d7c52199b3d47b11c55e7b70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc25fc5f095a60cc3ec3b188885bf065ff36c6165fc0f53969423a25f4916ab57c41642b2c5588e572a7f7af87bdbfccc23087c042045489a942a73f8e15943dc834cc5a68d952e6fe792404a357ef93fb774b367b5499ed14d48f06c4289722c8145192cb6ae77bbf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83e78702abcde79c8df0145fc909e3dd4a088c4be0c33d23b2b1384193ac9a28b2a7d85b106755b444c9626ebaef57fe4c530256e681c5c7c00c6929dc6a96fc9020b9209de0a8a873bcf891eed9b68e39d258bbe741a3753ccb3637c891663205b896c4ff5068234a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb762da214914d7bfd8476b4e67a78ce779dec9800a3dbf16ad395944b4817ab0e407969ef052a3b1bf8dd59b40d529b03e01dbcef0ae97054283813a8fb05c94cb44dd015ef2ce7c20bcbef79da01de9dbd3cf9f0127df5dea358de8234257c865ecee84873b4a5146;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42e927b9d724e4631e1ee848081fdc325bbe41ac520550a35f7c81b59ad07c5fc496278709c30dd35e7ff31dd2491111c6d557a645a769032d9a333b59bd0a833d3c5f210da4e6163a91b6ea4e5855c21e91d0a0bf554dd8954a0534414be91374aaabc73db6621867;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137b9483f52a9d85d746acf16e10f187a58ffea01ddb5e202178297a8227c357a07b9b5ec47c6a11836036c84432b05d8ecca164985ed42dcc3678a9bf4056205748965f938e773f3d100408cc17919922bf1afb50176f09dcc45cb61558f136aec9ed4c5cd5c98b3ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4212f462178d837cbc3a7aea53aaa60f8bde4eca88c120e79dba3fddb2b036360bd85c80f67f07557d49ceea1efe988eeba070a7bd7df29600a3467bcdf52f0d972f21bbdda21afc668e52c98b182e899d864f38562f4cb99975329f181da098bb78d89d75cf11fac1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h631d34231a78399a33b6f40b35363208820858b337d399d274381ba254db931dd8ab8c659f2e748bdd128d7944ee250cd1263af08425c7293d222b40d223776d0427c767e683ca1b32364d2e0d7f176e4e5ff0ea0e41d12e722a52f2ae21259bdd6e1e3ddbbb0edb08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16227a071ab8826a51b4e44b3c3e4ee9d5def6dafabf8cf0bd4646a0e59ca707abcb197dadbbf62f7586275b508d4d76b574f2918e5cd2fed6998a5453cd90f8e977a6421153686a987154e6022719132c57176ed12ce1e5b5f00aeaed0e2f778b6f5eb34a1e03b99de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe9bdb823da2337ad3be32daeb0e58aaadd63bcdff05dd52e0ee4c409952d581650bf24baa1ca6c85379fc00f2e5de324f4c560920bb86538799e1880da1d08a8d5c3832f474c1aee4065f3133a35ccffaec739ad44fc154a1fe32302c8b9d32d8116c947ca93a618b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157437e4d2f12d4922c756b9c3381e957c6beaabc7516290d5e451edf252d3b0d69195aa3b75aac0061d2578f40d7da34e494c55d582413e4cb374ca71aa16b54459032d0e0785e073dfa8f0ca10adca00b244596e4743920d5e26a0831f82f6ccf5201c6225b03e758;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ab66be6572c2ea33d5984692b6bb9584c1b3308ffa20ba68d3303a81508e2f5c1b25dc18e4ade903d714e5c1847cfd5d9992f17ea639a9a2e119ee867d91ec8f07ec185c6aada32e85e79dfa7e47edbbbb6cd2a19fd3812bbe79ed458bb349f1009cd92a4de56e916;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153d58fd63a091f38167d55384847a9e0187480335a4785c8c69118e7701a5b8466c794904fe5ee8a4d3307d152f4c5165b717b97b9e535f7ea3d58be526cede7327d985d49afddab4770ae823c3342f5984a96727706a3a2dd24810f97f431261e1c3f67c42b38ab33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f85427b6a7cf05d4b90e217910a4e9f56bb0029aa6781e2bb42ce2ce457e2694fb2d193ce5ca2248a98a0531cb74d48d7311db379d5bfce47d9b77b6338b263f9e9192fc3207f640653fe7f99090520956c33776b3827c3294264ab4209a832fa6fd6fa67b98e937e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25ede21a3f5c18b35eb9db06f7f3b361c1be5c01da66d0dc750cf2b6efa34ee5e175e5f458977b2b8d5da03cc313ee8d383847ff5f8b3bd4a85036e33b3c03d91691b2a20869f3d090d5721425da5aea0001c59f5abbb866b7d5f82d69367b1409f4ee0f8ff20fcf0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb706206df74564968cd64cd6a86352dd12efee479f1a6087cdfe203fa2d107555c4ab7eca282d021e006979448ba6dee0beefdb1eefc44d29d826b6fe646e2544d4b285a2ad12d81cdb01e653be13bd50cbd32c8c6b3beee32b2e9662f795eaa8ba8b76c772f35bca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156452c781b70cbedbba30b5f56018f78c54fba33e37dc332fa88854abb8ceece8909e52b0d924a6d5185e0818b1690ab4f2659a3423dec164d45086b3a404ee425bcac828a506a6412630f36b96108e9dcd98686ef3236556f070312db2045fb403b80600316be443b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70c1695e3036f9d2fc8a7c74c75b571db04956c0f98d1b95711bdc877963c227750345657b8791873f1f1cf45bff5ad770fddd5be9d6ea9ad3c2cf036df49d2ab522c1d3decc52d4d2729c1df5e44e476a0b5a3f4a29b75e7f8487a9193bfec596368977dec1d98366;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hafc2816f593b8a12b8f1800a7e5f3ad9bae677928e91cc1cffc3d58b325c48d81fe38fea73c0a4e69e719ba12c467fbbf2d12312ec1b95ac24d1f07cc4cd95165e4ddcf81f857f79fe0743929d07aa4bc737a36552d88dbdee99017bc4d65be8cae25056b66005300d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbff8becfce2e350cf4038328de3a9a70a0657b2b82bfc5bb3e724f98230b9d30956cc03e788cd6001d2eb027854aa5ff14385142db6e5d0791aacbf8f88691e9a1996d9e9d1363dcde85fe9b44c15e721e3a1ee516e9f9b2945b2db7801ddc83c03cc8721fe3c1214f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h947d4b3439802bace151adde8f9833f83a9d0ffa79ef8275a40d4cc8ceb1b81a608c97d72252291490be86820be83e788dca92e2232f56a79af4439d3ae96de5ade2e1dfc4baa6e0d086c473494fc68ce3533d337c616aa14c6960ff6d2850b61eeea8d616b40be1b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc47bd7bbbabbbae90bafc45d080d2b98eae7f09c673feab2c8bbd522186d579d2c3fc41c559c643b5031c3128eef000dc245fda2599f96abe47fbd0d8c4434d2243d79085762e38cd52bd89119015671e95da72960c4c587df654e7fa00641c89850ef2aa0f1e6c888;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e339718622d7afd12b1ab9e8512f698020b4231cc71d64321defd003244b05e939767c4a2c40ebe518501a832d7c182c688af72332547c06036b99c817913e06ff402383b201d98b5e0372d2f5163392f69161ffa2fde49a18aaf050efdda4b89fdbfc2f3a19c6a7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba63f54b9607465a5cad2f70dbda63396f4db3b29a0a702000f49be72c2798cf0369c90b573bf4e5d66716be74ee9d0d73447c3a0455ca0bd7e3d617992240e29a446a2448b95420da0aca83e9d8c200a26b012fbc6b8a9896614f626141bf54a79872312c13bb3700;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167d346c813a22cc98cde15fc547ca6674efa1a7c066c3d72dcd2317b02f8d8c6b85d18f8edcfef27618000032d485c2641a3c15d78ccc32c43038c1676c82396129426f6cfd3bab4bd1744fb0b68295e03a93dcb3a20a6adaf419e7c16552fd6580611cf13fd8c04dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc888711cae10377fa578787e5f11f2405f0343c84800c16a34b13014b8c099238632e4226673e3abbe0a03d28e15d7f2fda4d7022bcce644ce531b0d33f6131c345e12c1fa957a8fec06a2529603baa5b10550e289b9d9e17025a3f922decc0763e70577fc142fb2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72dad2049bc42cbe64a64606e0ce14ec2125c4b62bc5da7f3cc1b17689c9e3b2d3cf7bab3f4e439c2ad6e28f6de87379d6cff3b1235babb186b19c8b30b76208c6ecb24357ad07438fbea4ef5ad324b81a0c7ecc818d04b51ead3f28982ba908da119df5b44079bed1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8c1862de12cf9933477b41e63c989422c4e7d97e3438022a4e3bdc58bab20c69644cd8b3b880444c4f1f7a8cf37ec569a6c7588841f4d5e77b696aa6a69279ea7e88b7e73d4113c2b9fb094ac48b1bd1587d102553bd3a559024836ebf968058a24c9f2e3db0bfa3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c25e17a543d54b06bd13e8c8a3085dfe8187854a331ba0ce669c4d78b0c3456f41ce4a9eb4334cb3e2dad7b56826506a8960f186941d66376836939a95cdbbf412ce218c6a7e4d6d3d5248dc3e4ec01a5875392fe531046172365d42ef8ca3cebf83bb1a1d530ebf0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171b016f92ee90a715e8a20cdb1853f6521499537f2e5bbb0e59ae79d50e094d944f4bcb02da131a0bbc3f518878a38d71f984c612468f0b5d8a05baf23ace071e3a369b6e25da43d79138afa991de5c4382207dfb70bc67568a1c3abf9ce38f9b00d5e4a201818a5e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1407d07a8d6744dce6a45ef5b9da2ae49d39c5e512c01cae8e9e6a4bbddcc08ee51f38511b10b61347f8803e8e52580b31f6210e472aa2239e971ce0ad6dcb663bb44b86a6e03858b2948c1e24c25e51114bdcf5976eec9230b41c6aada6c772f51071ce6fbaa97a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149a6fd0d44717b40545ed74e0b3b346e08fb9b7e003088d79a5e9244954ee2815e668faa44a658b3b8e67a665840464c6bfb6609fd250c9019cf6b663ac3c94c38afd0c773a64819ad2c13369161121ea9b82d77fd5579bcb05bd1445cabc1021047223303a5612c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7b253c2ba4dc4928a3f0d042d549cb5a1ef4caecc7e83fe63c9b2b2445eb2a3895d8099fa598efc77603125f6f696c21002bde2774a17e85edb71c20d3223ecba66e2ca1f41938b2f7d59f9626cb0b0dfee3167ae2033bfacc8b774f7c5d202ae0de93028eb1b39b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5e893ce7670dca35625f58784d3f61e3aec9b9cb7f62dc16842f551fbd9b00b73b18e04432c022b3e6e945ed5ff7b52ca34abb55621e5425eefd130ab7716f7dc2601bea687e424f8d5320c224e9f31de90f2ee19cf0f60dc6f616f506f1136c1bca2f752a3211d79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdefbc7aeb85bcc565e99bcb90b746eea558c24c307b44d0aa6da454124431892cc64ed24a23e885bd7690abe284c3ed5c02f6c045d30285d40f840068bd0e3db1532a5d551fbb84a6672ce8eec0476628be52aeab8c098f7459691c1e858bdfdec306b474fdbe6a3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a20e4fdb89c1362196626158c8c81031790a6c9a795b71171cb0a8e42fd4012e4c31b0c8ccdb917c7823ae0331ec7b5f0d4c9b2c04ec7fcddb71776acda197b6c61babe16485a21b4f68521d23e7fe05efbb749cbe9b967b87ecc012b07db07037c708bdb3ad36f18e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2edbdeeea485bf5d68dbc9982d5a775b62e7db4fb4d2f601e77eb8681a4f82c4c629646131be0b43bde2b7fca1d54b7de82b4f2c6d993fba2354fdf7e6ea982a04651b5c9bf69954cb672247ca0eb3362995abdae47ad0327ec4e6e5be14f138f13e45f4e3fab4277a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7fbe2ff79e84ab92a18639ced1852295cc97149250fe7915fd80cdcf51df991d90dbdd5d03b84483d148d803062cc897665f1c0399218c048cbef52b2c20e52eb9dab8a37f90d064914a0be9a271b86f43f76e318e1535bf4480e2268889431402e228f4181651d8b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56bcae0818b072cc6079d128c1d8888a844ff4d7e5f030e0d5f45d689dd35c64c89f3fd7e40702e5d05226d6c5acaa6e505a09093e7348e61dcf7b7d61a1ca3e9d2e124d895c245a36e9e9694c4d04eb01d193ccd3646883f2998d20f8d342b1b97b1f5d0f9120c59f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84c51590d6aa0399d42f47d65291060f326481773c78539cbf0728a49d009dd75b2db225be981fc36707417e3d7d67bcf7f4beaba70fba5bd7e04ac985ac6de325e7daeb899d05351fb32e2508a3440470f2baa01b41a18905ebc062cc34fb15d0b279dd761be36bf0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9eb11d4b2e1f02b8e8fd6cdeaf2e8079761212c431e62ba9894e2aee93197252066effe67fab02cb25d35d9f8b0eccb7bb3ea7943857399c708474a06deafdbe3328991373f9a14e08325fccd1abd8b97ee814a5461579bf4ed532cf59f179a827271a99d1d0b00ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1205031a3fcf77dbe0934ac9291186ca779dbda2e34aefd13c9d50d42d52f2cec425bcf6f4753037f8213a751526da4b2ab1f63ca82affbe5ac8a4cde5bf54007a516892519cbf02abbb97c508911c890f6db0830683d31e7b15f477507c1299287b149082985a50f2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67cfc4ffb180230c22d85c96ded894047ae05a3c8a08d3432067e6d23b391c8c50a0af31da3ea87df1fb763f404694af953b223741726b1e0bcc0c0631a998158ab7682e7708b7204f898fb56b0e227896f6ffdcf00424072b9c04ab865abf35c5e14e40fff3fd1569;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18108d5bd2560c96d23a339efa637a0d62d3fd816660b0cc0053a06b77271f496451a1eca54dc1d487148af065254dd280d014afe66852dc33fee8294a09854b1526305c27749fee5cf7fd58c2545947b1c474da5845346c40599979c8e0e66cf149a52e88bf9abc2e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f059d4d238057dc7e01f6064fca98c0c14a90b538d402067bb63a5981135b2c88abb521d362cac11705a6c5218f913e75d49ad68fa4b4423b268b3b9386a264dae2a37c8788e62be7ac54c8778f1044506b93803deb96f75c049f3f83b533e8e4e90399e9b59a4a41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdee29b403459a68442417bdfef6391da8b5ed9fbe2a35d81e7f3d7e7f2a8e23e64ed12695de4985619e5c4b46b87ee205dc7d30c3cd25c9433e082c73b2765d06d0863b5552b3e9286889c8d89f35d9977676447852aab21b1ce65c3e7fce0b9bf7cf4abec10d01eb3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c58bddbd0a286f607efff27889dc3d817feb03230a160c405738fe6f45dcad73ad9d93340d1987e4413b1dabe9e234146d998389aa3a6bb835e572b361e5d16a0ddeb087f577d086023d4b7f43e0233c67906ddcad037049c168d6ba12da7a3315583ccff2f3237c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ec51817a8db2cfb428a2e062b56a76b40b7a077ec6b4e516d0006065bc4887c1e455a25974ae62436bede8335689303c609dac7d60edcf9c639a1c8aad09e78bae08eafdfd161193db84544bb69044eac0940dc12b0edbbdd9851609cc295c570b0fb6c931b5aafc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d639c5f5334c381610fcd89f3d55f5e36ab0e4c96d90c4f6f9d8af84e0de938588976a18366afff378f79ff96e59cdba1aa74b16393c0f8ad0353027e0c21dd5e622dacfa9a85f873c5b3515e3d21ecc5837f7e82cb834c58eb90cdfe1147cc50fc26dacde8de7e2f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6c25d5050b451b96ba7af28f7250a06b9ac12b7f272ffa21d0b71058ca773063c9b7cf2125995def0ddbb1e2d2ddb316ad9ff2fb0866a8793c85b6f9fed1504ae4aabc5fcbcf88e003a51bae5db647b3fe37ec7ad7ff3bc87cc00678a41d84eeb06768e6f3a177063;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42d59fda5dd05c7c2fa7561f437fa19a214c5b3c320d39c99e07bfa958860054a667b491145a7e8d732107011c94fbb83b213e62c0e3fe634435f81bf918c06114ab2e3d77510360a053af1499901efad32f0ad64bf9574f1fedb6399a6a4d72848f93c2be4061dca1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ade0317eb7127eb055ab39da17ea1ad6f1ec91ccdcbce0c92e7df61299695a478c2ff3a9cad4da0baca186dae91671f101cf84c83b1fdf6bab9972cb2f3416fd3e02f422117b81ee06e952dfdd91675a4c313f48e3ed5bdc372932e9b7bf85a564591797be5e37aaf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ddf795d213d430096f2a5b185648a48ae968a1394ff0ee221f940562c7ed0b38cb752e4eb47a9e65901cd05e69d1dca65b31df1066c93f42d5b27d61f3ee0c45a6e74c335fa7fcd6298a8e3588f1c1ee3c4573699e1c8a7a23985ac6a23a765cf43b5a5f0e4ca48da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf20b92d44ecde8f132b11280b2b0bc16171ff840823b0480369c41cdf229854f12015505c8fd6aeb9f8a9f8ec92d9c51b4bcf8df0d8209a99605274b78e542e387fd00d777cd947a4d298e8fe6b3333a88fbc677d0845e40d23dc47ec509171d998ed7e55a5f285ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170b5adefe7291be74fd6ca08fdfda8092f396f4286379b896938be8fd8f3c46a317c50c0af21ada0540b41ac9e9de2db2e8ce3c02943f483ce0f3f5429e1bbb39d74d5c93bca69c03678763977ab2c23ff61901580c94ce772f2dc3637fd6c98b8de2f634c2bb85d04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77c4b4739aed7fd34065c46267b9aa42f963440f02065a658d7f0c330e897c8f9b489107b453a6d4b538e1c791ee7c5f5d0536cc5dc4cd20714ba56353ff46b010797c4f5c4b564267c06e0d98fa5850d038859a07a14b863ed6139f36b86d22337c558ecdbdd5a4d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22b0e9228e5fb9fa902e745e471c85f69484933b2495148911e443beeb079d127100118ae84607a1627c20f3c41e0bdca83a966df0cb8a9ccbd7b77a883777813b05c19c2ecba2fa6da1913b2e6332082204eaf6cea15a01493a43721af5aa82fe9c1910a4222ceea0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b47cdc584f26c6b9fd15285f0b834cb110125a1b4cf47aea3894eefa005a552b7912bc963a2cf7ae2ecd55907b213c0a1e7eeb89c2c5fde3ef1ba6f625237a0da1d77fa66857b61779d1d2e472dcf2c70574592f836f3c9d1c5d51ca5821f4aff5019a3e4c2e0772d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a1fea69ca1a3f9f913654bae5b59dd7f898a2019e61ed253efd2677349b12a97cb25a22c9fe1a024cc8bb31f9ed367265d9c8046d2ddb2e705d94c3e47bd95b6beb90b5a40557726438b0e94f3a5a7d122989bf70148aed369c475b6aa24fabaf3f8da280f957af5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf376d6c41bc71b92693c8ac14d3f50d128ac45adc061e796d03e6f6d431a3adb6058cc053914ac50b87b0aa8858e233e1586a8b7030fd9f31185f2c00a11d832281aefa371380f30488c7da229f246517e9fd2de8228113c7421bb7e8d9256d4aee86f5210d1b8996e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e43d7dfd481b72b1dc56db510b4350d190b1be723d0b2ef47bb2368ef10d26c0dd484a2ba63d4763c0262049abbde9a62c9d56c501a4850093481debf203adfdd36b5ee177e6138b2f9f712d88b67223605e22ef7a4cfdd14d9f54717a4fdc29d46c3e6fc9753cacf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc5d16d2fa2f695663fee060fcd5d30b3d831f5068d43bab60e8d2bf8341daa0e79ac8fcb7b9ff099b77d60d952a5f470f34e90e63dc676a66d901f725da0454b3d2f2a6b1dd31805867f4b7ea7869d2c3aba52c5216eaed6cd47e16c9b3bbd564369ff6ec3cc15460;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b3bf1461fcaf77b79a5f3d963f8589f2304a8f9db683072990e413b21e6b9ad1a844eb4cd56f3aa38cab09e5f0130d1bec531cf9f8bf95c5d97b202a54b3f04ab97bf7b49f2b18697485de2f2587629c4c5663198b8c094da05179e4411b5db1dde10a679ad3f0875;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcbaacd6df16bdb10d04c59f56a54b7e22aad6f343b39a9f1bc3ddeed2a83f516d22d127468d3b1a6c2e71a645f6b50fbf3ce9fc33eb2c28c83c91f0e5afa8f46695729c01e305293c08857c67da0aec5f6e685517a7b5d21da0e4f21e94c4a0e7dce39a19e8c16ef31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144ff3f0bfd471537b880d7521c6e20f1a052a9e9aefcbec77e3365b39fc7bf0aec47ed16be8b086192cb45bcfed07cc2348f26f6fae6ca8168904417c22dc30c36b21f269daf069fe7903892d32d19b96987ce74d5f6a5e80ee74a0a0d0ccce07ed93cf4dd56aaaa23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3bac68b2dace350c4a88600634b3c71684cb916b736c332ff2b64ca0d7acd28f8248e0522888e537cb9b7d568c7bc8a163249c2e2ceef5f5be737a3ebe61b8d0c6e410b7fd05c0e6cac144bbf3b34ee2aecddd157ca9442d164ba4577003cdc5fd31fde814d6c0914c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167cb7ec569f4b3c15e1967e808910d26a1bd96506cb030a561154f915abc5578ddada2211624ab643afa37439306f807316552e7e4031bb7fdba4d4b0d816f7bddd9c5928564ebb93e3cf490a5585463119f75be4cf9d873d69c1ba7d4d77c2f60b82c5a3bda389812;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177e51e18975e0863468b689ac8f38dcee60206b24522744e1283855e00f9bfb34f96eb6eac0f11312c696debce770bc728132be934c92026e22cd879eef87cbe9ec86383489c7eab731823d4756eb92514f439c3bd17bfaf392bb6f53a703ace334011a4bb558fa92d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f306d20f496e188bbb58237ed4a5484445a2bda36d09f6f59cdc80fc76611b07ef5406eca3ae07a6c31efeb5ec2d3afff7d4be69a3c4db1b623499b84b00809194e61820c5d1a418ec157a20b190b91d1fdbb8d057b4955ce72be0544981d36f419c41db0ffaf0b1c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110ed6ad0476aed03c0b0e09ab39be8c994707ef8eb1ee0c424c3e3d34e0cc99ef6933b482cd4e35e2a9b7afe412d674479958a9c171b6fb781d457d1a720d2a3bba0d2eef12916fec63473d8ff1e4924f2925e04fc51d239f63bba2b3dd1edcf490f78c746ed427f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha62f9b249310073b7462251044a9cccd1caec79f3c41e7ff2780d162b4ea32284fe13e01555e408f9d70f354105273d05c2678cedaf56743beec4173c8d09f6dda5de3a73c90d88c91588010d05eab4248f90f2769c8d92acbbcfefdddf91e444e580d16e08a289861;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1039195f226da9be1d8113aad3fa41aaeded0266acc43243fe0037af87e6739376d4bbaaa3ed76c6c1892cc9d589ef7ff9e879c09db9d8b6b20d0c99a8e23eef40c3ef140eaceebcd71fe27a9f9c89757dffc3915343520a54b4b36047fff5dcdc7d01278aba90629c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13095fc232301a1c9eee1c7b997a42a8912f14ff27d9860f24e4ba2316071a21ea3fbd7d00c7745712b6aeb38638b2786bc7ecefc89a688ea94f371fbb63dd7487e92e58a8e5234858e202de97d9921cc2729ba00511b5e74b004bcda467d67c48222c23fbb94378cb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42f780e2291c2148ebd388cf0140421ddb05ffc33863a5a2f34bf8e1176f8fff90299e74942599a660d964403288016eedd5d694ad309c845984e53a5df74e9d5803769a173f3389f75a82d8a1df13058e63364942bd9d69af183b3d8b1c977be4724a16a843183968;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8009ad40d7cf9599e1724910402f134ef49644f2159fec8bef93e6c744d23e631bcac971f75f37cb6e87a2a0acc950eb547e3653e923734e0407f0191d6bdb165074b4c9bf3508325ae044f51d0000ce0be471ce45b33bbb42e6b86cced0e32d37e09e31f01b5dfca5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca2f758ed98b070fb47adbfdda291baff9aeb181ec2149b5a71163f59b78b40cbc08393c75e8ae46589968d2abd06e8d1186f4d7f7eb91ea4d1b2ad621a76bacf1c4266416dd63d05301c08abdf58824451312b0808e490235a8acbfa8d5231fbc3dc470a3dbc3b0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf03cc35d22d7b403988708be15f8098e29206eda9dde8640ccedb5057ddbda3b1916ff5aacbe46b1351b6b51acb905429eeb67816367d3dfe3269f1e4c519c1dba044c51770f9dd6d92b5fa4d9f2d8c09e333a0699f65c366db06c8083da2a280fe4faff3dc9ead21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5ec52915e5a49dd2205e8cb6e6237717ef4dbb9a14c3ac72e6eda44c549745a92bc003054bdf1d1eb9a9c0feb4d56b47434ce55b8716114ba05bf762b6622d26c42b14a17f97ce3c1bd821f0cd2abe330fc7a54aa4d925f11e5f0c6bd7abae0980ee1735143b3b977;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9dbb552ab6ea8e3ceebc94cbddc4dc3dae7e6095799b9e81bf7d891ca2290b04f5da4a6d78db647ca659f21d177c244d1956ba42341bdd6c59910b7ec4eba50a0b92cd08dd1aee41acb1d372056ef25449b47a80cd66f33fc0174489a6dec5430e7a465424632e5aad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b31b4b17107b14eb6d2f05b39beefbcd8abf69eff5e5035d7cc2affc0c989e8d0d864a075f1a23278512c77e6dbf41044cbef4fa68246e2e467e7a38469a3bd724ed97d92a6c6bc2cebdafd03060688e9c34b876b64f7f96864247c72f620f8d8331738a7df63f251;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140c831164741d60647fec10cae1f0188e1f1a923a0c3f9976504f0aed9026b4d4b7dd707e7fc4f49872577e7c8cd921eb885ee165f6191bf4d9e800c004e3cf818edab082b06b252f4faa64ae6c5da1288c0f232747f802572f0eeb3dd1d512643641be3023bd06c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b72a7f684074b08c51e132b03ed1b21f716484da2df492d183524b8daa4e0a9724b9177db5c64c6409450dca3c73ea166b75af1657bc968acfe986cdd2f06ab14da6b969d5656bd5d26432c244ca7cca52716cc93dad37e2291bb4c12f60b5c01efddad4084b808299;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8a5d3ad21367d53e5618c9a4fee9e5a3eb5cbb5d8960c349e16a0560dcd6744e7e6000c95f7a1cd1f3ecac0898d45e19ba8763602fd4e6c4bea43733271b3dcf1f9ae4b69f8b50a16cd50db833591bf33b1e0442144872afef261252a4e3deb5f94b4346aff4d2545;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e7fd9ae9775d9ad5389b4ce26758a5f7821efed4341be4597be2de793d72572f11cb7f3dea8ba0e1efac8a75689b2d5a2fec3551fe424f4fef68fd9a9d1123a128f1053d073105f3cf56de61bc63d430918cb4b52c98b821d8f5988e8feac46d110d596b92caee990;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc67544579c301c9efcc8d8ddf087a9e8491399662976356b31612f689e8fdabc33c1807bef5c97fcd2f567c11a0c4aecc060f7c90bd274e758958e899bd477bcf701f87acdb16adac4c26c5d8e954e6d8f8259d7ab118893b0a5d536d35efefe9c3e9e06b7c40ae9b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15683dd01c8dd9ea6ad3611efb8894c3999026aa078113eaddeef216e53b0d6cf4a9f31ab3867e58b03349aa184fd5a063be386899c856f1f6f822a9f687e1acee7e253899ef16f4878b4541781e0553a091e7c48f01cea2ba1ecb9806d146dd4599fb2d472bb134f7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e34c264a3010956dbbcc4a0ff7f088a870b7641d612c8bace89702964623043a04c2f027677ba39865370ba629304a317b11da473997b26da808bf09fcadafc3027c3d293ccfe5156ddda904142b52290b157096b54b8eb2202297a16edf12a2e1a90e793f7bedf4c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbda63fb80cedd070c0117304602999c6263b58cfe5ae9bd6cee3d878702ccc04794a9b11a7270a644602bdf672a75d32afe981f38496149b613e05a86f021937bdcdfabf77140b364103e97967b33ad154de03f910d453a287d07358e2d5378cb59ffc7e4be202305;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138e52a7994ae4a52f68d1a2dbc88cf695afec64a46922aa7743fc9a4b98c916e3ffd0bcb1aa7ed94c80f5470bd5b16ce30278d1c363b18ed6cba241f2821be744b341490b889d815ecd65dca0aaad1c9c14317c8671a765ed5fb374b615fe111f75548b770f9d9da84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfadc31066048db3e90d2086f0b5029d0894034ce34c083c2bae4e3afd63accfe334864c44e116f04acd2f43741adef957aafa0a7608a9eea8642fef17859ce891d6261b9239daf2dafd14ef767e328f56b5e82713fab0bab7de1f4e01a9e8f7cab1c1f5430704fe9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1507a9147c348f49e30c5581da0b68ff0511a2651d81b92824978ffe5fff7fbfde1748f8fd0476f6564937724c321e4da82a72b122a0728eea6e6a22cc30550f1516c197d9f31f046824b8a4c40517272202feada4fa38a13713eb3ebdfbffb3167046cee11673f4b04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb2df4e362f18f67357d323c6d677fdd4732e2dbd82b691746e3b5b3357d2d4d0efa372ab4b56555bdc1218666d80f57dbc61fa5865160b14e5ab0e02379e1cbf074c19070628461d365545467f81111071492f8f8ea48ea59d5b3a6e124701198c919f49f3ce37740;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16432e1c6dd2c7a33a5659d8ff2ef3b1564bfce5b568d6c7fa3db00b40114f516310b51322b819d0a5550e0a3320bec0d9294fca5fc67cfaa47b3a9b201ce8fd09d0cadb2a17cd1fe1f6800d08c2438bc078423b0713dae4b1f20eddbc4a79048ce90d5422fc1b8be2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c66eece1915bb5eb3ad0804fe32cbdced025570379975dbff71a09950ffaeebbdb7dd70d85bb1b82c3c23930469aeae821396838036b2b66ca5140354191831a58379076ae1208b8a4ebc62ffdada384dbc841c7df95345c328b51e4908fdd8c3d20cfb3587a7d41c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133d48085504533119e3ac181c7bc7bc12395aac7fecfb27189d2fcb18fe8e7f3b37197736f9c850e1e770155db29a3b9f54c4caae77833856b5ded2a63960c2bcbffd04b8e8b0b88c87e19826d93037f2ed66c99d279290f0c340a4a72b6a378ed76a5c1d47e86f0a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9777e9523724fe0750a48320528a5467a3657f03ae19fd93f4be3fd0c08ee76ce11c34db16c38bdc63fc78864cef1d423ef3d3aecf30d4908b93b9512a600ece1f1cb72e496c0d2d93618e1a86fa8db7b913f9c76ac174d98d1591f030f959950c21b76f8b9262d9aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10df1e4a8bba759802d7b5bc3abbc571c067d8d48a2330746f2a4ca120ba635a4ca13881fdc3a071c994178f9ae42a33220eadb45a1d7db99904964fcbf3c0cf2ae023b7f643ac7a42f4bccff1da2094e2370ca144a828d109a68fca7925a715ddfb78919b220d582b5;
        #1
        $finish();
    end
endmodule
