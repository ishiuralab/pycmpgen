module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [25:0] src27;
    reg [24:0] src28;
    reg [23:0] src29;
    reg [22:0] src30;
    reg [21:0] src31;
    reg [20:0] src32;
    reg [19:0] src33;
    reg [18:0] src34;
    reg [17:0] src35;
    reg [16:0] src36;
    reg [15:0] src37;
    reg [14:0] src38;
    reg [13:0] src39;
    reg [12:0] src40;
    reg [11:0] src41;
    reg [10:0] src42;
    reg [9:0] src43;
    reg [8:0] src44;
    reg [7:0] src45;
    reg [6:0] src46;
    reg [5:0] src47;
    reg [4:0] src48;
    reg [3:0] src49;
    reg [2:0] src50;
    reg [1:0] src51;
    reg [0:0] src52;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [53:0] srcsum;
    wire [53:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3])<<49) + ((src50[0] + src50[1] + src50[2])<<50) + ((src51[0] + src51[1])<<51) + ((src52[0])<<52);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b37bf64f0e7e172c3bcf4b3ba2597aaffcb46911021ace05c364b1096843c1972901374d781f61246a599bf9c44b16352775efbc4bd66c8bb6e9e006b713e43a2546e91beacfe080eb590225712c22df06efcf843e34dad20e6bbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc31de59fd95c89dba19660a0b132e391ff6a65e493667282569c84e4e45b1d24c600262420cb9a8149fbbc3d38a6b8b4370a66a7d4916333e8dcb633a4820405895485638b744d88e0ac536d235e4485eafe3e490692a901651f96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d4b681949c7e56bbbd73ec5bc102c6e9912eef1059f9deb360ccbaa2ac66c0006fcdf430d2b20493b56afa5826196d7e605fe9172760a3a194a0ff3122732b17cc7b322090cbe235e043c4ed869ec5a3448259c5ca823afecfa2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f19254565463d595d01e5b87dd9c4f502389239efd15a1c77790456cc74233b1095318a43e090a760052a1dff8163fa4ea1e5ad2d88260c52118319c83e478afb26a428cf5a063fff1ddb258b0e064490c19c5dab4eed0193d2a60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1492e4ee9f4267f6a01a52b28c44a6e9d7c850dc8c6929347aefc8f364f60027faa2536f2c8a46745d733942cf96f8e6867753a8f0e30c8e08c4d3ed34b446c337f1b782da34f3cda882c178f02ee8965db043fcdd626f89f435415;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55b20ad93a0cb08cef9c0d80d8e7c3e2e77a59c601523884cf197b1dded42526535e78717d6eef3a37d52b9fc8322e7ced4b54cc7001bf60b4bda13670940bf9a9a3d9dcacce12c0eb22f174ae6a595ca8492c24ddb6cbbf9b7abf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4d80d46f3021aa54101327f7e913f986ac5b5bfd612437f47844cbb429cf23ee9cf4614c8efe06a5d25e77106e0f38f1efe2175cb880ac2a862e25a81f3c641d8931946e52d82ce9f5c7f37110d7ccf40e9ad19ce01391f328566;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h833b7be8c105c1a179af5b04ad8f134899458bfb6afc9c9181ea07548aeefa6dab1f86babd46ca94ca76c25b93dc7f178ec1ec23daa627941326bd456ec5916f19c49d8e6464ff63ff5e14a35e869aa93655b5ebcc713a081589cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1143c04355d97248167beef1a1b4e099045cad9d06b9587b1b698535a64c8c9e7c56c612d8131d5849aa6ca2a9bae9bb919d8f9b16a921180c87716000df227f5b71f9eae93e1038c7ba058ebfb2c64b30272c913791d060600fce4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8fef069d0c7c2552ef1a885336fd7691b5be66f891c56c5caa9d1f44d2ec50eea23e6203388eb4c984c27de47e291fc09954d9a1596f2675b279eda66bcb00c3b06527354494bdaa6530f17c00b0fdb427e0ae5393397add11d5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he35e80d4f78f23218d4572f1997f91a6944d2dc9f29c0790b75f79627021883d281cca7d60d194fa4ffed5fbe2601fae127a498b01963de8a020dbb9d83ca255b8ded13b4de9fa53f9ccd746a743e9bac047eb1d3f48e73c826180;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h929b497aeb6dc336c05b394c5bd1a19e6a01af71c2b6f1493de6af33dd6cab33956ea6704bec71cbb0c172d3de1bb466861e01cc11f3f8f54206beeda0322fed0450b0c5e5afd73c4a0ebf96c39d28e22b0f5ac33ffb764941067d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8910fb392639e4f76fc7464da32e4d2e9a53f59d6054bfd6e31ed92579651c666efcfa198c72fdeab1e0a97517393857909d79ad0eaf646432c3a17c85afeba2c031e663e82fd35f04138f7ff962aead6933654112065f71abba18;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3222da3b0832809ed767d556f02070b82f9a8d0a35676685c696fa8997a001c71693394628f2cc14aa893727486fe8e0d3726fc9b14279ce6d8ad1deb5f91fcf78418f173faf1ebc5437a309ac36fc3a11980ca6ce352c0aa934b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79c7907ee0d38b3e4be47d4f9aeb9fb6fe6b1a8f63ca42e21fb0284fbfad08da2b7de829996ab0e83646caa763038f6a0a0185467921e918ee4569230459ce1ad47668118ce8214e39a209a1f3e60be0ac151ed90a16fbed4da160;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ddeadbf449695ef6d15d6d4d8429dff20269901658dedb1b899bb7f7c69694559d5382f482f2da5148045e7f3940af33c3d3dc3f5a7160f6c3a48debc49a95e5cf6f68ff4b68e83253fe072b94219bc1ab0409ca53288aec1e639;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1adff73b068cc6024d3d79310ea3c8d1879cc41eba5e3102ce30ed99636d28f360e705e6e66ce1d87fc8038093c4a655cdd5f0c7aa3b2a2ba9e14b364be9a68cbf768b112902252a0ea8ac0406ff31ab7d70db25b378b06de336e1c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8efce97182b2b0590b8d6b98e26f34fe0b8e6e1f66f6d72383eeeff8b3fbbcbef6994c7b36e77b4aaefcbecf5d09bf01efd864e09586d6d5065d141c3cfa843c32cdba0ef0b74cb87a2946ebb5537483f177c77adfd11b06f47c5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffeb5abcb8c7b82d17fb02eb61c240be793eb1262911e113bfdafc1bfaf7a49e69b80d700deebb9db98b637ce183eb7ebc75ac3823c7278c8264e2152cba17adcb33c8cb6d52a0fe72d1b5dee2b6ef392328fd02a9cbe343f7bd53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6fcaf5717578bca3738a50564c527647743cf3e3b98d80886754d347e159d3f145f586c9c500ebd15b61d7d8953aa607b0d77668c7b04f2635f44f819127e7754b87c08100d34014bdb2b1dac9257eb594f2afe87e12526a43652f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f3f3b428210ee4b8c4f8af1c2a7209313120cddd22e13e2f0e8ab849d3ea8d0bf81cc6a4f0c64efd98f0903ebf794994dcc025c7efe0723a235e5e24694bcc08dd507e7cd6c4593e45e5b6009f6101203d529a024d194735e2cc9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee6f8ab5393b1b7ee75d2a564fdb380ac2ef107456f6e4a88ce9382c2493dc5cdf66e473edd3c7451a966ed89acf83273645c0d24d6069a0637618fccd35b6168242357144ffff268ece79b5ab9313572662ac2176482ad4016536;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c82816e3e231e4597068a71bc4c869238564bf7b5728123a6ae4db79e3417f567548378c3a5901e6015d75a6c190b5d8b20527fd8397ac7e3900f44bad4a0c6da1fb8eb5157068e12640c446193c7d4c463e42913ea8f9e09ec141;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5a491649d93d47413bc8fb2ddbc1513e25d9510ce7e814cb701876f2fae28e7f037be1aef63eb1026f7007b3ccb3de3ba20cd9ba927bded19c6e74afd7f6f9c454daae1f1c9e608f680144a1a4d2a7e25016f0a332105683593c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8461dd701eb2f59609e0ef1a9d0a3dab679a862472ed722b9d6f7957348e015bd5267c32321936148ddc73b256eb1d2aa6e8405cef0b4f0d41186f89738e0506185e09745e3bdcce1352d29fc13eb862c46cb103b8da968179054;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h117600173c0a7776040a793535346ce61a5cda1256cc5d34f185c67c085606d633a573b8fd5fe175d8e15f47f5a4a3fa196cd913b13f9fe73352e76b937753400420e43615e1a4ea6b81df9b6811e446304134f24f3863d827285a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19550ad56a3f0996f89abe374b16db5f331943623093b15d669af40327ab6cf887884a3c21ef00de5b744787ed6a872529d3d53e3d861cc2d369eb2ba63ac77fc3ec1960ea99298c3ee5ee0a922f976b9e50e497086b49e7baa41a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e512955edc98ee59ec3bfc97ee9243ec4a38af70fddc32eb0b331ae44fffa80a12d54333265a3814e4fe9d6841072cf83857bbb6e5537b1cd0d05e1b230b4f88928153fb5c221505559132a8a070a256b1c7c059cdb18936474d3c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188cfa6acce3adab19cb6a1a01b03b3af3ab3843952b0a89d7489d4e4569294c804d06cd7ae1b58bd5cb4a006b2f8c3a84715f3fa93e22d9116b6ea7ddd242475c6a38a019d38e85f2e86221d7ca332ca9d525a7cfd458b6d8dbda4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d38e109e5497e03db7bb66880a5c153d9492af9377f53180c0e43aed2fa2d7e2cc8b072915aac751431f2ab26a2aefba22fae6cfa5b583d7175cc67e84341c1ab29b245479c5ba33cb5b8364db0f58d04066dcf3f09c593d868842;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f05a2c113b43aeb4967d87e54aa1ddd653c2be25d2687e9bf23eb3233815ecc4ba3ba54c7fa2814aad674b6ed978e83b6328ccd898540c70505b3f421e7a3f183375f15d2202bc07a729a23f3eb425b24e8695e4dfd2c16bb64dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1486e6243e5f83a8bf382ef45dc6ecdbd914ca02065349c4d04bc48be12cb81167ed993561fd0169c583ccf69674431319607dccbc03fd21b8f56fbd77c01592dc8a3c15f756c8bf6b3c189b3b0b147ec769e38de4eca0d4114b3b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1020e85324e0d35e4c90177bf6663453c72e5878d5a858ce1f3661b9d6f5557a336dad37ad0fa5c4a0701e07f5dff162fc69372a82dbcd4f4d082036a130509c3508e3a2b82e8cdf31a7543074c3dda69db2dc0ca5938446da357c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5af8314e50d2ed0bf32a787bbf3561d3d22bd5f7e3e24c6764ca274e001bfeb463bb115356b2dae7563cfed5e0e6000db91b8505167ac5d94f5efe393d0803d7eab9ab5ddca74cbdcf8b08d5ee21152246c3c78e13aae0ddb0c2c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1128b5054172a371f8ed59bc3d5c9b330d0e703ffd6a70bd0598d823d3db6b94fdf29e2244f4bfb29797043b7eae1cfb708d79df2494c9a08c6aad4e31df7c2476cbfa9b94beb25866b1fa7713c655e9408f73ebe9f5bbe8a62fd44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb22cc9b90213be3b28192bcbde3699c72e1fa75ac4ae078a7a57d74f2f7665577e3f9cba927c51fac357520c754de418174b262152c8ff4ab2b1490dc5b8771b9527b630f863df2fd539d3500c36aae2dacc6d6583c79322bcb8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16991de49ab8a3bb0254465c026f9cb8fcedafb7dc47efbd9ed55a769cd42d237ae8f487d0b8b487624f66c118d5357a9fb2780ce199e8a7ce39c727557bd41c4c10bc00a647c0fd90f3887074e2c1438610ed506a7a05f7f304d1d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a24070dbbed8d19683b65adad0693456d6ae7ed2176276479ed02b709b01d9398024c37f6135e083b8e53c83e0cecb92308e28265f404dae6455819d85ee5c0a13c5f02935cccbab09b0be1c4301da0c6928b754f83450f7c3413;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc5df20f1610bf4d0d21c0bfb603d072f8b9b64241abcd1e43fa1b3bc42ec7685b3465d197ec124805e225d1ffd8ff2d55b1020c57b2d33010e9feb31de025a4c7e48b0c6275c0bbedbae92e5a4fe24280a330428982520d84a115;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18feef0790c6df8855dbde6ce36ab56acf3fa9e904390369c6252e4a6bb69abca779fd35cb2a9909b7f5395d674517e297341b4f24aabf116a983e1ad25ab9da9317eb7aeb377e7ce96bb939e2e849e97d762433303ef48ebc4175f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7b0304c6efa256dc65ccb6ab41b14182b4da49fd177bded67d5be22acd07df7f2698f7e1465210f3a9ee990c13e07434e31e2c2be5d13a4b65c85fab458bf248a107e4b68fce9407c69e97bdd6101f00b4d10a1ac9b132f20501a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe92a9e3a5de3b6f3163ad214ffa42f18a1eea4e7ec2d564937f150ef9b98e42e675b8a767edf8221c8a9591d311cadafd372891311e55b0e59dad0dc82bc0a18f7fcda9059cb035a6c93a5d955f1c0c2eb6c9da1484a71a0208b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd7e17c1f8b5eb6fe372dc17676f1c8238bab4c950856f74e7dc81f82d9152e6467568d136fce76ad8c817e97d3d641aa91b7b4d10546f3e33bc743336affd0030e8e0b9fdfad79e1664d19a6bfc28c488e6796a05ce75b36f38b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11077d6e5e29c54e29303073aaab83381940c08f32ebf236c5be0e801b03eff9a34457d6e549ac410ce549aede15c2687a1ef72478c9f1fe9a4bc051a7cbc504647c91d5f6de3d5a9177b039d02084ba7a720294dc44469f1b4b15b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c457cc9b0edc16bd514bbfa74e18b5a24bc4bc0d2baa0b29f610c7b29971bdf4d140a619181d7bfa739465a929303d47e59f0cc0dacd0d8a40b1750c25e4fe9a14af1b22bd5f7d6d87c117df13902ab36f134afa69b304c29d9276;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f16e54cd769cc357d5371c923176deafcdfea094d7c26849545dcd156f52db2be5162f1ea79b47f2b23786bb1a429e4f90e124ba6c3137926ca6d4b51f7335a718208900fd9ba7c53ae058c2517ceeb3f3db6ad12ed5728cb0c8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a2ffe8ca617c1b378f0d2b82971d6edd873137b1b88044eb38ac27943b60834b13bbb4a6ada1c0c0aad5d1b76842cdb47179267c181a3f9a28cd48eaf9d15b3ddc79655b7b6aa5283e5fa66a4ba7b4c5b6fdbfcf4509e07a58311;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc193730435cfb4207ec3ed8d6b08b73e9420868c6f44572c729d2ab6e44fd4bb69b99aecffb2e2644a2f09e40a8562d55a5b0b7c83d022b023e33bf73cfbf37dfb7b3f3850eb709b57c19adecbe7ccccc2318ea79a4ff545669ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a06097715bc1e69f561a0ec189bef617521d5ac565274bce0f6aaa049f9623186fc486dc80d5e2c4968fe587dd81aa9976595c40a9b69a5ce0f4c6c1cdad4178ff336a6c32cee882103a83656f5621c3dab9365687713eeeef488e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de2a0930bc8c7b267f777665460c610a48b0c392dccb981deb02b948a32e9aed5ad5c149ce64ffafdf187bb0ec2ed3ce65573f881fcb65f4df6295554ce0a92be29a81a9364ae9fab4a64fee471d7be873e30c622e47fd370708cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c807cbf65ed594c355ce755661f4031731a269fbcd8ba8ac46a972073743d296939286650e37ed8bdbfb8bc153f85b70a253eb88e94531a61f3e456b9bdf9aa9b9c4b3bb682019460a4e1652dc6da532e26d5cbfffe9d062929b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126b8f6b367a2bacfe1455a7fd58098b7d55759195bb48f72f5749facf0725fe46c2401fea5d8325690151e2406ba320893664079de9d9ff74f09ee0e19ce1e52d11757c4e318fd9e5963619f9f572814025db0b00df2b0028f6dcc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2b69f851e9c06df73e31764936528071603b22759dd00d6c6fe3ad19eaa510976fa0c87b76d59cdeb45f01bd865969128e881eacea9b14e00178299db21a4223465fb53351a9dd4a326d1a06eb471039210d2b8961614d8ff43bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121271e177bac44836de6d2d010433502d3c6554a18ba36871af617988101c570613a01ef567a6f13dc2fde0b87976d08a5ea0c06030b988a37751a60942125a69c1cdbb8ef0d25832ec14158d1f08b2a8bd74f221bb0eacfaffe08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h931a252e1cd3cd76b40f5e5e68304762108cdde71184b68a72885b15fe94d68d2c9aa793e56c1a56e472a7e2cc62effaa6e78a64ae649a8b0484d6e5a96a8161c88e0236b70bde68403037bbc09e3fa261f3a54bc37516e72a53cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee8568875545abaaacef8146b83d36738f2452581d08586cefecfcc7a88e26ba374e620c4a4d81d3a04a39a0361029cf370c868ca8072bea226f1e3367d9d48cb7984c93837756869d12906065e64f4df82d46d9e2ec185a08582b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67129178e2322ed67907ea762f5e309fc7df2dc02bc6c2a593c45269d444faa1f0577b65e9c20197999c76ddfbee5706bfc29e53aebbc0b2fd4a048eb0843428b8c2a1cf1911042ee9bbf85fe6935de7ba4917d9d5dd871fe2796f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190656cf66d4c0febd972f7106e8f353837b19c8c20d96907cfa9548d7d65e5d0c326c61fb449bdd4a23928bde0e86a45d80af6f96b4f551feb84780f412fe39c57cee5ac78baec00d020c633e70b69d14f43f22dd082a4e4aa2d8c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5215f32c6e938275b971791942cd6658c1cc8c258716eff5428392ad61a1076d0750c359b69ab45f7214becf195074d2d7314425cd3a737e6394041a4fd8bc3c1de147d1dc401d66f4235028095e92a7ee4195f7ab2a411ee7e9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32c53752714412bd7079550172b55368e564afa735982d7f87a80e13898e1eea469d137365864240ae25557c33c2b49529da9ea481c1100a6e326feb01e2b2ea10d6aa4b9aebd6cc6538b092fa41d4facc40a1b049c1e4b11e873b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187d908de8420d63470a6c73fce78b6b5f70bc0fea844ec8680d421a18a3935ae445c81030b0c2e0e69e3024bd1035a6e6f04f59f09918b6342d5b7560f9b62e06336c94b5930c7536c3a5f9b2ad7ae89cd5c78ba20d28318099c20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3f6499133bc3969c172d6359d5ba3f1301e2c213b9bae0bce8801b91773505f7fa4559f71d4f78c2d580fe808c35426a9c82bcbe89f3c288db3ca312630bb4bd531cbba7507d3d1565ff2faa8e3745ba9de60451506f81f346aeb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14799a4273ccf0aadb01094cbae049ca6e8ac08a6fa617ff737a6eba12e1f6ca9cf84a1ef4386a6f6b882e8dcd4e0799f856f7575f953a81595e5632fdbf55908d7a0cf27e304d11714f4417426e2b46d4363032e438c032e3c97bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af037bb6acc8aedd7f5e1ba0a1aa566877da9171ec1568af1ebe5562f0964db94df46ea8378118128fb7ea88c896c256d373f861eedf24f7232d81d42e133597a933667c3b7d02c2a0d8d1151cdbfb2c820a27064f14563f5eb026;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81aa912940311ffa07f426a884d94495177d7fec0013561352e7dd181f16869352f66208874e664de6f973d39e402559d46415ea61260699e46fbaab3821146f942fbb24b495b2ab6360c3dbbba0117f4ee9298fe76528c5bc3891;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1204cdb1a5a5ff7d52dbb2b3945d7497bd33f7662fedd8a1f1b6667ca94ca7520363d8a5a9b0600e4d216898a25b979e62c7ea906b4ecf1c3986a7ff83a4d427a47a3f50c9aca4f3752183b7a5f5560c5bf9f8cdf3cbc211794027e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1698329f08d48be1e424b3f08917ce78f95b98a4eb0540e7b4335193bacedeee795ce970d19568fe6b158388b961fd1475c20c0699d22e86a290b8a47606686b562cb158366da3b6edc2e9572e27f04eb9aa2b788cc00d1a6219dfd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa230f0328bc5ec1b29b160d0181b859de2ecbfa51218cc49367b5dd96c7d731f3d913ab8bb277a2a02337b254bec820f0cdbf3bbfe2b9ba126762d812218e72dce49a21dabc8e35963f92fbe9b6f534539b91399ec1a26097f7ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1304a92a7b1dc8da3077884ea0429072f726f57a8f5096c6dedbcd16aea75b59aed4510aaf0a329c7efa20d94bd32c6f59368f97460b1d7ab2da28dc677cd61e55a129496d36fd25943652d3299852d591693f5ab2fa7e859595e43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1992ce1565f3619677cc622d2134c8689c109e7bb7074e760940c28a2a7aa0da557acb24b8a5dd782d888c05cb3da7a755bcea5224a295e8651a15f9a4e08db57622ad35377a1e90d51f3921c8161301296e97f998bf54df376d632;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h984011913ef3004e1ee88b8aad57928b7a44d0c08e263da9c161de456cb3c3b17bcdba06496face3566dedad7ea201d9106449132ac6c4882081d7348c8d009098089039113624ad6831d4b42281b9366fdbfabf904a09285b1dc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1040054a5cee7157459be9d0275a9cbbf8fd9490d99b7b7d46a789873694f38ca2a321767d4b0e0563f7c60567ccfbcc99b42d5f6d879d2de72a076e5b0edaa2c85fe3a381ba07a345041c3649ea15846d936a3df4d8f77367906ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c9efa0e13c56750f75ee46e08e0fdb487dc8d9b04ff755fe3ab1507fbd52aa94cd8098adc5438c5db80520ff1c6e2fffbaaa298c88d8369ea7b8a24d0175378208c160096c9a940e1274afdc291fd5a2d0673bf677d4990d579b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc2fd1bf8bbc30a3f0943ca6295174fdfab259a1c9a81c2914254bcabcaef0df5a224642c0936fba789275cdffc3a65bc00a19bdad359449732b44640c44102a21ae432db06525f66847003256b3e9a3ae4b05bd934e3417da39b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9c24207162158c25ef421a5450b2e81107aa52f31e3d8de487ecdd9773ee39ea8ac4b9e941c2c3a2f63282d42212577b5485bc856fa3945582a663434cac0c5f27131a091f334bb2726df6431e29e9c2956d7b20039a4fd208966;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f90cb126adb0f90ce1d5acd07ca0df4c93cbaa1b028205b5054054b765b6846c183d90e4e44b4c36c0f87b3d459cd9c51c135f620aae6b7cc9ad6b54d776c0d7345c7d8dd0e1e116419fd28373113ca8569c993bfa601ac40e2531;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf647d74ba3924dd0c8307429c0d37fb537ebc6d7b946e255c1249217faf4132f87687afb79aad8d6016361bea3b0ca76c107af4ab436f85ef1914d649ad5edbec2b93abc305a6cdfe7f027f2487245a0b06933e12e9c9aaec2418a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcff622837a655c4b9d0e97885d30bfef35c44a5468bf34f5de3096ab1ce0dd3c04f9875787a5090c931bc79151f752710bf9d43dfb3d5870d71d88d93703efaffb339ceec8663077989004e78a343699147557403c72b4536cc81b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122b64d20cc5b508eda6d4bc1280f1a8666c701a5e3db6da5230e97026541eb8d7ca50ebeeab417126efa0a62ba11ade08966e82a586b6f4afc817881b3120b7c04545d59723d4b76e75a5179eb6e994da62b791005ed1edb15dc8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf17fb3ef5630ed8e6ebbb614dd3cb7965e2dfc481900f210cb4860d5395e34acdfd5bb1de925292d40aa2d935ac5359ec114e255ac25c0067ff443eb1d09cf0bde576d601016de5849691d6859a1e0962d0fdb8290c20338aa05b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1049b325d427dd1658fd7fc34e569e6422e78635766b1e7d95a568a754bb8aa00d9ad3667dc3f366a7c63fc5ed991af19975f36838935c9582c422e3dea3898e4cbfbdb880e23ed06e120254ca2225e5402ac6577f3e9082fa3de8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31169b908dcc2a1429f4b97adb5173a58fc3e9100599e1394d8f8c97e0c63cc9c80d1af0c94dbdf5a3003acbbbf28aa56dc4c0adfd8d905d8b447b647a9af430dd3aaae1c70942ff08152ba338d347b945f0be803c75f97244af0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16924d203ed95572e09dc138362e9d0d81ac518a16aaa3ea625eae7995f52f640a3a45768aa563686a1fb5e97c36314e07e2b56c8544ea1c177985a7500af35342a04a54594166c83aab5f758984c7e609f206a01d192aea5cffdf7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135d492c4ac722d0a42d516cdca6006e8e36f1f7cfec12577a1bf603da620aa02559648124637c459b29269ee8de496a0d323080fd7f15dc0ff1d10237bfdb52033be04ccca99f5c1b1afb44f3a1716d00a79c166ddad09bef8d610;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2ec817f61c3aab2352a252d4f209c9fa12d2b59f779572b78b72b1468816289ca2e73d4935ad503e04d6f04ebd5977a59b0e79262a6a22426994e13df9ef9f03b548c92c01ecf7c800f99cac1ff481e40ec7b985c5dda0a94ac0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0d6ad2eb5442ca7440d1c8466c7c24f4bb7548146534ae7ef101a892c918579e7301b43316a01e0dcd3a504cb28827315172ae9fca5ad44f615dfd371d959df449ffacaa7c9584710cfb25db778b1cfeab4204bf5e70d66b06d74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da5cbe19d93734afabdcaf6da2bbc83fcb42c323af4757355ca5828ce4bb4ca0f2035dc30993a30f169576b50a477fa23ff03c6d9073d82b9b2fba11cda1f10fed7efdd1ed846af18b78080b91134e962a079f1734fba113b9a7f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbb60460beb2a2f73a49179a11b063083886d1bb149651abbcab7d6511c9c3b7df6f6a9f4a488ba02b071c5baa5c9a2caebb5dee02c0c94079b789e30c05d52933d8ebe0a199680101a63332e9f952289a19f41fd24ad40aa62d09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a01f18357755cbe11d8876eabc6963638a03978ff0fca9ca8fb1161ae9f4db5b5cd888340324acb8cddfc23b3bc74e58553589bd0bc2de3acf27d385f5282ef2a3c91ae4629b2725f4a40aed464148cd139530dd2c9dccfe089fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ea3c367c2c15dbdec2aab4fcd9909e27505e85b7b3f54c83b72bf7482e66387d1d0d0b11792a47f81c2428dc03e0500399669955a98d9d21836e1a17ab7f6d0fa05a078c08c19a0ce36394a2cfb521500cbec97d51f984d1ab532;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7585dc654ecfdd8bf7b4c92077d0df8c46d2cec806cc2339ef3b65ffe6713fa96bf57b887c6cd3800dfea756173094ffceb462ddfa4132f8deb6e221c05e37309a9f21b689032bce22252bb559138eb3e9fe134268d84c8a3ac52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd610747e93c047cfb8863a4cb122b4bc513b28aaa3a07d3184e246f924f538340a851a530dd96debd162e949b96c553982867c5730ecd8fa1aefba3b7d5dfe2f1eddad1d234075e1e88322313d69bac430e1bf67ac0e1cb5a4f5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8084e59901bb9c5f95c2ef3bf1164688d2fd5ef05671fd26abc2f16d34fbe88c07256ce0a40165e1a0017615b59edc181177bf3f903d00cce5da1db6faa056e3d693d67073e29616994a7c9bed690bf522dd8396d72b99aee78d77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a9d40472fd25df3413101cb5d21a6b54b110d58fb4befb67768cc04672edfda352d5a6400901641721a5fd5c75e5b26b075b64df45d2233fe9d62d14d864e23af05a59c941f785bed89e4cbd9887e33b0a3a1f26f443c16cc5ef7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc16016b487a502f77d7150bf09c47d2165fbf20bb482612e54eb513233d726014a3a02d84a3c8ac4820d6da3213405d4c9e614aa4dedc40809f492a6a543c3e929af4c5a4a07928cfa8cbd284e496ece3cdec053bd8b387258ed0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12be695bcb916d296aef93bcdbe4298ca7d1e290d1ab16c1a5ef93d76e079a19d3f745f2e5575674c1cfa3209c79dc6ea2203f65200061240b2afa55fb3de64185aed9cb46d1d4db0bfa8e9f62037399481b1313393c3cbc1bef6a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbd79e13cefba1d46a4b6b465c32a5d70a785fa1ecfc8d2e8dd4c546f3938b80b20145020209b4a00918d445ef6bd6d1e44de267e9b940a79c932ee53ae23dd53d07ec84830484efe4674e4d4c7c644346fa7d51099451fd70c92d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7dbefe713a6df35254cb0bc38a19fee6a46704cc4f58517bed6eedb3210d1ac7e5f47329c2c6460f666a1637491c0d6990d64035280cd29cdbdda6ea2a76932ca99874cbaf26f88b0cdd87cb14529e345ba1c9a492749c3ffc12fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d24202407a5d4ea5f4422ede080f1e009a0b042ac6b5dc4bfbf15468318a39db5fbbd1cfb2b29d9390e82540424706524f61edda56d0640dfa7fbda78eb1ba95a1875cc799f01b940864a8ea24ff1e5d481c5f189d39b66eb81c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa001d76469fa453476063f2495a9308a90edb62f77cc50932d3d4f04bd96bf5898014946bbecd77989f44647da97dbef3234841576528693e98f2c939ddbc26ef34c2bbd76beaae745473bb54c508779be25dff8ac9b162d6e76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194f3cd42d71bbde99bbc426c246fbfdbfb55c600f85783e618543463764d16d634168e3d9e7334c3ae3760865e02e68ef927bd3444ca5269c5ab7cb8ec52bf63c0d099a379e802d3104757c387c917253b1282d287852f0383b0d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9689dbb791c29900c21b16d42532cfbb05b582e99814ed2db2d07fd339e584d401722bcbc17a8644bedd1e64c8073cbef1644444e3cff6c7ce6641e31bc55a9aec2779425c8bdaf6e113299e5d4bec89c59fb4be9b0244bf9d5c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167f60364c824783bb2c1381ef2c6be6f2f9b76a6851fbcf64765caf310f4cc8b024ec0b331b0abe4935d4d824ee8fddf24b8bd2a38ed036309e98e7de053fc4f4328f8f6af45cfba04cab884d2dcfa344e66d007409a8d49276f7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd327ab837722891cf55352ffddf072ddcd85f8849106bfc3a5450b51e8e3a244d4db971afdf361af349d56132321e0dd253a26619e3ab5a8f64ec4d87bfd31d4790c92c2c04476b4b5bdc6ac11abd49263bce77ecd71ca7fe6807e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3553595d85993ad343038adba56ddf8f2182572dd89bbb25534e1ac8fe274e59993506dab4a43bc4bf27b20b494516d8f9cd88071ede7759d6bee7c8d1e531527967c8f4f98eeb52b53607e2b10986d2a6c2342018bc7c25504d3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ecb5339e7053b2a30fb99799bc1588f021f2825f030dd027bccdfca1e940c14be76df484e6eb3ab5d3017eb4e1e4577bf4888b0a52100554e7d8fa56035bd66d071a955667f41c2546e0fae92fd21accd91d23f478f2089cc805a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cccbef74c30e5935497f4fd45ec256adec88d9c8db0dcb45ef94df18c13446d9eb4d6857d489da0c124d72edf971af7ed2ede5bfe0102c9fd9c16a06c7c259dd90387a49d5ac382f9e2c1db53d9dac755a07d36903f38427a71b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e28c146e52d9394fdd79185e0f74bb32681e47c0f08cedfd401a14c5ad29325e8f962b5ca5d7582f744ae18ca6df9d1b6316d1399169f0b2ae14892cdedee96a04a4b72fae62ce6f1d760b86e0f44d6cab9699de17fd238866a38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdd769cb052d13a0c6f2dabcb174f9152e4c80aab3a42655907872f9fffb679120f58ee8ceacc1928bdb92ff08ad9bd066d39f42686a11365bcd0ef4219e9b2bfd450cc61d621391e0af5a072981be702fca75fb652981a46e3a8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aafca16a671cdb54779bb10bbc61d445c614eff1aa1b9fb1224e69710a70b11d420d76b0cc7fb144bc215715ffd272461090703ba8c9ad9fa6b76a09e38424ca1259de5f1c2d56f66587ccf2ac651b1d1d586055fc27b7d3e05c01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d466d05768d11d54fee2ed06381faeb175574a88d3c7f31eaad81fb7d631b751733b13839f4409bbf0853239768681d4531e6473f283122b6e92dd55047de59e406b32061f2a5435c30423083bc2a7a0f01f02c349c19077434a56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62a5dbb8af6c48313286b032ed862ac1ba812e14736ea30fc4e7846f6717f4315ca04dc015ef47cfaf4ae6355795ae6cabd1277eff28b3af0384e0645e1e4ead63b9f75fdca647e0d4a51250e18f6ae2ef2a51758c772c7e9dc07b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb179d99ec4f0ead95e616e64c8219b439e02b7223610a64c995600902214565cdeafc4fe74d9ea662db08a13301b6b8ff6aa9baa986b31b8f7989d3e45d544277901951f34372d9b901cc2de76a008f777fd5535ed149bab81236;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e7102e73e98c457ccfd584b59a7f0dee4920f92ab0a9eb25e993055a103c5d6e4e1c40cbb4f623150d32219dcf0bebb8dc6080de5d16d38d7392a693c7489a9db963b84d2fd62cb8ee39c934fbb10adaa9d9f2d60ca55e3b835d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165b5139696b81a3df1e284cea861df30ecb674e4d144a0e4164f05d669c30e80ed535ef62cef63a57e3a605a3aaa62aa16809d75ad209888423c86038dcb027c6ec30606f04cf291951ab9a276d468249ae9b9ff0b5aae8507ef10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d0b123c7ba96f08a99292b9e454e7dd8e0f90e8be415dbb983aa79611836b1d5ebb94bd25f1355508931edc571d9826afb9160923b8c81198d58825cc523c653701c88311659f537b0103f87c25d1ae19b278bebec0ea9aabee13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1161af6a34a4c7d21cd8b282bb550e3838c553c832ac4bdf10e61ba70726b9e63d222b70f270180159ebf1ee7d19949a49f91c1b117ea301e45c8756969f4c9b52d5b51c321147670eaeedab725e698449d9e35cc2bc5232c686602;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2c75437623ed39e956245a94e8bc83ba88c1f61a629c7e8198601297045d12a98a5201f87112f7ba798c50215caa7da6f92add002ecbbc8f030de23d7fa51c2ff01ab13ab1c1e4c1e80600af19f69f2519c4205876ddcd96361e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bdf19aec0b7f4d30a6c2c4ef660f95ae9cf2ada14a38d3d4973d7b1b5a8e684930e7299ebc0d9bd5f606e207ff26efee484b334c7113bae064561545ea3b8a055359bcea06321aa16d8d834930350b8460ce7431b5583d9b2117e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1077bcc24de6857bd300996333f57bd25bceda7665d79caf48ba4c0d6bab1b69b017ac92f728f13cb838688799eaa031c18f2a7cd163b6a85675bd563feee02488747e219355f54072da5d52eb2b86c50989e80bd34cf34cf13b051;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6799b5239aa9050624b62a00bba4b26670f7c8f6f2f856db0c0bfc555b5cab4c3c901962a0785e7835bd481d602e568ba19bed85605a03a03dfea8279da92642fd5c45cf956746142ff5e5d70f11640b56f7400db637cbed16834;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116b0f0b8f906fe6c04ca2c31993cd1b6ac478eaa2ebf195572823464809b138424193fa7defe300d66bacfa9ded84d1f4c676d26ffa5217e211006862e413af030df7183e68e6b772f897e6a6eae6bbc9fd1d0bc88621a7440a5aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71926ad49cf5b817e609bd0f70e830907af21e50652761bff79f621a11c00a4a5ede4b3ce8c2ffffb720369a855fc603b2a54ac855261032dd039a9908dc86a7b9fcf8db86a22439731bc38da3d536e68ebf337a5a26f483907957;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e9e85bc3947630f05e71bd887aa42d64e65ce12e6a3a757946a3273ef8c2ab84ebf279717d386103f68379db1cf10c5f89f5cdc9c7b79cd377d58b5d35a3fe555187c377e23e72c937bd88a93164e736e646e775c2aa06244bde1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7439ddba529f87b4bb67ac0ff196ebb08bba917c19277d55ca7d2e9a059cf7e161a92b19383b8b091d4fe734b4b21aae2ee2c72b22a3f2df4b582ed16ed59ad6be18a000e292a0f25c493c37cc255810759747df19eb7838defb1f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1643168441d489ffbee9fbfb70a17d5d4a2d602caefb5d8a3db35b7893be86e2691825fe85267e9234623c6325060a1068269ba903d63bee08d25b2b19cb010a0de296035e814629cee20dfe1e80a2144345d2b35258253669d2a74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148edc09c6b822e1f7730b5343472faccba9eb369cbd51ce6ff43d387920577fd8ccf689e8c7f7fea947fb94167879898e155ea14686c269862fee7c25f30c574d82acdcef77bdfb21608a15aca3fd203de2cef7d5b4652a3bd3995;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa943aba11b36ac4f787b484edee5fb6c69800300fb45d1fcc04eeefe6cc70c5784dfd1c270359aa965fd2c866627a37c7292a2538015fbacc2b402eb4ffe4441bab2e96ffcd5f786732172a4deb02cbebd677a395e9767e0037c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170a853486ee9cc5c822c3fc88e2659190e7e1a343d591a95742c8794173eaf73e3b109d67d4ec08881484f8012d94519e9b3dddceb4419299e5004d64cedae0576fcb50b866b7f9007937345985c47bf238a1ba20cf63941ed33ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had2b916b2208a505f80630276dd5a27c72a70c1d51229446e65da60ea5a8b9c566268a8d5f296c0002f348debcc5e11b072e781ac4f6ebb83a7d4813be6b81ffc4833611881e6ff04b1a991c21c18772347fb0c8aef71e40ba4fbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3bce4230fadb39f6dbddcee40109b5397db7d49dcadec002b64c123d23c84999fe005d7e64279377b78fcc7ffabf8d8a18bd0f9dda1c65d7b40afc782f554726111b62c83d4dd896c0350627f3fabcd5c6fe364d372af8212fb16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb6bf6f56e05da206e29cd7be1ca1e721e9781cfbfca185586989a54d1bc1e602469e12f76d5b6a32819b17f2e969988337b20cccbbf5278912737e4389058d3563f66c4f9d249b3d6fe9508663df59990aef83e82e962810fe636;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183a2c8b2a1c2f1c78fa862cbfc0a6748164352b501fac3258080f9e9e05a4b1840b2133ae5ba1685327ab1f89fb771e5f7d0e387922908c883682d97131f2d0c3cbe7818f180e2669c2a1585782b1bae88f7f07fa571decd850c6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cedb2a2f752ab4fa8cb13f20e419479d2f47ea314122303ca96d14e0f782405bddc40ce7de0b5cfab4deaf589550866da856c290e1b57fcdc4a96c80c7fae8a70f71112eb73e1e75888121e29105736267ae55a41e1e33c52d1293;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1975acca0f037c2023c7f2198188604876643f4e474e9126ef2e29b5d63cd474f7561953623364d63abe5b19538ec397227212862fcbd9aec0363a0a7adbc4ad659d8bd12bb9af751c905d031f8d8018cea0c026ad06e37c6799cca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4326d64590377800e67fa246ae2742c1be47dc8ddb27ad3b884aa8363b84635f20bca98b4ed369cc973966f52607852c80bdb5d1e4ce8fd5012f29088c7764fd1d3c06e226fd71aa4a02e145843b165531a7abb7d156d61f92c1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8285b687164a6be2169b96460fd2e6cbdb6408d62e693787cd50492c8b27adaef0dee68e842148abd94bac8cfab655cf612761a73720a1372cc9cbb6f2e6661f571009163386d0a60410d5a5facfb539559e176989bc8425b5773;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a62092e2ae3291820fadb9a7008ba99824c4c4b2811eb2751bb53332721db3e30d7fead2b964e77ff3e1b7b7b61736d09588a39dccc49505eae39a0eb0b56243aebb64b87e24c4712d8b2962f05f5ff3de964f433dd5329cf6b4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bfc81d391d75a4d243a0a646bcbf3e6e3c566015e420d40aa02f453963f859510d7f04eeb330ecf9ff78b89fe347ffd0050815cf7c7a88343f8730b6a5ee6b05a2968182f7b0398f00e448e03ee0e47b9166baa0c2ac6f7b933616;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b4dd720bfaa80c6780e147cb44e2f1b2f2e6f0b2423d8fd3ec305dcbf891261f223fd4304398cbc2352e4fc77ad98f18e6e8bcd9154818f35732c904d6b0dad88e4943828327ff31431de5ef1151ed21817ccde2ab963d12099de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a70ee518e7494e907d3199717e37846d4381acc5aab04a6d3beedf848691149eb327e05a0a62561604c3f6ce66280f13c357b773bb1aeb93cc7e75bea0070932aafcb5ee0630a9c834ff889e07e1b769e9d447545e6f007484d2c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a526bc145310c43270021c01e71841afd59bda7e84db89a03cde7255b575d174de925f30e59cdf68a75cbe8011b29ed22a264b9a41485159270822321a7f82bda5f9c8704a050a2fec29c519926d09d058b33aecaf8189b3b04204;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b314d482238ec86d4e4bb303f6c15d53d68c72c553e1f37508384e41a0572474a3831804f16d2956c30c1361d96bd8fcec5bb39c5197c47d509d98c73866f50019e17d54a0a95e67263eeb0e35c56bfadd3a050ffd297634cd62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfa78da916c10143ab58d1d1104c4e8ed5e66652f618b04f605fddf03208851e51137151788fe7606a0943cd5ec2028ba59055b1f6ec0de14892565b184ebd5cdc3c6e2afaadc6b6b7bd0e876ae906972ba5b20fdcec216cb3f038;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4de81208a0bfbf102f32eb0c21e6c7a44b91048ce8721624f35afd85cd3aea498c4ee3f0e895744273092d6f4ce5936e32ce0590054538266564f45b45d0295b0ff235fc51735678200d8c758c16b2f384ba05e6ae8020f1857bf0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf7ef2c3391d79cfee82a8e28fa74394399ba380d4378d8d00c4f5f86c9c7a85a31e40ca80b5f767bd3d7234449ee52915eb4b5c9792e9c5753d35badb625c9de6fc92d464e8a2e289722ffe45f2c6ace2a68d8b22ac88d2ee59;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a74d929a0f78e927d0a5b8fccfdf1976f91d0f5979244e634183d8900b8587d3f7747feee32d4940f3438fc9c1621b49af8bbf0856f6bdc1225a0debd8a3c8d722e693050664514d9cd727d97cac95993a0d1151df8301fb769d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51fbddc67c2f203db801039f044a8c80ed96f194c84b3ab66f922e609e5316a38d70f6395a516990b7e435904337d10662790d08f81ba1f495611a8aaf0c63fc834d5460e8a36f32334346e103cb8ae36f95538b80f7333dd2a0ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f55b2549b8ad39e581ca2250a1d3413b0d8bcad9f9a4d7a4912bfc4961cdd236bf5685708162c86596a4301f7a8f2fa3664032dbf959b7cfa1633d4c7a4a4f4d5a11c6ffd6fad22c1f1b4afde620d30b83b06a84f44a8f99a2a71b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd471a7ee85df58b02f187448bbed0921530f1236d84e1ed41000c5e39766f965865500c1bebbf8c09d93509ed3430d9a3222447497d4d89f5d37ca3fea261f5580b98fc1b75716b57b88ad93e676515c48ac8d16362934cfaed43e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98d2db0e4750035d2012e9fcd99f1360447f08c464c49d55010f213723b92aa806e2ca610ca830579ac1bd8859ce3ce70edc73d88a6331c7c50b43327830412c9a8ee1d94085080dbdc21a46e66b631867c4b13131c6c5a80a31f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129ccbf5a6f1203dc9b88b5ff1e9a22ef685d71e1c3baefb79b7d831fb71a434ec814942eb9a85f0ac15687a7b7100eb1de5baf92b44802c316c1a2e1da92711c438b79dce56c8a6a1cebae9c82235e394a408dc0fe1f24d445801f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fe642b578ed6eb65388761db1c62b4c043d064fdff850fc6018edefdf18052ab6d658759deadccc6b3b5f5d71d0cbc98367c09a517dd4d8292a061c464f318f79495bd063eb965c7c8d361c40f95debbdff57e6f822a9dba68b41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6adf9d3642eb24ba9941645549b5d368457ccd891f87a3a837a3185e06c273a3ce5fbfc5bbb991aff0d734c51d48a35bd5df08d24307eaef5439cb0c154c7d0d7170f53b951593ea9f8f60828834c474d0430103a420a8ad6e4d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h150145880cb7d3808699c27102cb830f31c10a7f9e9852f576ccd06ee2e4f716a572eb74b5a288a38d4c89f6eade7a155c8dc6fc00af5d580b04bcd69c53a1628ddaca8b1eb3059abe8ac74e1dfcf36e42cf35840893f71676bc071;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168c576315fa45d3240652ebd69cdfb293131666fd566fc54904581185d857826971bb0d2593468f7780789bd9eaefee7e3157a7a1f3b4f783159ac5b75b9ea40b57f6bbf3d4d085a405b2c18439fb9a861a7232673ee493116fde4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de13e8c4d108893d91cd37d4a9905ef8d95984cf9f7f7633601eb865f3c0debb4c890ab1e93612ea34ca94ea5b1651bab21c03e907ac229155ae378e718a651160914fafc432a4e62cdd88a5921b2f6793e969d6389384335a6db2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd15a40dc7f98d7087fa719d586533fed5c296c95e29a9e202f8f3704b62eb6c076a756bd6a05450a870044456664dd9a1a853f3da117d0b89e5d15d1cdbb26d0c2afe1bd8cb7481c7f9303c2478d366312a289524d35249d134a09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10472b027c085842ea10b886651cc77c13206ce6e6154e8e5b8bd26bc9b706c9e0e2945491709f415616283b0a5cec8b2fdb28f6f51cf64d88ceb0fc2c7d68ffd9291d85282f860e885eded24dde341cc47912ec584c8a9928f540e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111a5df281c89b374ee3ab6f11084b73e429051b2360e5bce2bf77a72aa32de1afd00b859828b2dbbcffdb22b28312a426f68784fbb976194878f05d75a8814563533102f366b2cce98500cdf02ee880e941966020a43e462572196;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h582618d5a4fce2a41db2a68c85cfa3ae45be36eec1638dbee44ac461f5e244a79a64bddbe4f41b2e846f0a53d365f0939fab891fa6a11a66ea6af7c29cfe2d3c12fc789825a9cda18dd4a0655adf91416e0e30e06b07a05622e851;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he619c69274056169440e60618815afef2fdc62b93ad61faa09c138464e4fdbff23a834d3cd88ef67d9491362989b39107cdca36250a43f56fc8dd6d1d972fd8bd92e71eec053edb6e9a81c10436b8238c2456422c36b206f040217;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7654ca383b0e2c6aa26e5e8efbc722d49ff146113e45dabe99a8fcdcc7a062906be69864af1d7f05818c7305a5417b35b3c3398d4f8db4aff8114c898d50e805236ce9ace31d960a35762f4cb52cbef450ea59de2377f3528dd3ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ea86e7baa71e01c321dcc1e39f83c7e6d83faf5498186875de0da06df201bdda4dd56c754a8103c1dbf841430e2db6d68abb1d8fd8f270439970969044f8fde807e10caf28cbb559c1ea388e2826fa9438f71ad1b70468dc93059;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h602ac1b33d55be6b12d3ce2401a7e11ad4fff741991ec6a714e8f17852202a48e2c1ffc4f8a4130c15eb7872144b3048d5653ff3e73b26a835c9583060e70cf32bebeaa9af9827084d4cf8524f25e8a2b60999e93790640bf8cf56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ccdd07fd5b61c00ddfa845602b5c9fd7b252df4529cdc1c70eca3247fac444b705221a9b9e5cc9d3c678232bce423a077dd3fb32aa94e7a14a58c2528e526bafa259fe8d716d524ef28d86294d25dd4908721df18ea48ec62dfd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d123b902d6fc282de0927f03d5200ada74eae136cf7bd0c3a91990e7f698e7a1f610d33aff6296c0d0aa787955cc7fd30576ab650dcfb88948a874c702ab953e96dccd170b38a118370442cefa1b84414371602bfb7822baea678;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10947799bce68758d0e4c1586a1a8589cb1bcfd3eb996212fa84905060572fd920f053d1ce3f32026398944365132b6b62f7390cd30924f1922f25851d6812e4edc0d4d196ca7c664c0302ebb9ffe4438a20e5227454a47a136b192;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e260ac6755bdc346f75d0816fe6b704b0b04e6515edd23084dba798d47b71e3f63f8d913eeee3a3683f88b517cc94b5aa937969fa63e99b28cc8b2dcd8f4450a50d94b517609ba437414fa5b92bc3d8b9d38f550dce26dc69d714c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f59ac91104823189b5ef9927972a68d6919790eadfef970114062f929409baf3b6a3865467c5a4196f20ecc01dab1f6f959c5daf9a3b7e14056719c36f4a2d0d3eafb04ce0e2d8f7746b567564bdd0aad69ef3e034bb5557ce9e65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaaee4d36166ec2a6a310ccf4972723cff89bf45357ad0eda2e25f1de9db63f68625e9c7b928f7f6a2fbb7adbd18fce2b5704c00225e16a4726e3d71320978b8043531f6d71f823320c48de34d4c3fa646c8b3b6f7182254015074;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4c05b7bf264571ade80595e8dc16ddda6599c761309a79ef1af66d80708d424730d599f981fcf88f5a925260b8f99fef45609eaa5f1809348a4cf4b62fb9518e9f4da85a58699d70fd1fc25119cea4bb89ea9071f36c280fd3434;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22be418c4eec6d14ebaec0f82247e6d39c17d94997786ebb7e33a44850743ad73f85fcc4c85e8b6bdc8fa1f83a968bcdd43e33770c4fc3686515917f5520f2b5b5a349d1cb3261c0723731665ebf38037495f2b160e8c33f2487b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d030db6273eb3308138e17e438086d7cdb470e24ea9bdc6a858f60446646a05329a9f6b22481308c62c39ee1a65afd70be5dc87fd576b3be0a65eb93002aeb35818954ca7631e2e4c184b2083a2aa76e4fa0f3be39c697784f16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b3652e53ba86c026baef9f7334862276f45fb138029d145acf17aeded8d3884e6aae93f145f73efc8cca9210598d4c09b7c538d91e3f7adcdfd5b85b97ccf3f4a86f40a1c4e26808ceaf449212000e9a38e75bd935a6c6e28f601;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1748d70c1b2a1c3d7af6ec0763e1dd2faf9769da3f05c2b294f1d5436887d86a16a63ecf71788d827062af4e2345c25692bec39c12644597eff575ffaa2e8ca0637895d48bffc7c84ad5d1005cf674ed22267d7de63e996ce04222;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he356ff3cf7ec6318f515132eda197fe05505959f94380c17b63b76ab98033283124ac0fcaf8418fcb88d68125f28dec415fef16431302bbd2a9bd55e78f975ebd4684cd418dfceb97f9b3e1ff777c311fd7d85ee8ab44ec94b15d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b234643cabeda348f7f5fd14583f14292590fe6e286350bf21252e8e6b3bdc6878268eb59f443d1d0e976a1e3e6cea1e63d1796a2c5319c05a0d86505ab07def8919a436f4fe5060545889365659655d7e1deb6ea98e552529134;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb155ed5e4a3090ce34ac98f838f9ca9c964caff356de10f9722d49a3518110ad9b03cd7330e9c8333d31ec46719a67c3a4f3dcfa028907654fdc849c9b4bea7f10f1e7ae174db514491a6a8359ce0a07fcf59fea8d0443efd83dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ea3ca96ac421e5f520a2f18feff1909cbd450d834e61e8fe2105a6f53ff1c2cb168329bff605354a733149388246bfc9914f801a66acf7da5faf73dcf799977c5eef64ae117727f53d4989673657d5c2d4eee18b8afa5cf988702;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fd34d259284c67a45c353af33169e83849c59e08d84df130c9c073222637ec0a5d466db93b06fdd48af5d296782ef26b408b818cfc1e2ea28098f94e5a16a54c56a17b43e1f5a796f1e60846b5568c17da763bb72f00b5babf9f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2716287aa42468d0bf771c9e6333c2be7c3e9a5fb94831c179382c9a39355d1e9005cfe0c1b006c434c157fb8d74d35d4961c73e40f7dcd85bd8c5dedce7e9d1126a7d6ba3931ae14c843e6fac442189fc5e7436b1695f261f1791;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7ca9be64b0cb6122076dcd211a27a41c90c1bdcafc68732e666b5c79a3992711cf37ad083801f06903280716680df6ac539514282c9e31d844c08d76bf59a4e4419907d12f34ae2342bf4428060f1b4e31a0434cece35c717cd4f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af87a0403c9f23ec9c0dd174dd7f96c6a8636fd4b987383e923818b6ac0633e70b2cf2051e0bfc9c64c41b951b123d2dc6b320833bce65bd103fd4fc6a381a3d433ffbb38c58db34def73bf77ca1d9d1d7e6a3bb3ebcfa1e60ea3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33123e8cf7ec71f69b9aa994d4cc9eac2a9154e969824dbf3f5f652607e779a7fd1af2246824c73d87399ab85fdff95d3c7fd5cb3f546e00662b3a62bbff74662b4ca3baaa825e2c4ad4f9c9db210ec5e1d91b7936006701cd2b39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8508aa09766764a93d502789d3b356f4274f12ed2ff19e4aa47df7fe59d04dec0164c719d2cdd973e873a3e5a4a0cec192a0b7efecbfc59e7cd7d0cd74c401feb51f847b8b904cf772efe483bffaf1dbf82e05ac4b9a7f2ce1112;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1842be959274d54d9661f604af20d694467793337cd0a2d1ae73c1b9d882aa3869e630772d090cb53b77f71cd7754e5f5e9d6cce5354a806cb4bfe05b6dd574db66197f6e58f6b9bf072b7688808da636e50cf9164fe357670905d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be9f84a0aa4062ad5e74e46655baed54b564b83fca6ab763060174f6045aa142fcc617817ddd3842540ffd58e02f5f5089eacb9c1b63d9584e3ee253cbe2a4b56faa8c987f260aeaafe99861f28509ceecb3ad0030c76021a68f96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdd48becc7c4d514c3e3dceb6db6ce0cb4cf0ebfa5507a37183a32d1a1c3cff9d2172db1c7981bd33f9e4acb6fa446730697a1a63cee325e687b3e32e3bd91d8d2f4a360ed9412c14af28670e24351242664d5dc1a374a83094d62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd99a0f925ce46ad0a0792599f887e305f6bd59eb65a45f0a1e0ff9bc25530b51881cbcf7ed4b56bab4987e9819f694c9266f0f0c37ca36bdaf49de8b47398858e3f525dfc0e4d4186287ec4f4694800ac767051cc27e3d972bb04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a054721dcc5883f6d774ad4667828824041c703d2e86732e4f6208f4051957d4c77de37a2a1e68a30af1224370cd871257aac6b20749772b8e057fd7a2e11fde8d5df065ea7e8a214d2bb22525de40c9795e3a7269131d60f54643;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdd2e5893c819ff7a04216e7313bd9c9dc65a631b014cea036f5d82cfc2b04e5e3b8957af56597e4492af02520070309ed9424dcc455d1d7e029cca5643780de0c4ad235fcb44e258b1835e8261157905ea65b44ccbb31a99eebb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h615b7a8872812c9e8fc3ec462dcfd8586efd7632af96a089d1281e61388916b52234fb4ea5b72a900678d143838a94edf24406abab590af812f61b94bb86c4da59552850a33cfd45aefb5b2a23e8a1111e1bbc9ef76d28b66a09d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7483d86a035e5722db0bb93ab89f6c04ea3f066094def19ebad4cd259a92f2367f87b73996885d7a05ded9030b8750a902ce8a27627270ad36e886f3a915a0329ae183b381bd0757f8b8608409adf91ab525bd9fe58f05b23e392a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f83a6a57d5c02ec61199dee3b9a04b51733561f4e2bc19b42a37d9449310891c0fcbc86a09c65b46157d5fb83b5a147e83f75865c780961b674435e1fbb07df2ee57bcfe783f5ae0405435d5e5c12326ed85b5f208950ad07f77e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc2b33c4c3807e43f409d963fc0aa4d6154e00bdc5b69eb296588441cd61c5b85e59f2152e78d28803f49eddac52f24d4f14a08d25d6f40352b963a5c725ad9f0fcfbd82d8109e9d458b47c68a447911ced11604314ab23e08338a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43566fafa048364f9875ba935f9d9a234e5b4b0f625ec4ca966a245fa9acfc03639978656ff7b8a700e72182c0a6e17b5d00bcd989f3c6c057d0c00d404098a3171450c40f90ebdd92a23aa33387ee1718d6ee50a69606667ced68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3376a914970ef21f605a66b2081fd70d2afa713d84dab142558f851954538ca0841cad540e51fc171dbc05a23cbd554426f583c18ea246fa178e14eafa2afa13af4ddbf82b1858d5a14d832409f29cd4605b03f03ef5f201a763bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ee5ab4eae8267cc9bf762a30961e1be4e1173451667453f8e86dafa5ded8f6965e5a2c1e4ae78268a50b5d10c7f7a0286534b8ef8d882a23b922363e07debb55df2c0c324df8fa6d8dff51af8150a758839f65adf0a639244040;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d27d9bc989a1b7707f6c90a0ebd47d8eb7a949c010dcbdf9396aa97042df1c6b59b377e81042299fbd0e48103dfff20fcb0f635cd67fa5cdb735c9a1ed0e7c242f546a3030b2988bbc8d87e72a6104862df7f1c55171017d3dd58;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1085a19b5a165d5776ead98a74e406a14b6066b40e1f58d2b276f9d38c6f31f8d16ae97d081b37d2485ff2593c055f64734bc084478a2a13f1f228c5e8dc3d6d3ef7ec4bd4cf9c515ad434abfb1d11b74dc1714ef31966c99a76b9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84c1687b334fefda05a9aa15d66b86b2ce909416b91c66e3896cc6eea7f0cb915847b752e0cdbd5fdfe2ecb87f3637830bc6be126c1df93dd5f1dabaae86b8f7f2743866ec99d180cf9b26b26611e4636e13ed77f8f4e0d618fbb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14379c77616f7583c4761640526aec9d729e753403f205d4a98565ebec04627d68233febe18df47aa0308b9346f8b50aa53d1032c43910d173615b8b62120903fbcda0bf2c339e80447d092ed99645bc8bfa273c906260786d732c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b8a5c1864a4f43ac3e679a49afbd6c88742d922bf0a6b50c77cccbbbe6cddc3b154d1e487170023e9027e41cbd2eb3d0d1287dc0498d7fa3a7fc133cac4c0396726285123cc3b7b2b5ffa61d34cf22bd4fc4b63738cd3d4d6b0c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d47f73724f680781c05ca2580c44e41ba761db4f2327a135fd1a81aa64b71db78391917829e51e6bcfca4e884c10f3beb216822ea137282b9d33f296660fa436ae6fe6053257d72094e194d4e262b0831b8b2768dd0ed9de08bed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4edb3ba738fc51ff91539e5cef3a6c964960a24e487f31441ceb634799b0f0e20606ba68da745cb64e130344cca19b5af16ff0f8f7bf1c3e0b71d464a5ee18fed449c546f62b5abfb176be581515d09c2eb65da6e9802f2216bd87;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5fbd75f6d0d19c8130bc161c3e18931b1e7376de6163ed7be2617184d7fffb7247887d6fe1f5daa789912bb1dad6ad717d62feaa21cf6fabe89e31dcbd0f4e92788e2b046d51176f053f12033a9fe7b51ada75e1e5b0fb1d8e441d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h120d4e1da4e6403614f007bb5456f08e62ab32e4d23f0e2709cdbaa1ad6f3062a0fecd7cd9ddf2da1e075e328bdd37ed9bdf0454a8f39536c0d76a17733cf482aee2e32ff027078202559eee23283cdf7487e6fb62d83d71e7d6cba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168e403fee77b3cee4b543b6c9a6db43920b188962f867db2390e8226e6408b4ee5fb00794b7d93b0241984ec1a5197ae17f19a844bcf25e5776b9d5f54143894eb147ad49e5eee12bf29d3cbf62eb85bf6a3bc7e007149318045f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1545bbfc16b3a778eaf16ff69f37bd7ef954af7af50298471ac6e097d30f03ac3cef1735a81c63a683f20849d923dee91d5daae9c786d1e135557bfec71c3656b9bf1daae93105579cd4fc68aeddbb98f486a629d4a7b39bad0802e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2b4b1ad97eb5f5bb36b498f323458db4e40065f91d7e7aa07356590e81bdec181c6881b091c3f1060d1861635e12d1ec418b502e81b52652dc400588c9ad4a130619cd8ef7880d59c28ddc91526037b958504269b2d8023d994a1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1906b31fd2b29d973a2d3771268df43888b4dc5ddb4df2ae89a85ec147bb9feb636f632048c837bd241d4064f18640bd18ddc08d7c3715dd63bf7b4394fe2ee2fb3f5405ea5f21217d91bcd82bfa1ec38f7ae672e1ea73ab87c3431;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7723e1dd27c7ea22468dcf080592378b85784419adc1fd990929333e7ad6f4471b1817d83269b71eacfdc91555d8e06033eec361d0439b657268cb00654ebfb26cca551d82083c1cbd62fe66b0262a6dd6e12f4f097c4eae6a04ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abfeb7e06ae9204115e88b687f9e9eee4a399286387701bb3c927863df913552ffa1804c03b11782c50fd56d2a4a169aa38d7a9d34b3a21f37b2a017eb57d5e1ce3c948655985cd1d27f43d35f7f6d3caf80b08bfaaf6fe2515182;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a25b3fc4c30cf653f52f2b16b11490f041b7de9f23a91e36d00cc84c994c1015e3d298fdca87913ebbbd5b1e75e69d0fb8091736741fb9221fcd54e2ef0157586688f87b2f8baa8bee4537b1baf6d5554a9c5e25133f34d637a77e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162f8d5bf86f88bcff36a33056ce0b5cf4aeaca2f4eb81e41a9bc3c42d8a5adf2ff7374e54115f98e9a5199b3ee7fb4e91a0a04b28bbd52ad63cfd8e16c79d89ab27ca0904ed1fe6dd20f74c7f9f980e2aa6732144d23618464506c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea33ebaa03f97dfebf8be707be3a25f703decdb3779d2ed41467d24314778ac538ebc13495474dfacdfc645281164feef2346e92ae4b3864aed74864ad4c2b71f8f1984e0606df5691a1bac164c6bd82bfb5281e3d52c945cd0854;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a53e5766dd57589c6ab13ab1d721d52ca93e45f1bc23b1d7cdd1df6d8ce1b2f8589f0e3a1250cd75efa3354db67107cc37169abd6e14994e4970801b48ada65b911d1ad0921d24503b0bd705ef47d86e88008e65445cb709e4eeb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha23fd232023b8906ac36999457feb14b46d2c3ba7190dfdc6c5dcc50b095c1e47daba6ae094ac8e2dc9ca78221f3f506710d57f25ea9a4dc77eeef7752941980270561ec542cec0a62d93ede7058b9554ff863c9518f44ab56f7c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec37bc490a5caef1a5feb9c805efaa86641709b485e2f8502aa2e217a0644f8f438f5d621a087b0ed9589f67116dadb45e69658e310edb7d8d13a9d348d1cbfc75f5eb79279cd687408b67e94c80649ceeb080e0f855390fd8e398;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c7731f10646db9c704481a77cfdca75ae4d1a42eabb5e2da3cee774898e303f7ecd11e540b19f863b02386600d0c3ff9a3cf692ac7ff19b8d4019b8d5cc892326834bf91969d9282ee76c03ba793c8dfb2ac2c851a0d3482bba68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1389f5ba88aee396018b3240eab9d9a6f420aee0af403b19be2e53780af9f7c24c88a7b90ca47eaa953c2eef2ab16084b02e2dd227da68deff5939d49c6103e42928c679e1617579e17463ba2ab36a757df040bd07db0dddfc9027;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b9ea0e0ce9cad374cc76d0cc3aec1175d69bdb98d0fe3c8b709ac894f272f500bb1d63a5a2096ab06a0f39cba625bf876f0b1495654770251b3b02f790470375ad1b26b263be3214e549d9cd3faa5e08db327194c0163d816f226;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119939e0a675adea3a9af68d3fa7d4c02828088b3e6569a6194c942139caedac6f8399695966ce1c269ab10697d0556507e0817a5bd1598e6fda7878919dcdfbf5df31ca347a351c07a9dfb7396912f8d8a104fc0dee5273566afff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h120ab70a7c8ab8076b04796282e11f99a807d8b290096aff51be993273d403a5580f648b198c42cad3d53f07658fa58fa25923a4cb225af57edb16f25e21e99a1e043f17681c75bb2c8539fd9de7e4954b0e437cf7b4c0a93ef2b62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f2dcfe44bffe7072521fe7d58ad87d576abfa7a546eb28f7540f74fa63afa21f65825dca20593d8574b634bc7476b3a75ac6dee2c1c61dda9cf801ec108576e5fe2db79f3c8ff0841ba60d71d10b3497c033dae96eb4efb490662;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefc6b9ccee00b5e43e7100dbac5bd89cb28021ed7a9ced11a2933238eb318e8dc1b5eebb71501872b30e734afe72fa1006f8f6ad3f3d10a2db80ba3357690e3f6ec7c80ff8e78326da9664c2232810f2aa57a858df34a9155edd05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7acaac20304b9858f47f78194314d77a9ee3df35599528b192a7c6d37a9b891b3416b9230d0b7a03719299d111db31473c5aa72178df07083b3379e19fd860d528ae8dbdfca7df32a2e7061fad1e9f500cbac51e1b5a37d13c5d07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad5130ba4f74ed005d21139000442f759c1ea29175f5cf9d5710a3cd1087e0681a3e9822afdb3c24d17d40dd131ed03ac1e2d92381575f25f7c11726aec96c41b8e0dd579f3df92e38f71f04ea28c4b3044d74a91a4447857ccdd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152236c3229d0ed347d87351356769f7beaac862d5cffa48a467845efdfc9899992c67239816d867d0a129fcf45f7b47463e15856572aefb9ef9241bc57174693a8bd812bd2406fb8826a4214a783bd8a1146546917e0941e3315c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180be32bb1d91f8de1d8ee2eeca42e4198c45652b49829a5ee53a0cba4e907812e15d41b45314a6db779f0570ff170fa660511f9c82dfd2a38a1e6faa951b329c66093577380a93ec11676a1707772f8561b47d5db70b66634ae452;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4283e5d8112f039ac4c8dd4862097ffd03d7ea8962be0e82c753a516f5847ed1488ad23b7e44409250da8c612cf03ba94538aae6d44c791a78ab7b012923734608388d74399b3cf111a27c2794abdaac1b9ba1cb05c344281be061;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c3504037f12e8e847d682a81d7106d87948e1e95aeadcf14461a1fed514f5926a63d8690fbcb7668b519a6d40b6e7f8425fe1b9f740c000f57e3fa5f4afc0c4b08298634a89f97ab81e0b21134915ebda78c2cb30df126c3ebd20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h363369d9013b56c5a9eddb50f901efc4212074b1cbe3c7fcfbd4b30bd656fbd950807fa924dd7e775bdfdad75d9c96cfb4107bbc6c639fae0764383c431f7bbc39932b625d4e5842586a11f43e6cb04267a9d4ad2bd2b04a7bbafb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf915b896dd38eacb7ae11eefe7a04f7364d824a0a3df788dada2a1296619f46c52c41389776bdc9bfbe59fb3817929f502de37420540d18c7dc52e02ef38b66c46d5d6befdce7df0b46ddc843ed0f6862befe6a3d800df0854bfdc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1025b3a3a03d76678014aa04cd08587bf0aa7572381244f487c7ebd09994e5e730555d7b3908eba99b228f2e8267289fa839522776f1e243562079632c6806a74b3a7a819c9b526f3eda5a43df09bb69ae364d053af41ccaccc1cbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146adf473197f37c5d1e12d99da1857e4f9eeb91e6d4c64b06192f76ba3cb8d20566b271b9c54554aee7741006cfb39665498c00744895650afdf5bc2feca50ba8883878efd23db2c56560dc364b7a5a4aac9218fc51bd3e1c2a729;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b2f60b95d88e134f1a6a6b9c9c0b43586e3116bc2f5840d52af5e3ffc578a11a97e887b79a8bb65c7d95eba8df533e320c2f7364b1ca6bc41d238a675653b0224c230d08e9504457a706a95603b7b44c486da553d2cf5667b1e4f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4b8b095863c06418c8f3bbc883589e98e59b38f0ad52cb499825cfc347fc9be8ea1e7a5598c122b0a01b4fec6d23e1a724184f82ccc34c3d87e4c1397c2e408af4e1dba273e307556eb1d8f88eeb8779a1f0b50ee2df8b12e9773;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6cd73c35bde110b0f903351f533964beb8f1ce76d7df9c95142f5e07c01751aa787191d20304a55d9f5be7c77c4ce4e604dcff1fdc6cdd5cfa962614266f7735d6274ce67a716c48b2d297488a4ab0430f530df55c885674f6fa0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b277133040d38fa630b0b1a3246cd4f2b329388fcffac4cde0da6df5c3ee8d0b596956c7ea3a83384186a2f1be1db00ee90fe0d2abccd5a3970a1eaa5191f675d6878bf78a715b2e1d624129735e4a7b8160ba2c24e317fd25485d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'habf5b0ac48e06cb8ea7961a33826d405370cb13ef02342ffa6a54ed16af90d5c7043bf33475afe342c4f378f2b3c2ed1c05532edbf1bb4eeda8d933525d642f6d131f9f17300f7e105110589ff633a0ca3c8afd61d324ac54ad257;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184422946a5724a3f0cef9d3e525ae5448dab76130e727114311d1d830ed1befa1926189df28873ca4af545f66456cc624a2dd30015ad978d0ca9e5639ed466aa004fe898d5541d395327f0ebd9ab1caf536857984269e05e008e38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115f20ca0394c0787486d1fa4083930524e9f74d62c6933ff5ec42bd62c166774430a0654fd33cf5fe7e771ee395e80a52eaf1cf47ef9bad7cd2709435353f2c1d13d17250ff0989c280d4f1608f0ea71950cafe9105b37dfe6519d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70c769c46258bc165045394aa8e7c4044eb67ddab80be2ac7ee771608061239c7bb5e1087d5bea768031abf6783dcce01226ea0f47cd687975fb894ca1d6561872d0db14a1e2f224c69d8b42075e9b884e08726594907f872a7d13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h209ced4f6f748d8a42d671862e6b3ec1a52b01c887586bf96c733a29904f046d2b8a64ef1e5194b8d2e6541009812398c2a03dbdda6b6456470d938be78f07d191467e9ccd2bc09f91de506261c8eed1536317bbb285ab8d4ce3a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6d50f613cc6404d11dd028ba6155826f5600f8a81efd1bd67c557be02cf9fe0d037778485001841b3cfdff18571e1cb42fbd97d55d3d41b467308a1c46651f6d30289d7bedfc6c4f23e9259f02cafc05c3f72709f8f14be5a14fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdc1f27f1f2ddd78d479115f0697253530668abb58226b5101cd2b285240ff372630c25633b3fc8400fcdd3b49c50c2fbe95a0c2bf6181210112e0dfe2ea8d03af6c084c630c913e2ecbb7f54b94a771ac95905788ed9ad1d6491;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116ed1ad9660c1585fbac96cebef4533c24a149defc74c720276b93cccbfe06252506f9e4ebeca918f5a859a03384aa1d05df37d52eea6d5fd325ac77990201030f2b1c27700144865e9698a781ba0e14f52e60a3acb3634f888554;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19428d37b3ff005ae4b6eff7298c79d1a988ac49e27c6103ee1dd2de824552b8dc2f86c671d73f2f51dbfa955daf65489595d46629a0c2e94f08d75cf7a6a00aedc862b37d8f2e4fa2650871ed9f68b99c2ee49fa837a3657ea7235;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17da3d689148ef6e3adfc30c075eaf47abefafdb06c09e52320fbd15d089624884a29f50fde00fdf50475cd3b5dac5757d2057a662a450a90beaee920171d116968bedad996bd626e712e4e6dd77d72d8aceb9dc565129064826589;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecc7a74e4c6a02b73ac43273bee2c27b8a2374e06a0ed35690d1fa6166da75782ef8bddb5c3250be9212e0b49b3775091d5cd17ee446d327c39e9f26139c1b3f9e90797110c2193edca7ec0f9a55b9360ef2de1b59bc97bdd297e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c8c6ca3ae0726358eb805b34a402f03df54cd1e6d8ee8fe8e64e6611022ae20da6cfca5890cebed3ebf0da28ae7ffbde18ed9e850fccf9b0f71b7fed1679e3b7dc9a78f00d83d9e3f99a078458e674966a6399848547a3831705a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14deee30bbb55d2a308f17cd99bdc5bea9ae747e28a931e770b58c84bf4624eb22778e77fd1216929233536654c83abaef2fa0e88cfc3522e6611857892479aec5c578ecaf0b3fe7fe30357552455e70f1346c526a4eb38d2f8c2f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105be3efc4dca80e05feff8699702e66502cf85b3fff535ee6f6842008cb3ac45debb3a4b0ee7b5f8f87ee04476b0700c11c7211b8e1520341e4182fb932d846ad463e2d71e07242788934f61d1273575decd26ba3e07083d2665c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e707cf7975702f0d5f216ace7dba502bcf826a4a58b26128db9c736e8ab56da3267467a541fdc02a9e67e25068265fcebb09d67d21062b5a9e9e1721e04226abcc4fffd402bc40e3f540759d46b33db343eee4d425ff4a237fac36;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11380c6d70981ab728102875ddfd70deca8bcaf3a3b6b5f9c31e23e4f42a4e4b90244515924d8afa0ad7821de86e122375c448de4fc0e34c09295cd070cc43f21dde63701b3e76d271f65a5f06575d0521ecfa6c848e8754aaacd05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha31d8a5288b8630596c56f9a13af38ac10a7a60474b15462b6a350858b606690f593bec00ca9b32870e66208c785c677ee7f83e33b5a16ff59cab6f98bd8e7c35ec2ed758ff657acc428040f2d7c6a6261b8d06c5ed71553c2b240;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8bfb52a52974f36f4a44439090b4aef0d3ad79e2c70e21e3abd25f5cbc2224e6fbc01768f88baff105dc6ab6666944c8e5db02e08644cfb1fb83d3a6497e86193b0b95d80524c5939ae9509f80b39faf1496a286a69bf0cab6796;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136c101c989f1fb74a18bec03c6fcbc6517df3547669e33f4fd3a5169af32010a5fe9cee69123b64ee3fdccdfcfd55423a66b6588860c4f8d2394a3626c561fcfa5bb2251ee1f0d59b833bfca335183aee370935b05a889b8b3f487;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2c86f416acb60f01b6851db20781c79ea99564beba862daba685046e9cad37d3f6bc9d26fc38c7f6fc9146ad5683fb3f223c1ab44cb71acb4a6b8549f20eb5533d148ea0c9c91713038637e783b34eec640312942e4ffa909e989;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1963e47f36a955739a5c15f7aab517b81225ca4f0643b0d3011904d67100a0dc19a50f10a8736d3a75ab7250fbd67be0fa0b9ed11239bc8202aacc97b6473c0f3b8e58c3bb839c40f1dc560d9d8ccdb81df242b50aaf69b0e308da0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heab032bfe177aa4b38a83888a26d3ddda91bd7509efb43aac17268479108f1d925b2899622a18b0664dfe238e09dce7e36f215c90321eca51943fd144acf04461da25177522b76429069195d8d3597db08bf3a496367ab745c676e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb86c138dabd78f327e377a078f36e2ab32ed43cf0f93f1005506ff94f61dcac11063978d958b2f026063035d9b456afa069bbe42813dd04f16a62707201fd26eb45d8bc7f60388aa33d611e2d478a85acc96ce5c2025de516af9f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b033ca43b1e89bceb9faacaeba2432e3512d0fda72c466e530610b3024c080f7691c26710efe9c97f27553aa5d8b9b3c593bc9ae32c648a1a22a9e545c9d87059d8e080f25a67cc8064bfc1fad41556836f5c96db2c53a18e7915;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b676628f35d4e158850d90c2babdfb7dbcab59f83c15940e8b747d754f0de9813b354f2566b7de2f46a970dc77a871c8819a4528276b72b7dfe51f07013822f801a5ca2bb476a00ac446dbada49b8b784eb8e5de940a04c354ebf7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc4bc1529a71e8cbadb2bff1a316a0a0504a65ba7179fcaba5cbdae6ba7595eebb96cb683545f10ff2a55cfab03b716fd2550aa8c12d63bc2cedeb217f9119ca5d7aff3e66ba126a7b6e1f291065ce34c4ac2580f22a1febb78d2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb779e41da7cd5491bb0ad45c3f53b2c20153928853ce0e04af614add8e260623ac500996c7768a49ed9b02461d63fbdc08a7a4d7a3dfa192c2cf41008c1481effc57e27812fb46284b73fd193b5f6a716ec43abcad25134e30d1b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa97b640967b3be97aadd157eb8ccf410e8c189f53da505817fd12869930887a8de878455215dfe75f244da2298da26dc4cfbd01eabe17b13b2159dce3c1f07acece5bd152fc978ba2cc5d02123df7f845782b4cadd21a5ae28538;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d553604beeb2f657c793c3cf446335c85fb68d64cd0cde2d17e683c28834623dd9304a8449c627831a3c8beca8c4e0a18f218ad174435c9d7528874893bd84370a426091b7336b3ce980fc9bdfe029faa357742c9e869fbbb9a39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb805313289055e54fb2f3ec1b1857cc134c3f976d1b35765e60dd4194c2846729f48ac8a1186715df1910e4ebef33d5dd585177f6a7881720d8647974fafc1721fa3322c99ece101cd3ecec979908677efbb3b9b761ea8b385071;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abd55ac50bc9103c4bf58b9cb84477598bc860bc230693f0b9e331241ab371f713c11cd37c3209a3fd7b2ea0fd5e5ba5757f3cd2dc860bd6d5cc842b73a8074f28f38af1e972276cc9a0b93ff92787154ca3ce7896e722046e83ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135c91c1eb295bc684592a779d4044925e416b3a1efe743019a0a939611664e9c1ca0a257963ef65e72fe8ced0a338535cc29b1bfb15497d1d1e6dc26e7f4cc34d48ba645f9d8565e03164f9b212c549d6fbd41959dc2b883a037a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h730de77f29b248c4814f01add9669fd2ac6413764b6a16c5f00bf0e81ebd4f2d8f31bf11ef970318dcbcdb587d76d9cd4765d7af81ac7c5d25cbb3aa9e322cb7dbf3bce9e7a190a77874aef1838e555e7da6987dc439870f6cf3ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158a8c0e7016168cbb2dc3be52458f7ebded135f021002f639de7d62262ef463c8bc327bab007945ebff0418bea92465c96391abaccd6983ef8bef17415a25f81af83e2f003913d55fe2ddcecd54606a63dab5ba6aac392aa0ef0c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105f0b7ba1e4c73d08c6fcca9ed770c83bc2cc1c419fd132df3c8780dee513c8fa161d95b5e0bdb2a7386d4d1dc0859cf299e771038bb87d2d592fba474b134043714913eb4fe600a16764fc6f94fae4197132427e67e96e523b0a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1d73c2632b34cba21eb7bd4571d62e316e963727211daecea9fec59b93384496dc00f4ecc3cf5a631608a482df5b0818e5c563de131e561eebb14d5b2b0f0884411dcc63d04085520a2243e6c1e11aa5ef06213068cd65dac7b86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af16ae1df9b0b4767bd011671f0dc5ed9e48a95c6cc716a283162a6a795770b25d3ca9dee95f1b8e6a635a8174707805ebc969bc6994891ca430714d601505da31b008da93a04f8fc969e233c20d4382808dbb126e8da65fc6ff3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b10aeaee0c932fbd6008fba9b97549aaeaa702ad7f58737776f235fcc455e62a558e5be6b7a28ea9d859291e97f7fe3a42cd898814e199386a5aa49f8b0a5e59d69126bc009065f8ee131a9c0bc35bf64fb0535f8c6ef6c0dbf10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h393ad437484affb6f2d587afd3dcc88a2d1ade88626c6ac65226b10499bfaae316d040ccfd3d5f3099a3d3fc6c81d30ed766f988ef4a6e2c6de050ee478f5805b8568d1ec37e744ba8c37ffdb14b0e8c0bbbd03ea4531824f87b93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67007f57ddd1333ca08d31061f961cfd2af763d919f462ceba3b79a8836ae9105e2517a6fd91306fb7e2af95fb7a25c1c6a799fd70e1f5b756fa414246cdce75398400828445d0df1a2da3b8931e3e54344a9349ebed94bb896cff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148a9bea229cd2504bd6b6146a10d6c83d0b7553889810f209f8f4c6504e22ad8c0954bd349ea3e9d82240699476db14b3a8be3f71d67dcf8c184fa0002be076c494436a6c8249977f2b85995e5cde4236d7993f0f9984857d588b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1718fc17e290f5fbef8cd1ed8fa2dc3c7388a0f0d9b98b4304129b49dead300c12e5910229003352f5efb43c3f9d6ed589ebb45989099d8f8bc147cd5478d9f4ccf41b6c7cab6cd368429d97b66a65dc2cd09e94b603125162a8724;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f0a199730eaecc02455d940a42978a0d340f1e82c648a419c63f93a65b4a93e8ad8719e873224c47ef0c243de24e585b8314d0677ae4c6445223469c84964c6afc497e0fbc440b1cc0defa73564fbd8e5acbcc2a3f9917719c40c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb551f13a68a70c995092b59628cad93df266ea7ecbdbc53185b711566542bd217c6f740752e687e6188450cbfd03c5ee277b76048be44fd9b5fe74490b1407b490788c5e63642d370b571d4295325adff9b706dd7f756a95357f7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd89e11ff52f2e3af49568c0a9d1f1da60de8805081f073dfb903fce034d06bdbba34005ae691df3ec76c71b3982d662182850c47e444a961f8240ff51c2763f2199494fc1acf5a00fd2788a120a5978f5717bb00c4b07eb855a84e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16972602f00a02bab9078626761d53aafc95d85664175b1cb47e957c81928728d88f371ecffc90a8690e010f45b1ff1f944c9dafc79621c6710c3a09f84051253085a48de728a46f096a3019b3dd5bed5eb913a92452775dc2e16d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94e40c3998145773c666c7516f20ea266465b14036568ee931c1c215e88957db74a22b492afbf44959b9985c80b21c66b6d1161c8b3a02253422d9ef74ec6ad513bd64a2d31b463eec1f25eca368c52024b45d5adfeaf55fd6c255;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101dda1a16d1be726a3b1d0bd74e961eff1e2e27403d2c146611024075ece34c76e1d4e2aaca61c65877605065cd3b45d02950337a79300356602338cce67ce6a53d3a7c988f628aaebecbc5ebdb115b5918e3632418750a241b13c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf554b9b9de071a35362d461a020578006273453477ef31cbb7d5194523530e63e836a795cfa70f78012b0b980a5eb3c808e8e327b12b7bf7516d36fea1233cf9ec37ef3657f9cd78321fdd2ad2e0fa4dfd1e43550b1acdbf6604;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0eabef96e3df18f32825a6033e1813a9ff85171ad3adfe56c014fd597844b097509ada76139a7371ac94b21de2048a2cbd9d4f1793478221223d2523b3b9371aff0854ada7f197b7e93c385b57e30669b2662e2733e53d17bba14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59a7209a54e64dffdfaf58a3f9a2bcb02b3b77fa57e1518b451b8ead094ad49962c2f5482b70e7377a55e45e6afe5e05025cb644f80a7c6abb3923b6666d07777b6d643e8a884392fa41158cdb4594289c8710730ee25e629b1a8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd07b32d198451a0bfa113a44e36161170d305439be370d4b36e01152206a3c22d270ab3833319673d713c944f404e0d078f337a7bd46dbdd49f0a47ece712994f6a90bb0687c7c3c404f4875be7195a1744c97b37bf4014cba25f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1399ee46d24dfef154c50c540a78681a61d030e4833a733c5da4f59a55839e94e9508b8cf3f6465eb897fb2ab633edcc446004c420513e16404d1898f27bae1db180e8ee22142b95feb601dc3300d273b937a5d68c84c8528de16e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76cc72402e5d4a7d1587eab29483cc09329342c6fb5c0ca8ce7dac78fdeae503724278182d5b5404e54fcbbaf46347bbe0bb34faec616e57a02f7fbadb8ba4547f039cf763d2a983b0811e2d0ffa92b75aafaa66545f355f5c7ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59885b838a242f4876c7e5761397899253c19a01c4aab912b67fb6857785f33177d71eed126d92feee38d636b8ffaeaecb0d4b21f0a82c6284fb71d3bbcc6b859cb378b6b5cb47d6eff484a74af467764462afbee17e01c25495ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144f42b73428aa52349afd8c0b2758c4678c4a3b2c4afedfaca02a6f122a944024080f106b75f57a3347e128d02e871d2774f617b63a0cccfa451dd68ca2e92911a7bc1c7a9ec1d90e0803e91aa779f16d73f2607a168692c477b51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164f02d0aa0b4827bb51d199d9a05285a3110027f6b9c0a1c2e40723800f4f0e377cc5d112f267219494b016c309db2c1608f38f47ae9eb07346afa5d415bd3e4c48ec7a16fca17169683cca6aecb09de63afb50f09bcba0ee69fc2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13693c216ba5070b35fb40b5ec13f66ed62e0be94039be75cb0537cb43dfd3f87c0f90df79e679eaacc94e78b566beb8c7ffcaa37be0237d1b8c6ae6614b424159ea27288f31efca30c2256b47ded8627db202be10b02ad644daa6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14df54637546085b4ab0dfa52d91441e212a2c05488782078a879993e5625e16b0771e903d5ce6785824f31850651e3b26f8d7cbcf4f90b7c45e8d1c37b7b09f074971ff6c418073e4ea1e85787ee1974e30c3fc20c7112789c17bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1894c524b8649c0f2cee4f55762eca2d6c9c815415cd696d63f7aa158979fffbc994ab82033beb7daa402c48f655a2a9adb8ec81edee03b4048b28f9b714de3cc02f17c114e605342693eacbe5b875684b76eec5af92e475e0c1a50;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122723ca0dbb0cdb42607e452b2a1a071d926edbb285f2d3f32d068cd8a2792e26a40b6c724128b77e0305957f0499e32c7eb5858e29c1bfe5b585d35ff1ac34129bdf0dbd1eb539b34872d644bfd1f0135d27868c2ea0a127c2bb1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc68bdcd28f20cc6992874037b0573f7da0a30eb742d0b575a740f4144511e088b20d0af7614e174c309feee4c06443d8cda1607158d95a392c2f2b9adf89bb18e7a32c6c25dc0f9667037c9375fea26c18fa610e2e79107683e35d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fee86ea0554d890787c6ab3b436f823874dc6b4312bdcd46512454ddda501349ecc328a0e8bc54a866b42882745cbd7416b5ab3385e6b2e658522a6e4cd50bd75bba3869af1bab2c50eb9dcaac8628c3dbf82f8e2fa9286e2a87b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7126b2ea194c1234b073535952e0b657392c5e8b9a34dfaa8a6209275d994001de8956a393db6de2dcb7bd9a3e3e2aebbb8c236e90a27c512eb30243750aae00983aa9deda8cd47eed4ef059ee67b1f033164b03f616214eace28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179798ed1e13ce8d3d23f959bac4b809d9899cb358f571c8f800a243e72ab23fcff97a540e12ac43ff349f4a5aa07a353f5723669c31bb417fd346c0eabb128b84615881b8fc6deaa27747044161fe67e69fe2d3de943412ed370ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9d7ecf3211587c97a86710fd0df0027de50947eef53615d5b8009302b02efdf71544e4096aee777bdced74ca884e830919808f54d4078d870ee279b62a997eb2929533fd40e5501dffc48dd167ac2b5d5cb223e77c82a261cc812;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h200111df33f93019643ea0b54b89d1dffe8ddb9e4c3288ec07b0784f7709a9f17ef734a86a9fef5a4726bce13e9f20bca5701ea5e0927e764e432bfe65f6462fecd6ff6a7da30bf4570b7e7856950100a5fe159b86a5ec34410049;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1319e6541c0e596b1ac32f9ecad7bd376af174146b93df30a8b30ce11d9751d27a79f19b92c894029d55f6f48a9f2fede2537a0e9519b06f76cb828d80126cdbd289bcc4d9b083cd21b43e276e72a360e8e26b58e3154bd24f86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h474ea9c47a7d980030bebcc75b6007664f0bcb86c2de9092b410665b9cfddb9d200ed3b595d8f60ba29e76d4c9874ee026e8821c7437f3f2800b9c41c6ccb6692be46a7017559012e9cd542c2559b7de9dc57851c8d251ba1d4062;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92f537158c987bf9baaa6c245b39e33172db8639fe15bdd363fe9eddfca4b3b10b3fd917182cbd431f5b9887f839666b763c86824d8e509e4c071db391a10cf59a4aa5eb611d76d41463da08870981eb14cd13825c2b655c3153e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d0804b85bbca8aad8ff7ec942e709e9810b25812b5a7fb726ce167749758f3df40d153094a9e278be5e188dd7243a6d75052505f45bfb203f2c470cc5c057eaae0500857af3432999a50efae9ec0db8cd823a25b03de092cbe69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d93465e6793311ebc94863a12ec8ff63a9c00d447f17ee4e911b3b156a1440e1c281b2513fd86a75ec12d1316e0d2ceb623354c99f954496c7bd178916a6cadc8fddb67efc7b9af9550c82df98753abc8b4d01533cabc723085d37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccce2ad73e53958dcb79de95d0a2f7fdd1ea82825413ea6e53c767174b2c0b07a32a5c1b28846b2f74041e9168353bd6adbc44209a0a5bb2df30928cb11a690f663e15122e2e89b9e87e2c3b91f2294151d4a926e9a10249c9717a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a405fdfb9210d6c6af4d2a011abf9ebf661d2209c704ed162f3728319399190bdaf3a3212ff37be50cd2374adcb0d43a5e345cd382a52083dd1c11042a8b15e0b4833f2f235486ccfd73b67b044b704fef6edaeba427aeb602f518;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7695fef6419235ca8a3dc64ce26a0dd422dc09f7459a3554bac08714bd7a508e643b7a5cddedd341c96cdf936bbbf4ecbb28cc588c502e1d1ec7bd64c119a7bf9b03af54273384370067005f8bffbe371f411d3c21b8d438f1077f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc5aae699cebea1fcf7aa22a35899d99adf0590501a4261c123a8c37ab2c7e0d55a39e8e86b4042115daba104fcbe79e23f234ffc123d8888d675630c80a8e2611e698ba467129786cb76efa90a5d64127dda4aa2ae40c470e8c37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h245c771a7b99abf33fde29f474579a5e6cf7602055d8a8f6fbc580cef9abe3584affd30a13a3e3b1865eccacdb2d807c650078c7f6fa66f561bdaeee1fb8a766d096b0e96c2f2861ac9a95d6da4a9f30003dfdacb23b95f3a31667;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd59f83805ee176f56b9aa99a6a66150cb46f3b9f1d87aeffeab126affdd36e90c83e25e5f54af9e04d3c3644133f03db1c9ff360a61be0647896bd89265e89e2eb3ecd4cdb05818ead07f9c92fc9c53564cdf45bf6aa3a8ed924ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed9cd648eca3bce33b19df62ba48c807b1465ab07552099489b30ece83bdf12ef1649ac9b92df5d0d07ee26016d6d52a07fd14ab50666e0b989a3143faab6d05986168fd78b9e5c64624b389055cc52931371b835fa7d1e33214bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e67459c17ff374d27ee1a1ee08be10ce4332f8a0aa61c44a8e973de0ea5c3bb2f1ddbe61ca5c756b1876cce63b4e13f7c6386efbfb476fe23443ccd2567bfddd576da1f89930dfb8e3e1eb714e4a6932ec5f4eee5e334b258aabf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d4604c0a24fc3e8ceb2fc7627ccce529c56501e2030844d527c45e576d43a62dfdc53e3a15547896f27904f1cf155a28676e22d73d07244c20687ec687ec32b5f69d47da71501ad8dc667052865aec0a84e6d8c3b38721900d09d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112330862d5a7dbacd52f350c1d80c71fe37f65085f35deb5a8a5d9029bbe432ea71a96911355a6c7e80b3039530840f1eb99eba0209d02f3d63d707aaadb1d4a5db2ab2af4859468dc41a0f10ecfbb5672248ec1dac9eb90e43ad0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1677d2a896e43452c39a0286279c8f0ca789fe6f787959abd09e63219f483c35a117703ba69b8a091805d4f841a59fa9cff1dfc950a685095eefb6ab33ee741b7ad6aee31b7d47b35a14c3caf065922bb452b80d0941a87f9d59b61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2082410d63f234656cd717d5bc39b113debfd50b55ce13ecdbee14b427d4b6a17b3d859557a20e3848e8c6e4b277fd1ff44ef86ee82ecfb1a6c0e08a24e1df64f81dba2170c11d2ee95c86a91c01989ed2da7412f1865221227dc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a6cefc8a83924ce593bde1361e44eab0b754feb317e43f7b97a9170969841b6f678b783ad54d7e0be8a75f96735b22cd0b57fcd77435deffbc3a69863731c42905fe5d302aea4d63b913331a94e16653db0f3ab53c3fc8b98fa57;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9a1694284db01abd9e47f3ecf2096190ed276eeb8bc4173010dc5388e0b3647fa2e5026be2865e76f15626413a6b5df7d008147e25bec0a7bcedcf4a7d5dfa78b2025fa903921f5547a38829dca1262d1650c04496369fca53d2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2956f77b913c4eb79a96e5a8911f46aaa8910161319a3e0075d027fab82b5ab5f1f0c0f6654ef82d54b3324a8ff9591e4676b84d384a4013959e79120cc876670858b2b2f5d32093059bf884b490864db328bba59d90f6b04b0e61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5a7c2be90cffbf3bc8436b71c669c1deaa02a53803867758cad7407f336c405d45b7489735d58a4e95675df6d7f39e1154fbd78d349981ea5089327303f4cff9220b0695c6480985c91f062d1a411e397ca2ebe622c743fb83b6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb497c5bd7e3f21b9dcdfa8e7617b45d947798288fa6d876f41c890160dfab35733c6958c5aae2eceacf2048b5ea5fe85dcff63ea289b34619931788294061a0396836eb10b0d5fdceffbcff71443b7eff9eb2d972321c9c27809f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb2eaa5d6d7bfb16323aa4faa79d3a1940c94ba5b681b9a47869f83a973d6447f965c1b7826919bae7b22f2121e4b0d8c81b006a474224f9aa4f4c57af1b336e2f08372291c6494115cd2d082c46f378714afef65b1b724696de07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9061a4a2007e78bb5895242e33059b7b22e4590d85270eccdef701f66c1e2cbf4b5b4b2329e16e4c21b5d5a6db5db175489495b211174e7b2c13a2e13af07cdd63eeeed48b4fe733461c6bc36d7b86ccafe88119db137fe97641a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc0a3e9d749a433aa4bf615b497a34cb715e5b26393f0f1b6bd47d90dd28c08f870f5cdcdb90f0c1b0f9aa8b014ccaf1c012aba1560a8c0fbb02a4c362545401f8ccc3472741ccc29b640f8cb36548f06a2c50836d887604809c06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe85209a62a156ee6c2ac3fda513a3d5c093e69509737b497c7f24d67f187310eea0312e8d2bcb1d18f163e6f2d6ce62ed1a52d6cbd8a8b8303cf853db3ac37fcbfdb9dbb22c925e3c7cfe083bfda675c711c9862e9cd6f88a3f67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbbe2cd3af2fcec4294ae619bb5b9ef78c82c55cf8474202e058f02c4fbc50862fd3a2a0e764deb459a0e0c5ddeebbbf3095ca5fdbe54fefeec91a7c4eed1f899a67ae24621487d7ad78316969307a4a908723e007db6b04bb885b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ce106a422d2ba39249508ae0a15031e39c1f31f4c8b077768929a24c413dcbbace0985b637d0905c62c09a1ffdb8e0a688e089d0c03aa6e499450ffd3b69d66488c966f7a25a5e6d49320e130bdd8ab76e07f63e31866e6664174;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4941683416d8506dc758531c224664efcb0c2117534112c9ff932135acc9f3c7e16d7275c12f1e0225f086abfbec2017ea6c629eded96e5f73d51e3c6ba1e0ede5b398b51bb84b2e120fc6d7db6db28476c8e6243c8c9eb99b33cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ef9ec8e5305d4e607bc6e7d42836c76d92933258cca5214a0d7fd6569ca082bc88e39b2e446cd1b0764a01bb7a6ca46c46e82efa206690e4796c97638df08a463202ba6b4c2fa9b967ad53eb5c5616d19b60b191155b22813261e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1467b03fe66629d6562e093820c399a37e3da3fe0db07c34eeec2369b914acbaca57617bb920e103c04fe4bf9cd53ca577cc6a655fc49ec5d567719c7b5679527fae8c3fc777794944f5da7bf7df53b3ad707bb3d684f52e9e9658a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14355c73bbc36c6e32b8c13f99862702cac281b669ddf55e2ba21f3849ac556c9b3a9ab1480914375b31f81641ca10bc1c35e01fb3065c7bad6f415cee76f4f29ad2635e55ebd7fbf834ad4bc28ea91da9ddb564fbdab457aa6f1af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf630fdd571ac3012f47cb893ce4bf8312cd4ffa33d3990bbeb49e8ee6d2f260e6326b1f597a9140b36a43aa84aebaadf554584efdd75b379fb82d7fa92aa6636bc28b74cd13cdfe745ee5fc68e51e55770c91180247ee7d1d48573;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae71e10e2ea7a886b2bfc6f6eaa18b79142e7e141ee82f0bf3311c79eddc79ca81d0fca7132e63a80dbc56260b2609991fd1d6d2a74ce88b33d627ed5bf763a635ee23749e3704e70d42eccfaf873a64c19dfcb8631c2b45e4b9bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25ca0ad6c8d35fc9541b6e02a13075f73c84bb121cbbd7d14a2fa2e59785d48bbe66c5862fd86722a09787a8531cd28e5ea8d097ea288823b2692e5b4dac1636b279d524d00bb8b7fa906dc4cb13ef0ef74c41789761b3699bd9b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106a3300beee136548aa75e47ac5fdc2912d3e7519d00a5ed75b60a8556fe2bd04b78ed9b26f5fae62167b7b172622bc3ffb50cca3c66136da51fa19f79acd21da9106041580882e06418ece53bc217955aacc4b96951d4df95df66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26a9d12accb3096a3a6a0b97e0973cb792bd84f1b031030a926fb403e2a04922646290cc8b5c1595fe472c6974cfd82529cf002de6b0d797eb43634457fdf4e993b3845c4caedca626c16890c9c0951cc6176ccfb278e9a936d5b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7301b1aa41b90397161d6eb323be592cd4c94f5ff7775d29f5e872c89ffa1fcd5a1ded3711bd8f849de9f219f75cf2f10a9036b4fda6603a138c89d027988288b73706429f56d05f96194619798d03ffa515860c9e345ee1f49fc6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b1b70a68fd419c66855cca59c91a6463f1a8b23eb8d5534a5ea119391018c4ada8e1bdb6ab8904cc1f3e099f08e9e9533ea2a22a09754f9396004488750102cdee933c09bf8748813a9dd5b80bcf4d10dd226ef929d6a25be8a67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18535e276d559762e4aee87cf5fd8b611b4dc241f37e45759a97e8020c3734f2dd4d543521b565305938fe8c7fbc12c82736c058bc25f43e7e62f670be6615c5247e0cd8b1e1c01b883b5fb36c5d58d553c2cc1c99653a847cc835c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155efbcacc7e5258b5bc1a217a974d55d5f16db43460fdeed654b199f63009178e61e490dcf25396bdd28e03308decbf1fea223c07cbba35a0c934155fe3d98c20f7d6251d500cf83e3fbbd557e61fb9d25ad2af170d908466efdb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43ed8b5426ab2e2aa8f8b99766bb678f9ca5b8de944b59bfb57cbe4ea89b22eee8a4220776818fd779aef8978cd2dbb94343a4a943715d06d6e163e34c9b5a09dfc7e07fffd169e7db85142c976e7354e86825af7cc5ba6710f5ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h577b99ccb2c86f4ef091a6f58febcc40f2e09988a69681018d39a596a7795d60f9c708d83f76aef4042b9f222d36114c0962f74edb8729ed19ee289636e7b0b95041e61b9a87875eca476990140b088410e3864836fb78cba98d1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167d7d047b85e0df209a6e7152ebb70f163e37c244707fc9dc3bde5a2da0583e12b81c6f3df2892b95234c2bd5dc4cf025f65136ebf5a348d5404c629e83a9c27c103c94d9ac488873c1a2f0d0f77b8d828c452ba567b8195ad0466;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55bb3c0d82cd22fa09d2e0cd0a9ab1c3305f90009da75b28b9aee95b372c8437854564ee25231a0b0ddf0735d20946e3bc7ccbbd5b50bfe5a77e381a8b0ed258ead976c539b2787c8f76af6f8cfb8531d24cb2947eff91304fd127;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100f2b2f3ad98b218f789a5a01960f73d6b69d927c6beb337f61c489a5cddef0f61aef9fa085ab48a6dd48c90294c1e2c6c8fda5c9d3603f4a99b74067982320a21f57c537023e1fe4523121f36e566e202ca0ca0cc7c16a009c46a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112f76c843c006e14e7588827164bc83484fed3494a764cb2b8d404c598e11aed666e9916b3e69047aaeacde84478c4984d2d03e89d85fdf0d94e7752ab194087175e99b612ad4ed690941f65beb3287ebaaffc9372cd6b47c4570d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd55db5e2dc7ec58de1a8f01b1a19fa53e317c9c5fbb8f46751857543cb6120371d9f135b657ea6ddf7a567e1c7cabfc7a12738958794ecf5f90510e4751d39009200d43f5acb7877f249e5d8f9e3372168af0ff6d8857990f3d251;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d87f18250c2a5dfd41e9d45cbc0625f3cdb6d5d72c179700b1ff2bc9b0e38cfb926472248583c1104a3d9e9b6e81256f0227b57174a93d3bf923861090aca68b5a5109e9db18d35501576e6540b34e1f6d02e127e26eb99f69ada;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14111ec50d9f32c0de437b71a47a379fbd09694535dca8a3bd81cba07d0beb8a1c20dd347587aa36b9b6bdf6e298908ba585128369254e6de4ef8a4b6b085abb2db8b2c6594d7d80f67fea982a2e4ead83694f34d69f72a2b6e55c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11eace8059aedb8e72e8f845af4acaee493fff2e7e4aa43c5849b20120c58c7c271b0a971ab82daeb790b9e50e2fa30619cf6b7e91265531cf1406dc3df17a009b6c902ec81d6e1922c6e510230144812e67756bf39b9639da3c456;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125c1f8d5207907ed69ff02441c1d18c509e51006f3092e0ae559f7109f2cf30cbd07169ab1e8a74bf0acc939484aaf2e4ebca646f8fbcfcf3a68c79af5bba9ed41509dc5aaad2b8ac79b1ccc9f9f1137e6263cdb86f0b0f53a4a6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f2e98fa0611c70653206f189334d5c7c8fb737480dedfa36e67a7a1d9c4a3d56cc07bf9ac5a86362b6cf465bd77929eef1205767d7a55e2535f04184d6c51984e18596b598c5cbf0e75627407c10af7f578dedfd91901f3be8558;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19268b2d7d7a988416f587efce13571d93e39a5268c691b10168d6465356a2fb3b2967b27eb142019d42904ac48b0ba505f21a8a48d71f1f479b9bf43bc45ca7ba4541b9678e23397ba70f20bc587bcd2b90ffb905f30f7b64342d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f3406da00382be7629c21eb24f1b22195a949ec956c075117ba416ca6676bd61bc692408df0a096aee8c5928a3a5dd34c49ef6ed13c966211d269b5ac77e7ccfe30aaea231747662a1016fdf55d4a95601ae1eddcfd242a77d078;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d6fa98542b5c7e321f93582d2f64a39eb5255d58a2f8dafa71363e9796988cb9bb99cc7718f476bb38ce70cd480386dfe81cdd5298ef8fa353f149962d375ffd0a8c4d0e680e18783a31789d3b04dc77ee7291b91deb184fe17c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf092afb14cfa6e534e49535c5fb962ad096bf078d67bad63f08c89cc20da7fa8d81ea381ba8eb80ca239dd0124b8bb8845d16ffff40c7c2ab1a88532ef1717126950897da0694b1a2bf8bf6157456c491982b8a79da6a73225d288;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8857cccf4c317ce20b7bcd447717207694c118c02073af21f5ed347fce540149849a6c96a38c242cfba7927caaa3df6effb92879e3d89035c9deb60af56aebaeec39be7a95274cba476db1424ef8345283212d794aea1843e577c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15200bef186dc82e4f5fc5fbd2a4416f63a1194948e07e2cb6cf4944becf635d70bf7f818d16f551d05e4d42fe9da8fdcfca6ba812bae13c753e843a809146b03e8888989f1bb7c836033f22b396ca5200d090fa9e4454d2c31983a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e61c5f765251deec3f1bc11ecd535bd256dc1a7c77fcb9192750c2cfb81a5f0e3d0a043a3e6aac8235cf08e27800ed673dd981a7fb6a5baf7674030f3472694c2f5731a9079fac2bc441bdd90adf90935a5c80778185fafd25d2a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc39dbd44f92c5fcc5a452d234d2108d62ddd460c690be4ca37fc9af446ab470d79b28b3513917ffae49f6011b1bb1bda04715d38172181a410cbc816b10b1f4160a152e2c6dfb3e6d8197764490f1b9980fd6328797d9a1fa9fb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6c2ca34fdae73d9cce7f63f8ae83a167b3fe82f6cd4cfa6314e27e1f067e68d6972e854e2b496524b5f543b7c7eee14e5199a9fac2ddd4244f37842b13cc10fb2d3fa85299501b50ea65c1ccff0c0e73bd6a2fc2f06575a335f13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5821d961093fa8c0a99f2882caebc7ab76b7e409ad73b689d9055ec7dee87d9a3b4f3cf8f0ad358f4fe1de53b1bf92e6dc5d4cbbf9d30b5128ffb118916e3e07f68bb8d4017d806c751bdd5b97f8d59bb043bdef3d8432df001e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1696a23d46b2f5e67d700c0ae9064b4dfa72b2dfc055b09c3f720b4eb00d11fd4d6b0e7726230a02176da4989c67c7a4bc63654a0584009a9721f8ff393d30169c301bfd164e31c13517e1f0f10099609fde9ed9443d757e93b1fca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1deed732465b45bddc370fca96136ec498b6a9d7bd9cc139d520395e87b2a27063417a8d0dc6dc4d3e4791e41cf175878419e19a4afbbce1f7c513471b103ed79ae883041961a0be65961b85928fc4a41a53ba93e347f97c610f19a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1970886a86234581504d7880271dcd04a2870a32eb3db5f12f27ceecf0f4a725ce0f793f3a0bc428c0bd4c4985ce75906082627227694cbe23425d41f3ad7275fb53fe40357a42c7f2004fc83df1fb24cee5c341513b08e5b910856;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1432fd3414e4f36d7a3d88cad55a0689a073018330afbef17938bdabf187b31ffe69180af49feb44a547c29b5c0380e86f7eb46ca4c12bdc0855dd80dc1d6b5dd32134b3e9836077cf5c920f00bcf36b120c8f2f35d1eb0951b3b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc69cd69e7b84aacfed99e057b3ec397302fcacd50eae918e9f7ef5d52c30db48cd5c19ef7d099e4715669e204166557f9a9dc667ef492c178b641474b2fb9a5f0ae4976300c664c60d79afdb4cd80041459917cb958b8cd4eb794;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1600230033ad972bff17947d9404b018adc3bb8fdc9ddaf3f20fc52f4b9d16b303e82796ccacc8d6bb182ad27698250f7e638beba83f0f2708bd3eaf0ab0ae167f2102d1ac5afb9170db9bad24178b65cc43446224cd2ba124832aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74824420982ec3a6b9bb2e66e9096f2bd8dd1990de7ee1e24f32f3e99a28aac5fd7ceafea14eee49047490b350b82d17684187ffdbbddacaaf3996a291129b906acda07ad443d15c28ab893f95954676d5179cbdbcbab35c27dc61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15876f892b69c3becddd3182a072cd844f8ab54543065138b1ff8cb54b48301b691cdfb5c49ba2e30d8bed3ae7b09cb472992fe8078a4936d99e4b859bbe18456f8a771e56471c51ca2926de4c3d8d2aa135ccdaf791c02e14eb44a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16303262222c2d79f881192a5652c1bb9b70ce3feddc7fd9d52dddedcef3be934c6990031dd98d3e0cb3dc5a6996e31dde7122f44779f1bdd7626323649f14c47725c71bd82b148f2699cf106bef909da1d695333681402546ef7b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e04bca82cd87ac40272034a11a846ce5cf8ad5632c418591f5c2b7f47547f3448303f84bf57b9d10d33df056da605df2d92a6278430b00f33086bad12616385474e03c657c9d201adab332b04c0bbcf6b4d5d314c8820a60ebd80;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3878ff55ac68a0c340f230ddfa8ca8c331960aab4c0f26fbcdaf4383d36cdfc1452735deb798f2479fca396e47dc147090967dac56f440d90fde39ca68826eabe4339778533d1acffa2327fd0a4f4966d07d164bbb41b65b263ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ad551c41410add2cdb9bb700fe9b7ed6c371046550719352be10325a0cab809afcccfb49e933925fe4f25bfd74f01c8f6ae2c3cf7ad5722a7bb2faa780b642164e71f9c0fc4b5de70ca3d82dfe15e5241200b08a5fc9267eb0842;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acda3cbd84eb3a618220c5c1480fef80b5652901987494fba28fe546f7d4edd571b0acce42e015165e16fd0acb4f11d0bdfc01cd7907ed3bfecb9bb42177de5fa2ad960bb795bfbc21c0083c670b53392491da19257587ad2d233b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131e64cd45d988277818804d03eb1b52709cc6ea7bced7bdaa96a29b1f1868067cea8a693ab2b35c0b33f1aed312acce32520c7f466b0b3082f59e552694a22b79a28fbac56e89f20967039686e4a8b639f82cd85e3215cb203988d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13638b7dfaeb1e1ccc13fb7c89357dbb8c4964858a7c607569665bf998e120bd5bb0b4899ea74ba4552acc4d8e32b34d669c40bf2dd97626fef9d97aba94e9cb8b42483be55db13cabc631fda68ba89d93054b9d9ca61e6e9ed93fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6455b76cfcfc496232fe596fe52da96235d3b0997a9f78cb579f416bb5c3a0ceeea264fb5a9ccadcdc4298b7ae38562feaaeee293c0a104870b3967a9bbe81f0ddeb2b59eada7525496ffcba65188d2e6f8afefac63d6109a29033;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124b7cbc9abe94cfb1f30b25bdf6455839cbfd34311f7278b873932cbf3f31c2944c7815b7c1ba1515daabd8d093b7d16a8d8d76304a23c7814335d5afa0aece9d57d96f088d5a347ddf5263030432010fe6add822e5ec1ecb59917;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6dba39626a961efaeff863b30a7bec8bb3b2f6763b101bfb07784f9738f8b5a065f276de3135f9a8dbfe1447b8411a89aeed425f33f121d1fd3f7b346abb5deff0006e94cb27e915b96a2e6a2a9c2e2b978c114bc80d02147834a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2aef9a2235ba6b58628cc2f7856f8d4c3dc882f67332829592a4ec87f702830302bb2524983a5d185a3afb12894d8cb1a1c0189030598d521cbfaeca447b66f326c6347b4e6f2d9b62f79a73550e58ff6ff24533ec1bd037dc169d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf86537366e80fef6ea4db8625515bfb5c87d185107cc872dda7d1c9a6b7c853ecaad747c58e017d25b21b0e0ba60357be95e987d8110b902d9f1461129440ad2650ef4b9608d6486d1d4882ece815dcda0b3ec92ab9ce2aa079afb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4b56241e02651bc976a61f50a9b5f45516b12b5d1268e7924cb932b3428d33ec491bf236c263ae904f4629e3dab0f3d9245a683cbe582bbcaf65bba9bfc0024fd82a87967af0b2c7cd3256a81271b36dca945b3bcda9d1b773117;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b307f36d35ebb06726bf7b8836daa00dd7f3383edc8a523156641a6e6eee1b116ded45b76a757aa566b4460cc881c073795f351b44a48feef4911ee2cf3b63d1e9c79a78a2ab7c20489170556eb8182b2e5f45709cd83adc34d711;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fe66a6bf93fa2562c7cc6b4b8cd2f9dc6d89580adcabe983f97896d8ecb3545bbc62449fa3dcf57719c2ac65d818a41e6c46e3bef41ce5e3b38dd8ac20c96f5e4131bab16d88929c2a13b8e53a355f63d9b7fcbeb2ed37677fcbc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75885af3e13bc9eb226721c6016aa426f4da2ec4c4d3416772f6cd53fca5f759dec743829eca582026568b5576ef3cadd739bffcc22a630a9c8aa1fb73a2c5dc0fa6f44d98c654007ec94378083e200c2b84f5edf00d21e9b3dd67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14fd82b5cd004485cff5cec8d777e2f1e2b7ba22fae9991285dab0f047c47aaef6d930bb1b8e99fee8cfb8ea2731178fb9b64f9aabdcbf6168f9110e2eb88c22603d6db2a11d5913d47c4a55dbde413d43c378ee65ab27d7da4843;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7beb9bd22001b6b204f01f05e6856fa3deff42857ebceca8afc40f6932db6fab715c7aa06a66f3ed0f7e9912173d7e173c3476e654d67b78a4a37d79703b2d26d0be92bd840bcb5a58c5714f993c3a6d5c984a975c9956bc0ed98a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92b32a89198aafd4804f8ba96d1b22c25ab9b368b7a107445195c04ed9208db340d437e38aaab02177015e420b6ebe1c516d2ce1df12827f5f4d2ac1e7287c421a7461a0fcfe62aac12c54fcfcc2caf98c9e6dc7182eabf35acbab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h145ef4a57b60c3b9db1ee4a06d8533710c886d4cde6ffaa0d793cb06209346e9cf37388155d57586110c2637f2da32ba2eeb15169710624af318afca43c65780a8c804ea8b6b7ad1934cb24b8a7abfe116e1741c9dc1be60f235753;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f50c4cd8af23bf1b8398f19f621b554600498c1cdcea303d6b50b9262ac4f6167d4d4e692faacce784dae68caa4d242f65b0c79fb4c9a75849d462873f1e8577453f9944ddf053045437fe1fad4a16560d80867be9da23dc2e9e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h494cbfca23b4e39029bace42075afd2a3fda5e5f8d67d8ba2d1f7150495bc20a2bef295fb79e351ef7e89a580e6a80c9c620140a2cf246c6c634db88acb343e6319bd19f2f55d73e2d77abda427ba70fbaa497b8c4fbe11ad2f801;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69f12a69418897728b837e71670f457cad12f70cd0c9c0b09bcfb6fa79b45fa0a741795a33943d3bdcb32dd678689ed030d727c71212dbb646032b16b7bd6efbc8eb965c2f6c6640e68cf1fd362b98017900c66610d3ddc6d4242d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a8a5eb73f560ac873093e74329824d54bc96272c14f5c895810462834e3b2536a98c1ffdc42bb9510b3a1478718b38d6e3a26e91ae9528ad14de9115ff65b6de14fba5bd29269ace5b008faeaeec2706525dbac4616858cc802be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141c7bd559c4ef897eac58b02938a54e4bceac74596c98f774957bc602b49961cd067081f889ce7bf039f0551858a0f4e19335be3ad03ac23bc721cf5ff7a0c652034c7df2e5709249ee2d0c180f17443767b6fdd6e084f29d3862e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46582a27be5f9ff15d36afe8add5aba3584b1bcf5f5df3256c76a593cea2e6ce5fc76c5d5575c1ddfa11a4e68eaab5a8fddc79446c0d82f032c23b2b9139bcb69f67cfceee661299dd508b4ab011f24fbf2ed76770ffe95a22cc4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148fe7874c13bd74ec741ed9e9390ae5356218c05e386f14ab4f037c5a8efb2fdda5f933c3a0590fa0bd9d58f362fc1bab91a00937a305c14fe2a31fa117a6bf671bbd464625382291961771a8d88786b95a95fcdff9ee16976b402;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c28207a07313dd7fd57253bb4ef9e1bed8c70568ad53454740c0494989a82ad3a07097c58d66602d6d07e1f3889f19c7d06ecced9d506dc780276b9e04875908e2997114cb4937e994960507cce55775fd71b0d4c14180948e6ae3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3987234aca7593f993b77cca5cf7e6a4c8137e702cb423b3053c50b8e035e30bac07613aae906cf04a52983d2311e80149d5ffdbbf208f9e786772d209f9ea9fca10839df6bc4485739745c57f63c9292da4457639e790e75bd2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcba1154c25f38dcdc22e5dde749a9f884642329f21090adf508c7867d875b8dde25e6316cc3af7a141846a1b3f79cc63956ea66ddc17999225cc959d8712c94787aebc918944c7c4cc8ea815e67c3a0519d11cd03e1045aed330f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9112e6fabab3865a68e1f9754ea87cd2a260c8ff80efeaa297db9b51db78e934e27f886ccfeaeb2fc5c07bfb3d01697bbde73a1527f18650938562ed90690a22502d78eaf1f8c99a1831d5690616fb8c65fc0c84753539fa8ade4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed341f3ee00279693c7d761d6ec7698049a6cc3fe21fc049644cd655d0a7a0d684a5836d5c1950e995900c2b0f6fdee465061c8529f278b8723cfa3401f4ec6b2a126252e019a7a070854a646bc1753ec12f17bf58ba756c62c379;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b4c3dfd38a2b61703779064e1b6dbbb98640b67fd360881b62c42180568c0fd9bd4dd73a7033d24be983c383d7179f6f1d44ba4a9d0ee638e1b5e7d8b43ea89f6c6d3e5c013176c8c65fdfb81cbb574f9cf742970eb9faa0a4167;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59072a384d4b78cc3f848f5203bd19cc032924c89576912194b1fcebfd8fc0e034a073e8a83cc2f484870d3c81c1b440857c60ae84e6f14f6b544ff0964fb14ab3b5d732a501b562cf062cfcc284147aabc20141aa88f091bfff04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc5414c80639193e879649219f8a54cc580bfc40eab9d4e068f8c2b5ef9f309f72ebb1aa5dd40d5d58061306a68cf1116ea81b9acdb554ab39ec6dc0f483ba83911a90a76b2f0f32160ca53676f560e168f662d5f20ebe8271efa7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h918e60e8edbf85b5a15ffd11c60df924181ee853fafc8ed687fd10f76f005185d73ebf5c5dcbec25eedc29efaadacb4b414ce329bede5e7ac34a007dc6375cb68d9b3fdc4cfcb52f206fe78e10ea2fcd895539ea518d7a93bb0ab2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa340b209d03cef543649340204431ecd71f4504ab681d13714bcb49ab199307ae15e53cf867fc0cf84264b2f2a40b3452190f9b4402a02ffa8a323a1e48e4e880cbb92abc05fee80ee4199fd35f98789390a7966d597dfc895294;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7d51ed69b5c4cac5f8b85a2098c401df28b11f06cc71ac564583d407cc40cb4fec70c585c35a714b211795a71919a49b49ebe2353e1ffd1270e661bfc9a7e2d3a92b8262484ca5bce7bd74d1a956280c24b623e102d7551892697;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haeb0a043a9e507cf34148e03ce4da6eac5967d38967ad436b1c917ebddc0f6bcf24bd11bdce110617746eefc9cbdba549b858e0ac08317b68f63f267f34c05db32ae51d5ffa8d0637dbee26c90e162f33e64b21a057df89e7f136f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db01379a8b8adaaeb4dd475f529be19552020c6fbfc0dbc146e763d1024feefce69863b2c8b4fb0978949188cf3b4d4445409e51484a78d6ab8037eb43d48c73be6a900cb00068222d6de43c5140ba31d63af1721bcee2ac4f4c59;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f24c10cc430246a162157bba3e32ced65d5415221bba4a6a9cf4e8e0d69deea675ba87c89cfed5efb9ca381de384df1013b10a1c9ad58e760cb90d20bafd7177799bbec29025b3f51636755d7b192e788ed1cac0d4ef6d91e7100f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9cb21bcef869f1d2ea04bd81c7a26fbf98951d3a0b5871c7d6d7ba2af3c8389ea42b67b5eddf187c61694caf712b385622b320c6bcd26b6c222a68386590910ca6aa779ccfd5a6336275a57a97514a964fe21f93fa9a933c5cde7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27b167da36e7c8c1110881c243545e5b06756329d12e387d84b7efd33fbcf155818c0d1c7bcc00516aa0ef8ed888b30323a2b829f3965eb5714603ff16be4cd00866e430ed8ab4340980150824ce9765b59281c192f669f39d4a71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f3afceeb440bbf4188826384905b9b1081a8002b4719b8d12c2b8b6248a28c75053f6d6ea494015d6bae0dbee02e2469e2cd8b23a05c2f90e236005e29c71496c6965685f70b72ec70f2a017109921501557f664399e4cb8ceb3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8c39deeb86372602abbf8d23edb3d1150bc031e8b36d3ea502d93d799829d51e0fe1907a407132718f5de5bb636ffa25ed3aeda003ca4cb9e1c80889adfb9561fbc0dbc9253922a9fecc8cb6ef5f2d8357717667284cadb0b0124;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0fa92002e198441ed86aa7f45c90a6b25605fba239b84cdc5d6151f4d0dcfff04fb5c6240f49dea6d32c3350bdca84ca219b6b640fe11c6e1e5f2596ed5773fa49494d14084ebd5dadab133c9e71f1bae78c4c950e1c065ab02a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d888a3024a9ae5ce1ae83077e323c3bf8cb5fca7e86ace57d56f1d054065e9e03de2b8b371a366721b1e70a1b680256ede1f2a2f4af2b41e829e8de1b0fa0b27d374ad1a9bd88cf8796d5f606b89671da9dd0e6e590fde937f9e2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13873bab379239b24e439984432d9025db9814dbe1901f6dde715a930787d9956a5ee06063d9ebfac1a8682448ba6d56c9ccae14f76f0fe54d1702c9660e2e78ba8d2e8190fd23ae789d5912ab1026d8f4c1d0085fbc31ceb6dfbe4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116fcc7c38a9f53c211f33794e52337b5f575e8543e314459f3925140b2a426d6ce77b8004131e0de3aa230a5a5a6308abcb3adca6786c4abd99314aadbf21148566be5c861c2e30252cd718d970f789058d542bd7d2e14b6e6ef69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ffe0fca8cb286003f22ed8e0f7331691e57a48fea5ccec4c06dd4dfda43e46896d6cb9faf056a05504d6863b4990a77841a7ddfc9f2e08953a6cdad2d62b6acc3f0a10e4db6e7ebe492c90c38205b4e81fd0fd83a32526b36f501;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h600723ee3c313695cfe6b8ebc2342f7f2da37dd0fcc6f4f5f7ab99c61713f1d741c43471744881b14155e01531fe0c740caa55a32c3ba75cb3458f00d4319a151b1d930052d001ddf169c445c37aa297674f18b1e72d01047eabd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8cfd0477fb09e6c9153b5815ebde55e97ddb8763bf204773652aa81f916ebd9c5caafe77a47b37773a59548f1b043381f42c259ac8a8c3430a3b72a5a87fbba0f535400f75df2f3278da9f35ac3c95d78447e0e6d12d3a9442104b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he755a67dfca027355c5d62d61455e5d9cb21014c067ec6fa730d5cfba98479a2feab7242342318bcea36b54b32b1ec4f62c7c2810f27c1b552e63e68a726510196a3efa9fc098fb92e0fd135d7615c61da5bb722a85582e6635551;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c89b35a94bb36c7393b3598a92691c79d8d03606b3d16120b419a6ec8e999d9499d74c657e9ee4fb0113e327f8d260a35d5a6506ed86e5ca5ad59015439513927c74bf7c389f3022074544ae323023fee8e755fadbde29e6ad00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf473435204cd9ecfca8438902e247fc2b576f6e3f04afc475635bb5295bc68102822b80e1d05897f5cc2d5ddbca2db4de055f9fd12cd278a72a7f225ea487632eaa5698732aaf572897136bc24ceedb115966b3fc102953ac084b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haccccfe61c0902e1ac484142f44e516539b3f78170bb2ef6fd005eb177e22422bfe5dafb7a8c1b0814566f2b10da6c3a481c2a48a8a9a4bd11b25ace92f2762cae3917748afdc39bbf0156b5fd2f93d696a1da1da984d63c6d479c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2fd12bfc1583c9b9ed2e5c395ea0089e8c3b890bdea35298d69542dc5767e9dc95c476e2b8a8b15ab49f334ffa7d8f3c15cfd10a84834786c2b27c987e8bd920a2fb2453436468e3cdbfec69ac1df25094502acdc39072f6bfda3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10078f5da8640689cff3165cdbf07d34343170efc718a48704b54b78999c77e493d56a8d8ab68fb9fe289c7a0fe8fb383051d5218a22a2b3641235df62bdda7ecddd99fedf4e97f4ae85fade32a2bca60d2e94f40ad53fa6dab63f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h618dd444d96232e0bc2b1ff46585a2022bb69e3b4b6fce5e4458ed2029e1989faae22b838c2b2fdb89240d0a13fef9684c15840c58782d7a5de3e0ae03c05a956bb897f6992bbcebd6d14749784894bd525c4189896259b57fdd8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98c7baa82a98910b507262fdf96f2380e36dff1209a5c8c0ced564f493b71e4fe5507eeb8e02f08db24e2a6fbb8317bd70efdbfaaa465dd4362dbc7525e44a6f68708743ab814fcc297dc954c3e802a93e9518143df6d494521faa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14361adb7b490466cfba7a129a3ce015a874697d7c0dcc1d96ec6b6701369b3202f1e19eef714093feb3b5a7ab1e9ce0be3206350716e5d49ea558d3392459a58a8ffb93d54c3e370c391bb6575e9401a98f6598e0553869de49c6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h584f8e7db26223dbc96495d29382ab806a4beb0064466c9223648827e2b3f8bd79c8b751c7a23eb4be9b7740baa817836bfdcb4fdb62610f29975f94a42b303ee4bff044b294321fc86c5452a0f8e6bb0174e0afe85d25a414eb4a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e805632c0a816b342c213781a737848b099edb1f1b354c8f8ce75c8f4bc9a1ebe6ef14f6be6c69fd712681dd9c3c81b49dba15088bfaed2a4ce5bf222869a467a35046d24e15f4ebcec5905beb8d5efab073903be4501935d7d407;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7f8829f6e1ddba990d326ccede407d6679971cccddea6f70707f3a28704527a8056c9deaa6d3c5edd56ee7c081e80a3c51c1f718148a79d5c18a1f637e5564c59fd38f14b49fbd43d97d73efb18e1716f9097e44dcddbb2973f0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13517f6d1d08a66d6fad1de2a99c204da5bc259c07d465d39899098e378e6f7eeaacacb0e19fb7bca6cc4691f8646ff4332ed188f59998665053599d164325f7ba4e739dbcf58a99197d3b2771aa957bebe9772d6ef6d4602cb8bf6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he252d77d69389ba0a66e8a7ebdd48cdd122d97d535493eca8fe87e19a785f9932e1e7ea84e1444ebef5d6088e29a1bb0cc7a5fe70b324aef43ea05e8801f0b4d6522585ddee0b63dcf8a04acb9697a06a9a37176d7d4d35cb85484;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7505dc287683a14c6cad2c026ef4b8738b7f6b2c212bf4c4cee331d736d55e618d67ee80b5fd0293917553620efb6642e57c4a343343a4db18d92cc75fcb1d12775d56c1ba945f52ead17dfa7ac4ed71c59b32328ffef8278fb19b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6dfc459a2c5f142793897d438eedb36dad510cbaa6ca07d625b018cad124972002b1807bc7eccd3e801b4fcac6e4b463bbe75b58afcce3fdee3e3a3dfb82d7d092a685bdc9644c79179480944c9a5d3979568a2ce32aaa051715d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ab2625f9e48077493e50778cd81ea050de5e9a53b2010595d20696eec5f2faaff4d4035b3c1c63a7d76c9db6e75c68c8047f94516d2710de63c2fdc6ec0260ec2ce21d1cd7221890b2d70c20454329374f6126b52358368bcd62b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f22e32917d6198c742f8306c89cdbd5093f0da6b4ef3fee41204a853283aa59311e7501653cd35ead0e00e6a7ec64e5ae58251d12ec1dd40bb118584ea3c08a1eaaf779ed8c4fb9d41fe555635d11803cfc4d0489f2cba18f5eb04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha09e617011165d8ebd6c507693e276c88c4a813d70e5090d6940029df04ed81c2f43fc17960e027f60e4ad72a5d18f8e6185237d7e288d455c4457bdefba9f3c2a6ac6f3caa85c0e45a7217cf29f7b178ace3b909025266b77a703;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10950800d355288052a4803d4f14e2898c33bcea4fb70cd31411baa3c63e431c4add1cf069fd5a667d2b5d7aee1f31e22b874201719281eda84693667a232753b835a66d27d9cd906f5eef5fe18ac6ab71a1f4de81f331056b32539;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6cf90e63b4180aa0585a7523d3107d478972ae301c486a2c3eff1925fe5e4e55384ced96fff41afbcbf63a379ebf26566887d4c101387b7a7be4e4dac57c9ba503b3214db543ae4534b4437db3dac7b3a86a66652bfc6da24f8c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82ce6312666c035367b42b67d799592bf8ed042a12a98337b8817e929604b0ddbb4ad38635d769a505676ccb7b21e2f9690616128f2568a7fd7f38f26fffca15f95f2e971057de1a1558471dba936a201ecbcfacfbf45bf2ee75c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154ca77d634b60f90599cf343164cf5437260f6df07e6a43edcb3e57a3816bbcba24dd0c7ffd6e307d3c686ae3525004ddc62ec2ba9702239164084d0a128ac9eb2acf6775aa3d658434dd295b6d6c7811e8e3a689ab463e82d6f29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0bd584cb73da1d8f4e25b35b480af88fcc7f8cb11a6243db2a70eea8934bb33bdaaee4cf95ece4fac6205f49ed6f1c7ca36596394e113e7348d789f51b4335d366bc1030fb386b2ef41d09ffc5b14ee2c5d686ef5558aca3a3547;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d384c9fb6cf38a92064db2a3d4af1160d9370efdb17c8bbddbcdbc5863656302f6ee86b1a2a9ba012c64b39ba44148a06fec47fef799111894d8e8616c2bc9fedf1989d3cde1e66bc683e984e703317eab7a360de7ed579691732;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fffc034daa2ece89e41239ba118b18dd9505fc5466b663e17b666c5d54f2ef8010e56c9991e06e6730206efe97e5968157f28694c22f367d362538fa536fb15939368fd962c2cae0a77f7baafe13b6764b32e911e841b86e7dd32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16711a220dd9a1cb97b30d7125d953bc8650aa51ba285be526fbbce427e3610c845f5e3a03746c94c49367f1f8340fbdad27ba562471ec4cb7a765e72e21836974db4c301410a63be10b2fa4e93aa772a2a3df4179ebe0bd66b0027;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160ed049046f983ba13409b3eca2cf8d9bc1a256c55e417c495adfdc342dfe1e9704db7c55b08ce03058323ab02ecde167b4448695f799ea524c4e204eb1eab9212356ac355987dffdcde89f7d7adc14074569a39229c6bea01289f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a64f4281daca92638319f0ac3f4d956a665d65d583daebc7ca696fef67be0ab75bc41c3cae9af7e261c561f20b1d826434ce084bf319773e91a9fa5edfb4dc2bfe44cdc1f27cea6eea958687220788d9c09c590d48255828bce08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcd0b229cada4e0f54864ca3fd6f9e2d0ac5249be65166823308aa25330b3424a972f5c273ff15c1312b94257876796015201fbb8bc5b55dac3f096a32a300a6aa8504f2be17c59241c22f885569fb2581d77a0f5a15c868d6a0ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166f17bccd888569d5562df46818e17d4fc86d8a1f353ed3fc671574ef20270736d60a193627c411244f1c1b9f5533b1d7e5c3ab8d6e53bc3605bf82848920acd6b86344b246de06c6db58872e244d895c60018ff3d2a3d3fca9792;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf84fd5281b511dc03f8f48aa0859c5ace597149e09adadff647281071ef3d02a1a1e737a60d3ad9644b605a60730498735fba13ac9e77e1c23790ee89c8049650fae213bf2ee0cac7fb5bcf307ceee14d40c2cf79d3e9a4fe3e1cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbca3a3a5c5619ed198c07a7ea080225ef4bdf957dc551fafd8593f8507e11b75e476ef2b3cec3fa62834cf94bd98c610e6f5b470beddd44846f6c93e364ebd7a4b25d0092308e9c4e4e479d76d6b729c96c0181625ce42de56d16d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5c35f36c259a8333e3e7a1f14f29cf237006e105060f90950139c992cb717827ab8921b2014a0aae39bd414cce464332d2bc852111dd2e33da2f21f776ff71db36a3f854c16ed31f7b56865a5a21eaf21261ee66f3c2c51d922a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae4c4f91b9d5970f7c8f5e38b7ebdf5dddd4396518a937d9412272b14cdc84ffef41f0db0bf3555d8cea3520665ca1665a974be248e36412ebe69fed47ceac8c6872af6e6d7e183d1888a3eecebef0d62f3c404ca9b4ab6f9b9271;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191de31e2eb092926583a1ea471bf9b9d47328216f7175c4cd1b3a46530d97a751784765850dd4a3b6552b907158e344251bb12d112dd170a112be623b6fc709956a22d448f498df3ec721596c0857d89da55a5b6e7c98a1bfe1a74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37afa72e65f4f4a6db01963624112944130b7b74eecc5dcdd518d92ee5e011508dfe00d8d169b805344d84f9a8e425c991ad3810ab84dfa36ce7438180aac4134ca3f8318b4515ffe79a74dcd2cee3ca1a42ee9f33596d3d232d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13780f067a471ef1a159c003eca782049181bf82643eef4ae158b46550931152286c23545b042f230d3c6805fa231120d0699a3ecdce25a6808e9821e5df78e868568d5402b6b46eaea5edf57fce40eea23629e2f730d53115f26f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9038ca62a9f6bac9dbac7c94ad52111c6ee0dff429c46936d341312f8fd6882de3dd81169c81dd06a215da62ea6c4aa17a5d1aee7188655f1175a606e600a1a812b327c0c0e0697832c54f14da1a80a5bf9bf4c22b417b527e1b8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a91a6c6c1546309706415218d50c41648591ca0238a46e64d0e3d53d1ab5d8f52a8c72f185198ded59fe83bffae21634370c35a7f8bcdd3c6d3893fcbbf5c73a5db69545bd3afea5d8ed5d1d2ad41c1dc9c1b92c1047dfff052fc2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3fa1a9ed35d4c415949a9f71269d3fa450818b4d842bb5896fad4161a847ebf9d4bdb58f4e169dbc11f08d12d74dea3fd6336754700d5be3d3b71c9fca7f414f3bf0c1a9bda0173010dae0399483d92e2f5be9cabcf78b152fd51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22ef4f9534d6762b0e990aa06dd8da921e12c6a6a1805a3ac4b42c080aa01f591c9d977c0d8f9b4ff3719e6ecfcb6f8e402a9e788544c6a37e28b5496071eb3f32a0aea996dd492b699fdda88fe87abbdb7d790e513c2fead3013d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heac94a1ed3cc27b8553960eb9faa3d52ecb27152ce17859e196ddacdc57331e88f3aacb5b3e2f3ac54bbba85c177e2c69f6c25cd281afe2d64007e4770fce4c49ba9091ec76ced3ecf306f42ed525e316d95af250f3d76b9f68b5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d38152549bfa9fa718a234c6d5af3bc6606650c920ac9a69413fac9f1fa9a4e2933af8464f4a047d4e34c157bf3846c3bd2137b4dfcf7dea4d39a3053cdf971e7a443139390e568a7772e2ba5d5735315e9817bf1bc2287dd2376d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186485ec67df73f87b669c33c62189bb24ac72913d4be505bf3e56f1d1e9bbed5e51317fb3c4062f64da5615839551f7c4d5e82e5ac5021c341ce8aa2f28034df0ca397a3cc57126c906d221f621f05766c075f83ebd9a8c3c7a4d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b63461d9a3491e234ba7036f7b204787a8c61a2d0bc01319d3ff7cdbc63b8d9fcf30dc25c79e249d55657dc55501be2c23c66c15c405c781845741cfe451dfb8765c6fed39fb04e28d112985937884d2646f67b71726e5db8efc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa2f2b0397db8f491e277cca6e447185c74d5cdfe1f20b2955c8e8ac0dc38df45ca6ec5d93e9ab3eac53ba4545832c0ea3aea288afbec1eddabc1217cc0eb0bb5c632641715d63d963632dccdbda87c207ea02c28b88e5fc96e526;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ec53a3e03b42df6bde85b811f04498a911cc0502f240e89794daf8df96e773b5eacc848d84d568cdddfe1d730dfc18d91437aff104ba7b4031ff1efb1c32a5cfc246093aca239b8454414a4d510c16ad95c830d38ee59c4daea34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19644438c4e3673fb09fae42dda30da14abd8434f4fcfaa6e5d75f5705c0a581f1fc12c3a2a068032aec2725b2c0668eb0ff59a3d7089b6792a647f80a69fe085620b3baf08eadbb2ef6ed970824141919350608e5bc239aab637fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148054f70662372da4587ed5bae5786174091250e19170e8105bd8d3958c2946f4599dd904c11fbc707dffdb75fb8507b8cfe2782bdf54829a64936cf8e6b5902af6dc16915f62594edba94fe2e8014a76bcb544073ea8f7b76860e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fe15e5cafc4d0032e312867f6bb980efa8b6928097b8567043430f3fdc07f3e9821dd17abdf980846192ee00fd76325687edb8c91206c72d24af151263fce91057ee0c99daad5a37cd6d1313664ad5a099394e26ffa01a5a0967;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59db57168a15069762beea900476cc459306a38f53d2a8316bd826dd1bf4d7daf6ff017a28cde5826617739aeb65afe9b659d83fc800b3ff919499c6325deab379b2aeda9e4fce8775e8f4f87dfef7524f6da61a936fb9d7d7a16c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h424d07b6b998c1970bb73514e5c880f661a1b1190f3484b33c7f9578cf239dc13d1d7b0c55eb860a149c758037d652f20843dc3daf66f5432e22039ea65aca423ecf65ad0332f0b9b2f8aba170bb4ef9d7b6eb0a9a17aac275c43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd50b90b1882ec96b2e4329669f4e842139b8e0220d5cb527a7445994e2adddecfa3f659028c42f931eac9ada41852dd716579f7d98e7d3f323bad60648da4ba4ae4690c466234f7959c54740f0e787490d536d2a01cb06343ce967;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125025d1f883ccf632b4bd1e459a794fcd844d67f38f8a2a3fe62a5e10b9a4095f0dcc4862a2f41302e7c5e9286486ab5e15f4809f9a00be6455afad527ddb3441ab7598eda2308ae0315d0298280f9a63e7e38fbd8de8ff27b1c2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94e1a1f2f460a4a9d4a73b74ddbfc1a221d1ea58701df6b9b0bea58fd3975a38b72c763af17d9851b749d6c0e23e25d8b30542ccbfbee2e3b6dbe261b5af502de3955c19d2851cb9fcd4ceeea9794fa35025659f19da5790fbab03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d3da0ae079d5ff03f10a1ebb091670717fe9f141f61c46ec0dd53d04bcbdea79d7c9b5989c9c3fc6ed52fb8fed36f4295db1b4ff67f7bdab8c8e5b42ecab2f436a7b3e24292f57da2fc67cc37220a807ebc73b9c9a2453476d0d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h531ff05b2d6df4a6c4027a00e06052d0d9db20b0e61663d76a22ff4354ea481877d481adb4eed9e201ee9b23085f7dd11bad62c3ddc015bca01b670cf4eb78abc3d6ead72cdbc9f478bfe3c6285c5dea8bfd693b5bbf2d40535bf0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b382e37058aea6f03f05e8b602b92a3b60a12d219f33aaf0fe2767ed5e664382a47bb1df0cfee6d42e00607e7229bd97ec71b2036245795c6cba908673d4698a25918d739608f5de275e396e095baa331778663c1209c5fbe26b45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ee1ba0aa0ed00f4efd4defdf2b60bddde7f0ce7ec8c4ee7e15b56d37f7f4af22902bd2d7d79d48e700d8b35df58c9c89c332fb69a03ee94a26dd9f5ccfe366328cf68d27e9c4bc69dd6e3c63e16b80f2764f8e596dc0c85ae4e00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d46cfe7d71a06eb1db84a33e8c946aca5cec0716a3249f97864a20354526a5f32398284b82f3a1a4727d9bd9c4fd1b80ac96a6a19899a353dfad6d55d51e865f3e8ba38a4959a8434418c2d53d4b016feb94edcc5fba657aadb48;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebeefd22c78962b4bf2ddded672bda3e751162a68000a4a76177415de26c6992bc45c51af1856441cf1da68c3f8171522e42133dc70e15d6d9fb02dea44c5448dc4c9745662f9f05bd9d7dd5742d1e62d71dde556489908f63bd6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bce4810c3b3f528d11cc8624688482c3b0dfd2a79d022e575ff869f2d20e0a17e9069565367d98f9a46e82b7eeec90c83af45192d8fd5f0a8b9085412702b7ee9f80cd7f3351b98ce38b342a9a75bc4b3cd079b4a3387002bdc7e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4672ab6cc6e555e304fde31df449e8bf3c2d3b62fb32f9c9819790a3017c409c94a0187421f73fe645f40f1c047428e5528d12463a655dda0fc862cfc8ab5b3cba27a3cd9bc3f51b5e041715b3be6eb54ee927ebe525172393f0a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf0d15f60d64af3f11a5d04f266d9179d45e6cd490e6267aa56c6b38969792cdb220bc1d17657a1b56deac63c15d32486f70ca4736e5375e23ba8e90abf4a758a25498d1612a59239470a22343b32c517532eb60b65f2277ef5cc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64ccdc968015facc976891c73d866dab0de2d641080d2bc95f3158e5d3d18e145c471db8a2ff6663d153f71a51bbc00c27deafe7fdd2a26376263e608386046b801c0c0fc2b1e738bb08f9d94299c29a2fe680d324aff89a254b51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h506525e3550fe3fbd9b5472065942ac16d9cac161912803529a47607f96f47bfdaf486d6035c82f309a7b1967210e4e789e14335c855ce1d473e4e1dc130729de34954940ff0733e3e3722335f63bbed5820e0e70a9efa76d052ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d503c0b0333e1879ee7e1da5ddcfb5969dda6150a5c39baa47ee832e892fa8ef7cc5d06fd5a15d893c59c5eb78f59ba78867d7143a4f55afba6a145782d6300d5953e1d8770c3e202f8b3c75f388250fd4f1aa81035945d215815;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd708fb69ff91d9586a8cdb2c3fab3972368c62cb3ca0ef3c147e190a6fcb6eb93104240da0075e4bebfe3e56b4cc76fad0879efbb4cb00a2a4c956356430c1d61332121d951060e65581a53ce53b7250346ebf2406a8a0694ce8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d090f3dbc880a32ceca124e6819d145326f2a1c1ee686bfd5afc151a2c64a099236ad5098252ce976b87ed87f535427301dc9fc75185d89aece1f5b6d7a81cf4d57e96d3af9bd527050f08588baec427553814c401a6901df54d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132d2dd900743757a322ff1c0ee57f7be71a6ac998a5fa2de618b5952ed784933803eb03cc274977f57bd8a87d9abc083914675df3f4677a44ce80a26cc7ca3ce565c8a0c212d510d63d6c57dd3a1920b5c76a1d2d15fc29bba934f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1927703236542e3ad25da7a4338c5e16392b1125e9631296a1e4230a9388d7e73f2a20510a6933774a6c3ededaf06e67f8da9384954f10ff3fc7213e9472691a134324aa8ae312605f837d2fe29753c6e922373b36ac51df76741d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a12785cb14ee8b2d6492b724fc4a17353a46429762a0debe962f6805c8832ae2c743cb15394b444dc1a362871aca794b246c670b3c5d43a1bd7c734bdbbe2359b18d65f108a3c70d189920ffdeef38950ec1d1abf364af04d0971;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23da454853e52ffe3826d8f998a1e12eb234e7c49ec79079925a63a3ed96a5a1c3d9549ea43e2afb258c42d39ce3330b11e7f4fa8f19bc595b15be65ec5dc1457b73bd047723d2fd6f5ba7f86b9f4c37716588947536e36284299;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1874a117fbdae7f9880e9f2a74ee3f7b9574c004b361c5f7ec8edb2ca6ad8ddfeee86570d67296cb58d5d931364548ad38415b744d81b106a4737c99bfe4286026ddfc988241117abf1c9d7499af12e758bfa1e4f7a69a5b0a67117;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1611ef97706b3b1739881b37ca5eff123c81e60793e3b2e67ca647ccb4bd2b2a20c8b3a67969333a62cfeda6c3a3643acc3fe643d62389abbcdcb6f7ab8d27c0edded0efe5d04ccc8889039db31bbc53194da379d919462dc181f5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f16e385ffc073baf7b0c3cc1aca5f0acfbb30ee6e43b1c4a61dd714f384ab0343308853e6c75f228c27d5426a1a8a000abf530ba11ab2781f57830bae1dcab40b625187fb1ebfd5dd9636be371be5312c535f4199f243806be502;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127f383c9c52060d881c7657cda75a58ae03ef545fdfcc7a3b83bbb11a026d2e91d8cc15ef0a539c4df1046a069f883a4a623a766d9f41f715624a685cbe5ee1a2b0bb9eab01f9e53487ba38df0b73e0af93ecec4fd512136dd6b47;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ddfa6c4f9c99911a9326dabc289fe1ea9600ea6292f03f9caa632baaf2817a8bb683c01b3b7d93477eba12a48f59784095c9ca1855501a95b513d430ab42975833f4ebda941e28b126b9dcc769eaf33b6dc44cce083c84fddd606;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31f45584e344472861d124a4b601d0833c8dc96415a154ba3186fe05a31265220e133bb3022940f73b25291b788eb3cb5524ddd4202a3fcd5fa87dceaa71725b0583de78bc9550a33b35d3bd984638450ed14f8ca5eeb5a0530871;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb6916e96c7031b949d6bab8ee2e571d77a5ac808301b3d29f78ac9f7d09ac6b6f98951055535cf576e53da204651732448488aa398473b596a654d13911a2c822e8cb472c53bcf05cca998c36377074f2dc3b85a330aa51696650;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ab19d7412c7314832bee3a325fc7924e163f6ec9cf671c5ea1d80d1d2156288f83066525024127a202ffecf95c6d36f9c567359a34b497741e8dcc3b5b849409fd2c09308b8fcecb03d4e189407fa84428812a3ab47226af0e064;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14855db19fbb33874b36705e863f80e3995042760a888fe6bbb7a598be466b1a2beacc6e947eb613ab6d21cdcb09743320f0075ec3fb8d37704a68c54e7720e3a6f0d4d87c935463c7bfa45fe8a9f243dbea98e5b71d44de8a3b108;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e95d75e3ee599e1cb751b4c8304fba76bceba872f16bd0406f9b0d9eddfe8194b94ffe869cd7aa697e1a9c425bec6f2e1422cae0971611e33b0bfa0f5daab780e4ab699c9aa205ad4f34bbe7c730a2e865c514014261da0bea717;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eccf85b28c621b4742e247f8072130d715581c66aa8d9f16da15b061b8a5d288432328fd52ea944ceb6219d0d6a78bfa16338a3e1b3907913836271a63c1f8775a0b653f446a5fc9ca3d750ec3a759ccd1921090efd25b35e04e70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e164c6ce32d24c0d6c3e211f5b6440f94b6bc830e8f948109fcbb9a0e6b83b5624a12139f92fddce3880af74d786b55d77c122a4b1077cc7d62226250eb9b420061a4b67084e9640c491b8b98b3a9e5395609121588c5a4833da4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e06eb9f4e5bf2fae6854f57a9632f47a0521d3baa9f966cee945aafce59456c0ed593d9c3ac22da5e8b73ca2d8ce8954eed16d692f87b5d05577c8e2398b4387caaae9d05558c1609fe2e35c4bbe4854f62a7e29c1d2ab6dfcc2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14df20abc7ade45ddc1606bf779e6e72936293c0b9a31dd51d1e6389d708d61713188beaf91aebee879db9122f859cd674f6e83112ee2998db268d8faee5d4b3aed38d93194441a89f87a2e16d5d5ee25f6316aecf12124f16d30aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf00deaeab41c7876b44000fe0f04c71de44623abc90f2dcfa67ceb3b00aee82d59c7756cc73fe7f495664c797bb8cb4ffd0263672a74623c8f81a7bb12c27b334ea42bda879651138cba16af10d04bd52f023c2f7146cb948db83;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf7ee603f39a8e2ececcd1a0c86be513fd5aa0fd8ae3a16af8fdda43d09a8766527fd3c4f0d564d76a9962ae64b5a76acc2f7f29eccc0beb6d0e3d5ab634361091c792c946a4c62d8d574be5eab97bccd20930fe4bc9328c0517c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155d4d0a3ca8be692e40a6470513e79caa5c0148937ae414ec13e73d84f743071ba5b945c1c4e1c53e9de6ace461d6cc54d0766a76a247c79a626420b6ee3bcf94f23bba0bdf1853abac02a3a2284ba4ea8b604ec8172373496c04d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf223f50e29263760e84da42f99a93b4bd6c8510bea05a35dcb952eb5040e634204bcc86162eb1cbecbae670638d898b13d6cd74f349592053383566fb756140cf0440e1621cc082af0d68f7c97245caa8a11181f3d5642d2ad774e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d53b0b6adca13739c7da6ae1aa7a385ede8bf2d9e337d8f3c2f88eb032f7a7c401ab8d494a548c00cd12bc0575f9684744bc1591b799a56d208fedf1bd91dd5440b9c23aedb5ad7ce748064e66ed4fb246fa7ad075a406889a2a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b9e945120f19ba9746c392bf4b4924bec24b6361613488f6175e58b82ec6ffc0a7f01da6aade19bdbdbbbd89ab91d5e3461fc8f0c20c0b6973f5b2409635f0d75f96bd7ba2a1622f25a63975087235fcd2a0dba1b757dde57e48d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb561447283b1d9967d0d29d27fd6dc5a0a33fbb785f98c80bb49b5d17eb90232d24a8ae1ff1462e57e075b6779ae04fc40e28847f7d0f59fdab1f5af95becd19f9eb5732a4ab7c339d47f4e500175afe310d5c39fa2554ab6eeb3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e496b5de9f551cd918d559939c4180440ffe111578d145c9da687e40409ff4f28b493bd3d66242961594e0831f2d93b2930b53b929911ecff3b8319c0c5250524decc37d057e9909609ab2efa65ede065b45739980d081a5b0110d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14192ebe1687858f5264138178a50014d8d494080e9a616cd621040ec65830c4ccc9c789c8297d9ecf3957d8c5d4718c8258e8207b23e9f349596cd43a5dd6f60c2f9814dd9aab6944c80f8d0773a914ac299d83da0673b4d4024e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcf1859aefccbcdf3f83141fadbf1a712511ebd865735b58d97a7e0e8b5e78aeefc9e481816825efa0df07bda39739682c0514701eefa0af66ed369f54c6bfe0654805cbd763bb5b2e9dfa6a28b33109452a276ee4944650300db1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d82a43665515aea557e4e43c6de93c938428e811ecbe8deedb24775ed13ae06033d3de6464e3d26a88ae3464b908520f669f897ca7d2b4f6e2c7e76072974323876c76287fcceba549f9e6cfa19f0d2fa6b5b79e76dbbb88cacf6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3d81fc89414905b2b6f4f3a89e41a0404cbd0d50c725df3c22997a1eb69513adcc701a559ca6e7624d19aa9a5056300db3fab0a63ffbffd800bd8285daeb26b692d4cd99d8112c78aed1ce43edb1b9cd30e915e5dc7319414832b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e111b1fa2d521acdad021263d37c9f642a6896c47acb12db741bbb088f2bcc85db0e7b66274c173c0873948e5fd303d22b9f3950140c1079d1b2f827788ec67f7298ecc9099f95f13dd9129eb3f3ccfeec3909a022e8c679aaae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139ecb74676e955a28460bbe7ac2653baaa272941920f30bc768134a3122c4ca1bf35edc927791404b1114fe863d0d0d71c87b9f91e7c70997e01a0795db583715a1ffbec82bd149343e9c866f0ce9e55b91329763066c3be5a6388;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f263f1313d0de7c94d08949d29fccd85ae0965f12d84c6a0484c81354cfee77250e29c4f0ae980d4af40cfb2a8b123d3e34310420abfa825a4c36e88fbd77d6955148e3536786fb8a58a606ee4b5ec5090068b92561a7b351e09e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b354341f3564e5f9c863d74bd8084ca6c49b6d5c43420aedf35fb44c4c811f762ac9c053b350c2c85b23d2d8bf93dc13f868dc534e13165d25bcb46f7e10771b52812c5e3f322cc37c598a9bc62d296e19d8ce3e41bc3123fef9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3bad60064d8275ee6ccc3ad6b360d23e30ee3c48c098f1ae658c757ac572be71cc78948a0d6deacd3ba8f852e3bb3c87af0613cbcdf4214664c55d787d0ea64b5f26e1433f0c1fbf65867c27bc53d6a51649d418077ad7df77705;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h527fa8b852331fcb004b7bc72dd5db7aaa389d686e3e968df8ea6f8543d503830716d3426e5e47c96c27b2fa7847b2e0b1777d36c376cd3afec3640da3d1afde4edea5914107e36c7a5b0997732953e694c11069105f2b5fa1df23;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a817630f1b35db5adf06ef8190c92782d1e402b0ff863325bbd1673fbeca4dbbb29779c27abe65d25e7a59bf56d74fe13c39c73c63eb88835e2adedc894d991d1a9bc89ac163b919c13bdadd881f7a8aee0349e3b80cc07fa56b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f0bac3577a834e24e900f42ac96c1c4e8cbed723a44f4735a78a01c83957c964485977f321b09bb5b2488604e65d5dd2ec13165ca35fe7f02199d90f322f3fe4e3f3877e68c15ce6847a9983e8582ccea8d865eb61bd2554aac1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he85661475303b5020542372fd4f616c34b954b7c0ba390c27002b2989b1ffb8cb7c13af3e5ecf77016e1eccf7bfca0db85297a81aa3980b38aa7ce95e1d632ed31e40e56a2c1c0d48854d9cfade9c527d62c149646bf52537c4649;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16aa41cc2b6b0179165da5820b9fea9b640c385bf45673a2898d875a27eee92637ad6889b23dffedd4b61924db9a5ec2b53c000fb90ed40e25d326ca9ddd1604a1ab7ef7d7008e38d73bc4dddf7f86fcd138b218894e83425d0942b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114beb94390e9139999285e4ec8772721a202e5cadb34ae235e367b1f89437b85d617e491a9a70740ffaf5066f627e589301b6e33a30d3fd96aaaf4d6e762ab8171215b66ac6b07b16eb93350cba2f46ceefe704935c18b7b32cbbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3122759faf802c2205f08aa7ca836a877689cb9a84eb7fb7c43a0388175a381720e690c3c9c92eb78deeb1a912cbdfbf11d2a709bde4e0b5813020d0b7b6b370aac23ed3864000b8e683a15aca6f1af91a1fed4ca3633a3c860cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c8f7c1fc4be629d46de82560d7ec56600432fc26dfe7ebb31cdaa64bbb5d58b4c2e41e85668208ad4040a14eb4735a51be003b143fd4c6dc5e66edf96de3361758fbb08c1bb9377e36f5de1675b75ab554df749c3864226ad308b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91ac6db580e2bcb9afabca5a9aad7a88318275e5a999880e6e1239567e9e88433a59e936d3eb1fe3899e92f9ab7ad383ffcc230d0155ac5bff2042e5e555a80184f99a96f5b25cfc94b577f0a3228f5371078e0ebb8dcc9bd91dda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc101ebaddbf416eb3049c245e8a0eaad2d9f0eabaeb230fc46061d5e80275bc88ae5071d1fdd01cbd26166db61e4dc00187ff6635b184389c38549aa28197f8e831392824f66eb41046ab0330cc9be760a5d3d507af05b14f4bf26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156e3204b3148e7ae24091f18f8e2e475b1974f2ea46c9d13555bab3963155341091b4135957162f52dfef485dc166e37091189569a5310de67ddc3fc2b5983fb4879a825b21612cf8f65c9957561b57b22c01e86d5a64b28c3b7b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a50b330404820b0f61ef9a828eb1425fccf888b1507022e3844719bf48fc9ddaa02e9cfa72b2ae57400d0980a4369ce4eaabf1736b5d8b998c75f3d643d35de1fc4b9b201edadd25a0d5552845d30191b4940c014cd056f41e1d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4961731f9722af83d735e3b713cab7c124a61092c470d7dc45cf007fa1d25c2b98b2963b4592baad9c28ed5c71f0aded8e3fc89bddc72d4e4029f61009241822aaa36f9d1240dca01be6187d824de829495671cd80d054c3f9c80;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hded80f3903a14fab2105f8f4a857a6d492fc986feae1c5552180f0ad850f2afd02d46f162fd30b628fb180526abbad2f5781f0caa64e3a0076a8071453fea3eb05d1a2d4da6e84f735462f612894969b975c2c916d4c7f42441d06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1290da4bc7f5ee9e1d46e67d52151d69ac5296d57063777d7b3736584af6c885ca556b9c851ff056df3aacca4de7851c4f83ff3bd4349e49243690054997d0e95bf9190b2656b0df99ed0a5e9ffe669afd5e2bda03cb65523434adb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143a9fa86edb07ca7347e9f120e5357e8cfd486ab201de3d1cf5581efe87623ea07ca3ab95901f60432c5e6c7a3179cc10521a2f83d74a9fb9735af4db2f5552bfe83dc7898eb8f99b182016bdc1f44a8657bcbf26e2ba4519eea2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fc86a164902733db5de8accc19a9dd13cb2c0a45f89eff6d9da8cc9094628757949e0ce77880c804bef338683055f1172bd4a5443c715f65bdaf4fc2bd2949f8981d4d9429be8f73537f2416ca8fd068d0c4a001167a85acd0e5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h225aaba05b6a2f9c79a8872dc6687b6801cb674a97d053eabe0ce01f40a305d81fb4d925546aef832c10464d5d46b76cd0b4dc1e700d5248a4c50e914f4f17d7c3a96d02d1356f4dbd1fbd25ef1c166f13e02abb77421a3cfd5914;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125fe895fdf5b209fb03513b91d82ac3b92e1aec86bd0212c77741541d77a5a6453f893b11977e72aa0f34fb9479c4b6e53f6ed9a75692096b131a5dbdecb00ac23dc8a04d4ad38cb109b45be32cf3ed951cc8c3f7b189c0b86fa4a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4f64f8126b1805a85150248f7a51dbbc306919e3da7ecc9ac8c868b16c47c6c27ef8df555d7d85fc23d9b0b98d16bed38fd08b991609175f0cc720b293d0abbe9b31c5bb57974d616d14c80c4ee37b4c6964d1881bab8cb6ad438;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d52f2b41fb869b99d43ec67a8c67642a600f8e9f2da79da3688b68bc42959447429817c39a20bd7cc851266ef4baaee7d798a82652063fba5a4b4c378d170f5cb1e8a6ef80d0169accc1bcd3afae2de36f53f9d2df728bf640cbd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4e52ef50f33bbd2f1b5e7ee3779f1946f78236be5921a0cf5006b77f90b4cb82d8abc5f81489bf8501365141fd84573032e00a956824994b2b96867640d3200d0b1007d7b01331d0c7a070ca30fe0c82551d4656ab60a4d1aa069;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5337c33c7fcf3a0a5675dcef02655bd1fe8a1bd675632be0b0e6ff51f760e0317fc5db94e27f0ff940c1f2293d2cfebe5ea14a449843d53cc769a6c00f0ce7c2a3c15bf19db7d15b4e67faaa82aa69e90144db7d02cf7e3209df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h976a2ab7977dead1cd5c739374bb7f17e95f9d8599f43ce4ba47187ddfb012f55ad0e727cfd38268232d9a3eee0b46f72a3987e172b3c7cb0682a72056db768c68056eaf6f060e40dbd0377115f91174d11c08e32ed37e21d9ad9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108d929c1b9ca1bb2c8278139e25deb1839004869ac5bb92281ba672b94acf073b7f1ef1276d7dc332f8036ddff0490b211761b158f6cfba906b08e0e77f1715c404cd54df5d2a3beb971cbf7b76369d420e9e0d839b3b4675a3720;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f56a035a381763062576294018be111f1054abfd2828eae15be7e714389523e6492df2ad34276f3de701695c27566abce5f1ab99ad2b5508d48f7df9fde1f7e830c6f68cd675e1ac1b82908433c92a70e3747e52ce2230e1eec86a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ddec0993ac4898a5f5269ec1209c3726887b01fcb3413e8286d519b327f28785eeeea391cf6ada29d44e699252d9ac449667ed94144334f25a79daf0df6f356ba28d57f3a048a44b9ff99aef48e76e89898940b977724f2d8faae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c32c10d09ec42b8f331db18d8857868c8b89d982c529f0ba298ac10695a497152e3f207a826e5ea56a61c2ba70629e75455ab9286dff6caf44ccc8f0af002e068e3e049b813e76e6d2dcfb6f2373c3f5970e02f3447e1a884c12ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183c2b1bfd138388e0801e4e236e6034050b2ae8fada8bf6765c6469ea5c01234d31208fbf87583f2c9efa8a4bc02f827188894d79208e83e6ee6bd0d2c07b0af83c0db00a39943a32e48a0fb3d7f734c7a54321aed50d6d86dade4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f4bf488dc5497fc30e9cc33c771c74d67533a319a06962fde2dbe5c28caef8b0c4ac6e25bdcc543bb1fde9004a0bc79c7464964b2873950cd32c0f57439f1bf836bd8f85eec9c4c6c1848b4536cde1bc2b07b56cc8e42c6feff06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h725280f8a0656233d460bbf12b3b44eab88b0deb4ee8acec974f894ca7b0d43f6d0150627d854e02af8dfa2cc241d847feb3d7a44a187714e07fe74df62cd56aa4df1eb32b9d98ac823f3575720a59e2dad1b187cff0c5dd8e3f01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11343acf6cf2c867c07a9f255a4a62f7ad129553a77c759bbc9b37c7eb1a8f59ac679a413ff4143df5bddfe0518301cd043aba69845aad0023d93f3431095573735034ac5298164e7544ac9c685ac6d5c462aaed153dfdddbb932aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27cabac6924a5759a70cf6342ddde98e6a542823d268e8e543f7a6dfc7a9988a9d946f091c3b0b0dadd6378baa703f08e7687eca089fcad3001d9a28d0c718917d3fc87466282abe1f9f2d373fbdb4f44d256d15b290ff7a239c79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65c336e07da70109b7b8520d546d870034c5cfc2d7661e75cf6cd5325e91c4142546d2c899da9ea9a4f1e6b20f956ff04816579271da1c51a677a8cc004beae74e86d98a79480e3f1d16daa655a6d36b5915c845564f5d704374b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7f7cedf8336ef7353250c7895f44245c8584181ea691ef9c3af8bae9ca6b837b04a2c0856bae61be6f7dfd5999216b86e89cd95f9791ab3245a1bb9b56d6c51c32150b2f00c3d38e2733f5aca341fed7100f32bd0a15386d189da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc6180e727e05c56d018c3b008cc06f91bc2c25c0a9430a1eae53b52ab103c72de9027a7bd0bc6ef8ac1f8a7ecc00f44e43a409e9c5f461b8fe0235546c482b7269c0e9d60d6c765fbb5425df8b9e67a997e6817070d8ba0663065;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16522262b21377af5a525d91b73807b1c536bf21df2f52b786e3ce0ea8b5bb7d7ca3288b0fd7e128c2d5b020a3e8b7f5bfb9ce3b66b1f89ebf1f34e5f411c33f6ca0fb07fb3f1f6a87b208c31e92d21753c8d6b627475a47f3e6869;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17bcc7169e705a2d86c9c8d5743057f2828ad80117cc33bfaddb82696b96bede2de39fb171b49e10026a46bf3f13418f8f6d98538126b487488fd416a53c88090aa492776df2da25ef053ce6cd5c681b0b92e2a1bfa2783e8554a44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bb5215df3638fa01b727263ae022702d5e0f928a04458cf80862e8feffeb9d87a53087c72ad55899cb88ffe5081002495f365554219b68da62dcf82d8c8aeb6f4e5b8a45f329b048d3d494e332c142a761931dc84169524ef2205;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef4b1511202f94b7920bb62b1fc6b45e247ad3871bbc7b1cbe9004266493bb2676a18055ec39066373b45fc08a295ce4dfd6b77a1ae93293b28457b043751f0c278f90d300402b06062445843fb991c0359aa6d1a3d8460bdb9df4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe8d525f2a52c13ba67b13137a4ee4abafab62b793a1f1325a5648ce95257bfd5bccdec0e438ae9e5f078b6c6bd14b63100e80e211bdbe4125f2eb2c43091e0d8d6480fca0bfec0b527c40202cc4510ba0117cb5ba076dedd55b9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153ed12c12c3d14595503bea8939318596ebd5b145583d0947b0de7ecacffafe56d087be5653dc0117c9d69c865ff16ff92ba04c314df5ebabe108210c517926a399b5652007ac5848eddfd96bc82f97381ac5e3c62e90ba24171ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12dd8d4e75ce09e8c6c8075a25141d4e24a73c278e2beffdb6e69d9ccc7b7b26e9f9472bdb7f358ad13e1f9a70e51a6bca60bce926427dc1318bc7755257570a0021ffbac9d1f6a97f8d2a5864e8e3aa4c3b171dd2cf4582ef87ab4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had2254a6204faba6f3057ff0f95e6cf1c4c3f9a2524d587a1aae4605042f2e2392a3f5e160f67f7ccbf7d129aee01047f31760a5a272e81d18e606d46a329413a102a213e07f0f08f01855db63e41336e13a99481d014937bbedbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h363da0cdaec298ba5652ebc2b937caa1e042504bb0cdcbd65fd7d7cd17a241546e53f695038f51797f06b3dcb271704b81ab6966e0af1a329a128732054d46ca0fa7507363e3da81d1ab688f50316088c9ff3bc8bed6ac0e447314;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136051951e01f7c06ec2f02ff71e6edf1cade0d499f1cba009b0dc94b15d4ee14b51118e03f36a1e183839594621f693e77d788f3eae360fe33f423946c39baaf6717fa6b5fa3d8c60f7f611012d4f5a959df7fcd8cec39ca9d9346;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5bbf71c82afab90d957a0cd623ec238af12fffeaacdda2df0941cdf47b08c8b708c955bd0fc9d56f266e87452b207531c4a3f999adb825752d76d5ce05521044769fa3f4cd60c30d8d228cdc02c94a714f0a5e9d7600054b3d04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6737299f19c715dd1da8c91d4031b39577ae46fe64322d3237b1790d020562dfedef2157770efd4dd6b6b645472de0b719ddbbc46cf57bd1606bb21ffe9d48a0a179f0f27b19de21c88f2e03a89f0c9918e0d5b6bb558c504b497d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf1cac342701188e5ec5860351fecbf5f72ddd1cf95274b4903af96248a952721beaaf1bf0a0aa576c611f7ceba962dda25bcc6818b533f5362bcb308b29ca9cda89cfc3e9a8cb7b390fc89374d7fceaf9b569f8126ba2017814721;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cbbddc5ae2a06d464c3b054517276e47c9a582c9fd2ec7122ea8bd918b2c85bf54b2ebaae3d84f9aecdfaeeb76258908c6ca8bad7e20192600f37515be126334ca651cf41348790e1171e74399f714b40b5bfb1dbc92a7edb1873;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12daa48237fe9e4f59d1abbb5cf08d0d6d4776c9700ef521bfb8c3fee730b9c779a0ac8e0dd5f564405c4b79b8f204c57d726778ad49fbcf30f1ed0d1650868ff335e6ee4bcc7bf40f1689f706447ff4cf013aa7d3fda5573046f39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2300012333b05d148c71a638cad2de7475d71e910a3726e797dcdde132aefd88c0f3b6b72bc797ee4ce9b27c90890758f82a56fe80ec1f3ca8aa89503b7e7c4304a242f08f7fe6c5d8eeb11bf6601d03b8a425bf201ae33570ab98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63a33a7ab482bead39d246468d327a50e6ce6e5faad6739f170bd99b881cc10089f7b1aa0f829a5ebd20aff81020382954655bc7e18ef85a2733fd5cf28b288b7b148a157a58d2158fdbcdce5e20b0f64acc86a237a372a144f11f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bdb0a6875c24dc434ab7aff28227e068ee43dea088c6bda9da4de5a76d1e79147b7f44b4885b4479980991c1ecf35fdc662b56d1db926dbde93bdb84a059a0a39aa24ecebae658c9f53debf9618a7de24bec6ceac65e5fc5b2ae6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171768c42133356d722f21bff3225f476a8f10c147f10c093263b431d8a08f53041d6aa6ba19f30f7329e175a9936b54957a1fc5eb016c7bd42f4bdc8bb4f1dda4e0c9e6d69866fb62b85ea9bd4634a6ddee789304433400779e7ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e907b4434eb8b5d864a1e3266ff94063cd86fd6b354345fa97c66810d6a18d481bdca328a898c235fa1d5245f1640c123483ff604ecf617886ca9c1959ceeaad72d683aca42b4b50df2d42f0b2bc194732117ec32e11d5ade1869;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h481a8629e09bbc62df8d43432c7d7c4b4314e6dc50f960a90b14404034377c205a99c3f37bebf246e7cd7d58d5f4ee02d68759ab8486e636b953f510480a51a6877fd16c6912185c71559ab8c5a953eede8bcb1bba247028e89cd1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had1ff16d564a5307976fcf855575fcb10362cd97d414e14ed96b5df30308f42979cfbb118a652c1348d0ea27d71be0a7369f0d6a39d0a1d792b482740003dd32ad69bf2968463691fc46d14fb18bb14088dce64a8a5119dd642249;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1682cd278856e2e2b58864a9e7207658b7e6e0c4a1ec29c0a655f42badc014bb8f606b552220e70d43031284062ba4005bc01e63b33e4023d746873a197e5e33620038e53efd082bfff7be53f23e5c569d22a0d8978317d8e2e71f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b820c2a85a05067a1ddbba3bbb843d4116346a3569ba117ad9d4f4dc1d5d67267f25513df92f1414ef43b841a371254cc455ec890813f5fe2ed308223317d9cc44af43227722cdee2724749e2a321152c247556cceedcbf26ec33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a2c47576fab101ff3818dfa0e3124d8ec3e09bdefb8440eb925d05cd883135525508feda5136c06cdca5823062666b05e8616af314b56d30644ea4a68a1f23494ac0ce121fb36bd5a83fadf60260355a195c6aae819efaba01239;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf5122dbac86ae503b3eb740b8f4dc882aae65a13013c13fb974f5d7fbafec4376b1dcf65c83d89a083a70a035569d28702211de4e2e706d53d45374de0fef2cb2f538190851557a8ccd322940d5693093e2866d7b353a5b010972;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd81a78fe4696fdfa3f4989df56515e1b8d0f4bcf3ac1a57162e96c8eb767d247c354f348989a64cf9be7e00f13792b9444f65a963d63f9417be28283a988944e160c221006cdb1f0942fa829d663d556638f25cb7d3f1555875f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17646402023cd1f3a69ed031f094ca602cc1b1dee1a0194cbfee82fce6fca56dd55dac66916636d4b77cced4b85247a35794bb162be6f7a69011090dc41c1f27595f2f1768a533a734efb2235ef719abcbcecbdba8a8982d6814f6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1513ce69fdf537440b0572fd298d7f71fed1741f391dd3b652c3418a720e7a07ab4367b12315da662b7328673ebccf661bfb0a8dfca46918e43e5cac6377aeaa08547c3de3e63f8489c62c07b1839f50a6856be6166d4a340aed584;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1d1f33ef5c6d7da9260ddc0214911c801b178566f17b13bb0e7bdd7b445edb334ffa74c14f0a1f35b3aea607c03e260303f27d3af8f878b2b602c7cbc4560cd13a9af2c9674c91844b6f2dc2c0a88294eeedecfde1eaf802acf13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6e22e0d18bca03f9561db8d0a46f3ca1bacd686637305e9e784e49914c5c8d3be23c80571152dbbbdeb539a84dac3cd07f3a00beeac7785a01521e3fa7e496f2598ec77dde35233d33cb6a35e1065bb0fadfebdeb266e93f6ef12;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10164e2fe8907847b35116edfbba3fd00c03b7ba771b489b5216c9f5c1bce2ce26550ce00ede4b5031e1d334541efd38ad3c9a6425535924006d3df3fe3cb7fc426164b3bdb0d22914409a30d528e4a2aab20e81f565b36d9b6164f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b11d5b4628b4075042f00a37505b5b7c07214a3f29f27816a72e1bfb7e59ba70fef7cba18535d6c8dac6a8e30567d41723c70f0b5eca54fb3459f964c975f46193e9c4d3d6bcd79f6afcca8e3aadeafb9dec6c4f18efe499731ca3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5cddfa4730b205585d37b73202ebba35a80288c0507c80414ac8f26842e36e21867344969e90b1260bd2e565b424e85ce338dbf35e8dded3ebd971f90b05554ce0d41938fd13a9ec1a2282413ce1263f530d9d3ae823a1e8eb6be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8073d0ca205e7ddbc2a198063b284d734ca43ee4a7624d21c4dbec6e1c3bf32649075f063696c1cdaeb8929fc5a70ff81399cd834e43921ab14acb6554d546f483ca16add9fc62737ebcdf338d6df4a06cf7ceab31edabdc7edbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85432e458c213677dbb47b1c4cbe7f65c403fc371d474aab403b07c20673b1d8ea2dfeaacc71fc99feb8b2d9095fcf128e75cba3cd7ae4eeeb6773a2db85c5c29f779e954f5c5ecc315c3975572d5d5431dfa9edfa648e45fcea4b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10989087fd4ebd85d63cae838aa4e25d2bf34b3edd0c4a25798e6e9daa9d658725f06b6bc687505384165836ce04dcd9f42cf709e6c70204f7e28ef6cccd9fc3ce26d4eee17286baa37d26379fd06cdf543369b1fc685d43f67b8a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0926a3bb7c6ef23ae78a530e5ab29673835f6aa33b62612066eb76a9086168ce79e6eff30d89777db7c80049f3a498bf059750cefd0bd5e256bd68f0767b13bb41ff71e666993d86731493f894437a55e9e8f7ac13f57c4b04021;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144ad0a907ef1ce13ca5ac3cfafb6c3c4f2272ae904c7222a4405542cf8fcac51e3fdba64ea41204b14eb503293ea73877f59407292674b0344bbbf6d63f46edcffb437ee58d0e113991130263df75c9ecd8afc19b3c45d0cfe784d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94fec194a89c0a119c71fc900b42a08cb3ab5ca5e1575c390f9af529fd40b3107ef49c67ebab19fae36cb65007c9697bbf8e0774592554a7119456366cb7d8b495550e1de092daf543610f4c29589354bc4d3f81f5ec2776fe104e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1607643f175f81dc912b687870c7b9c934b537cd4fc7ce6b695b167d2b7dc2d52a63d1063a2d77eebfe725027632ad696af93705700588a9e77f715b7392a95d3e97980d9f28f9943c42b824f0c1b97d3dc34808d08730c5fbf0731;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f06b56d304bcde5346ee169eb65b0b5e869ac0f518d1d50a9b6a8bcddb1952883ac0d0b4f2fc0b3655838544614104499aee778f2abde3b1bf6540d66df8be7bd3196da20426a50d92069f0b2e0dd4abb91637c1dc22850ba7ae57;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd434b4f59f37e71e89a6c198871326bd5a2715211f4b0f87c27dd27cd90d15ad18ffb6677fef4af7d42ff6cb6e78bfb9f2032b682c93f00164dfdf50422926496927bc4158ad1235d34fd781fdfe8fbd87c298362b4c57d67b9439;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1225c7b3fbf5edafbaf2d9269cbe92583dc071bc78ef2e0e775ac81849e4f8804f77fe4e43c95097f8a2af4471c89709eb2d96fd3e64a525d2d8a144c3a0a502310cdb2a1ff8c514d0bf39ff544eca9ed6e2a8f59b0a7abcade2fc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab62e12084e4abee0b2a1d997dfc735b8bd24a3dd8b3b526ee62d1e4df83024443039e6f84d79db7686b46624d60d55441973c08eb567263bf3b1d2147f87ce4f5e18fb69c7667879080f005880eb4a149827becf52c4b8f402f95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be3d12f1fe6e97ef479a2aabf993400624fcbe3a5abfd90ddcc99fa00d83c8b2ff2f5315a408eecbae2223d6aeda26de679a3dd2448d5763662f73628e073ed062234ac86bf52acca9882e7991859fa020ad99049c42debcd870a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdbce4af792d0d872761fc6fab8b7d7e3a148870f31c92082d6d8b43545b1686f3b9e32de457ba0e3add52cc7c7740f94520df7698bc490e314807ab27ba5b0c600a50d469e6ec3be2b7f3469b94b83f93468bd227cdb3826ced7c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4743c818eb474da33b8907e3279a8b4ecf2f76b6a6dac1c8e54467445745f7b9e78923174b861c76c33b6cc1b64315b7e379488218251d79c744ac52a9975104582e21a59050e93bbbaecaf33246021a35534ed4a6af26aa2595d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad08eeb5673edc7acd5bc86303083f3e91cd2f16721a9edc34b5ccff239ca609d5fcbc4f9910ce487570b95ad02bfe96a89487a9051b71f37a30752b07c47d241f466b25203420df3ffdaca77ac8a970de6c5945970bb8e5b2ef1f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12db8ebd385206206a73af8750809ffe67a3f66f34806018dcc3f1f69ab491fbd7959c632996c6af496800c5d8b902674692311d2afd1d37a5471cf219fc6481b24ddf33eeb1712b77e220574c9c146856507c16612c1ce2bdc8d33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb87f41df6c485669a90ed1f7415b114024488a2e1fdd8ace2866e597246ead4f594edbaece6e33cee85648d0ebb4f1521889b10efbcc90587bd005c83de60e1c73008ac71b29c98543ba6e3118fbbeeb3ce066c2180b60ab451be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99c049859e6638efd30d8aeb137efe4fc712a9cc154043d56e9155ade03df41e7f832ef9f544695f15d07433f5963091d963e52977f2f9dbdb02bdd2a88103a1cb7edbebdb3ce71174db9c416bd492d15ae319b5418581f2436010;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc228232f98b226e7b67e8bc87a6211ef9baa5b9ee1ea48450be757dd0956c5155d07decd6c175ba5e353356f85bb9585888bb2becf1f8eb5e34c84150befdc739ddc4fda959499da3a6c4e914a94773adbd5a5b649fdc2b51b858;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba2eea42716c599f18e09db61bb4ea0e9bb8389e463b839d14ff14570a4d20fc3319239d4a39f8ad052ef74c1e2785aa8c62a53ceb58e6a18739523a86fb7060adecfb08cb846db4f9d63ee0eab4a6a03736503266069943b0acab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8b77118c418037c0564a6e4f35ed29d36e2f987e5097f664da24ad86602c0e7f63811387c164b3a2c467c0588170bc1aedd75de0488cd74094548a7cd6d0ef0e61feb5050ea591997754c03cff2456f3f4af6dc130c73ee9feca6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1019d104d593a49cba0ff541ab9ac960deceb17db09649a112826195a916ecb9af04dc50f2159920f4c7a0c110f3ba485e315f00d2ed11d635e997fcac2d61593c02f4a79cf82cba92d6187a4f170c98ec41afefb1a553bd4f5e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h765c20d177643158436265fbdbe4f259addbc0c5aad0a61e0cfb8fcfa1a5cce7214deb78748d00e01fd4dd40c52b4246d46127b1b55b816c38d599e38d259726ced58b94b4a2f818d1f45356f52fa011cd5b49afa17ae7680c5fc5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f85bd0407240b5fc5956bc03b552877792bfcaa330609e1d60a358c711a488f4660c8104248932116ea4f0c3212b6dca392ed5f489e02a5eb22c39c0561d95bf3a40ea5212c87278481daba34d37eaee40bd02b36787e48973bf9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84b09ad3eadaa61eac792d1aa2f7790d767ba80ad9b7ddcb8eb5f3745acbef9997d519b03ec555f0ccb4e9ef3369ea541218b1fae7cdb3bf4c8c1dfe254cdd7acfc1a0be33fc546709fdeccbfb5d798c13caaa6d72e397161c5330;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcdf3cf5c0717f7b6de1a48405934e00242919bba9708262f3f53d6d133df4b4f1c08868184331d7114b6a6fc12ac315d645e8d1ffd5969bcf41512193121d779708f3e902adce6e63e568cc308d46d033996c05d1273eb08b32e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12598a47576dca06d06ff41268a333a0c76ae8d8dd753f51dd2fe5ee4157a16d18da316b8141e8c2b19d75941044db97467a2a63ebab23b3e3b47bbe14eaedfe9c76f7b26c1bcac2dd397f6338e8a9102482a71e7e9fd9ad68524a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121e6d3f99aeeb65cdccccf3c989606bb0d2a70e4c62d1ebbbb2e786e557fa3570f0bc3768cb95928ed4f5c7d4dace94937a16508b67b98ea001aecf8f24838c4a0a0437bf299fd862a2c5a9f4105d42b6716d9051b83331eac81f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h421bb8d8c6ba013b6f80d847706415513214bb3eef6a6ef0ba2046ec5e47b8511d118373543334a45d40f18a93290be5757fb9082aecdd839ebe48728f7aad57d1fef91f01ed160104f9f51a1fc290e6d9f9eeea48fdc5dc8c17ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fdc214ac513ae87bba56bb0e8992c105e4b334539ebea896b34fdd4646c2546b6ea639b40531e62527944c2c7e8b52a69b5ddfe7520da7c23430eda630f8c3bb3ad1cf3ad287f45954c00f7d088bde38b376c6cdc01c0f692096f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f88f04db1b754f8cdd4ca77b9aa20142f63d061f821541e668461e531bdf78582b49c78e1c6fc06fa7126994f41ce4bb3c20e82cde2ea9de0f99ff0353b75afda1e09203fa1884bf94acc1f7dfcc22ee9bdfcaf93d6b31dfd496d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h582bd8649fc149be73b571157f49ba12a4a6b24e01ed305f53ab72d2e11f41ba2047fa882c7d30359c6f1749685f12088a1041bebd9b92d3ef880035b6ec493e87d3ecbab9e8dc741b6401d86b1460117e549d7057e12b02578f39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1c03b5e0373a2ba3973b8c37a03d6740293858f94d08729ba2798e7df081ce9abfbc53893519dcf5f111141a29e357ef4871fca2006bc02dcc9cc57cb0dafd5e24b236471ad1164d1c4b3b4ba12c8acab6a9551bb86a89ae39ce6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd8c0563b824e8c7e04f0e1798dc89e4a4de1aa5430209729691f3b857130d0e0fe8fc052af8469d18f4452dd9ec86f7b373854456f1b1fbd90c7176909bf54432a974345baf7caee4c116149bbee0f6244681e99e364176ec68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad02da482b6178abc7b97ae5e16069391f243f33703ccd1ac781c5e080e51309ff64a3ef92446ed1ec23a3c262d8733de4c284e77444869f9ebbb981e9846782c3666c5e28e28c18fd4871d9525c605f854d24e60bb9c82d629ef2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc94ecaeb9b070638fa6898a7ed3d818b552393fa2c1e0c555a6f24cdae1ff75c9987ec9b0e67e20958f201fbeae012188e89722ac1b821f17e96f330a3897e59e660f1cdb6ae49be4f0d2158b2588bfe229ded6d0a33ac4ed2170;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d1ac80d656626530c4c05a42f98d47d631b5f4d4c40147450143d4b7796478672aea9142108ba4831ba578205ac523c7f99b80b25229c224da0222773c8986809c6e2563c5e04f4dcf46764e0f0ece9451dcd6147fced88854797;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h400b97e416f922ea92ffe98b7fa750d97dab14cfe642ed3865513915abe0cca6c153c4dd7ad3555d6051a11e3ffb436a2549388bab2996a45afc94890802c05652dcda4bd81bd08e16b227fd9247070b3a350dc8582f025044df40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18781fd3aac3a7a0af0ab89e936b027788951870906c06a6ab7ceb438a67a586f4dfb9221e9c9f9187e85d1f1c158f7e1fc73e8f446984c04348ee6ff51f520bdffb8a2b6c2732318bdf9e4fe295fdaff3c6da9c799ba0601031dd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7eb5822358fe95db2011c39ba6341fec1631eb350038b644762d3f242f3cfe0e80351509dbe4a7bc8fa7d8f8ec86de05dfca511acdb47af710cd74f385f17ca4990f641a458f41eb40bf1f09dc5fb5a861bd44296572ca301941;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb806b664fbb6a2438dfe4cf13a5e68125864bbad841e70d0f943726eb420d159e4e1a396d1e2c66ec0753bd2f179cf8b2a0402baf10373f51c28870b04a60e1a009e784389b3d67b4f9ccb548e7d9dcd599b38d3efe702cbdaabb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h428222726bb60939caf7c57aea5ff5b3d42b937461f051bccf3d401ea114a18e42df27af4b28ba1bd837e18cf32b4376fc20dfe35258adbb16d6cdf771b7b84fa9fb6bb209c4f500a6740a218bc79d928aac68254e974fecd9449a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hddd9a2c2ab1eb37cc67c166e9fb313cefc671df0083ea7336be02c5662d1f7282759dc722dba3c96fb674a7195fcc7c6cc617977605bd0e5df0ad71c26217a5adc7d20be9d27f809c02800052e768d47d881c0daa4fe31f014bdd1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1886a01d62dfec1b381a7a998893f9624dc8e7b4f0fda2777c5676e234a7323ad516c869a233e6f8124fa66d3ef1b4d831d8493f82d374104a8e608244ee62913a39c45a1f5225aaecf8305ffe5e5a4ee962c30ff547b47d1589643;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d8e8d9c435d6c7019559db5b94f64a0098371c98dd391740db6d886ec7c1a7031f5db2823a1bc04623c3e30f13ea64fda0ecb5cf9aa4cfe715ec73b32ef627bc45e0157ac1778f401110286c4a4e8d3eee2fd5ef48efbcc22c86b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb13c13ca5ce616d8b5d8651f4f38d923012f00ac813410a0a944e3f9f8152e9ab8af38844981e3fc1a9a846ce049bfc9e82e8c0b6cb7a3ca491e54c76d7661925032a0dbe2e51e21e2dd1a5cd8c1fef973d3615b5746f593aaa0f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1260e41991691849a47318e579a178f646384f468921da5a5ceeb438154d9e3c0963ba23e916b1954caad0b65f4fd5d0acea346e409e1acb32b2b775f7547f3d4bd7d45157260f68a4f881c28e70143af37edffe2b583c6e033722a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d74ab1b371e333dc31dacb4b57f9fd8e3662e18fbf3ae9735ae5e1fd0ee94f7c6e62d08a04509d9c757a7c3f9b8e77e38f6eda848d70c608a2123be0248aae2104a6e3e7d051d806f8af5e2c79d56d9ca5b7c6061beadbf5fd6c15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7669b13f9e745709794f134dfb7f21d1d74e09c5409ed7debc5a1bed5470fb608465a8e7938dcd7f2408b0c73bf0d0fe518e61709ebc157017106610f75273b854f645ea2c7e08357ac4bbfdb5d32bec4784a7c3de5f4776f84ac0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7fa98c51a014ecf2fb1bc3d03532af505be39bd08e0344148f7701bf594579007c8a4bd9d090a67afc3d888c9b4478198d0902c26861845abfe4376da75ca32737cbd5e8c358327d97d6ca2313f59aeacbbee9713061a879111c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca1d5dabcd65157261f602534e8ddaa55769db9b35f656399f5493909eb01d1f4e0123b181be6ea891df0b204ac7957ae5e3cde7e6dc2228e00cabcb2b668ca550a99385f99589d32e6ef6f1b136cf63d44701ff0fccec75f47ae5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115bc08194644c47bc78e0c23c34f766fc35a54f579c5887b87eac187528f6061bb2bff7a4b1e47a843ccc5dfc0d714a7d36fe4529b75205b7ad16dd2b9abde8753a2fa74fbe485d9b62de3d7cf38be0f88e9c38f5bd1a39abc530d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcb9bb8c393b0a12c8b351a66c83207bcdb7c7ab0f59d5d3e648017bfed4313544621fe798f1a2e5db1d32495c2aa7c69a4c8b782b6ba0f0c52d0b009499921004e173a5541304202e4d8a50cbc42d10cb103120bfdd4e974d2880;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb83fb9b8dcfc6a85251ef69f5e8cbc8121a7d4fc89905d27f2d1c3d23b83b416feb131e42c46202ccc3d2e4de6041583ef8c440b0ba8cf1e91d563d1e6a4a63b72222d797bab896a71b969cf58b64ed4e6a816cd7a64249b211a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6f59421e266e64e7c3f253926b3e3161979e492b18529be046dd6ac737598e26dd4fa2dece73a16b90452b128273a60abe615c1bc70d093d30b6adfd959e535114b7a785af63b472f6532308e4ab7af248386cab3d8bc56f72c2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f8c0c62df333cd9c7780fdc27857f20965bbc10cc605c3ea6236898041c10feedbbf978953a00ee590429f8916db85a05a9e4c4629e7e3709c748778cb54ffac6709fe02447cd3600e367fe179e44fdc4ff2c3713b1393d7e483f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc158a75551c4e4433e1e2f394ecf192c6bdd65092466803ab1b07454ca030517c4fe415cd59e3755fcec4dde310ee4fa0922711af714873501d28bc8f63a49d0ae57182c523aa52f40f054808fdaaeb7e34d9c612ef3e37a9e26d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f23af4aa072a61a2b54f1862ccf907e3d3073d98cc79b5fea7076d8150ab460b3da5aebe91f55c908159ab2e06bb992edc6b6b368eb7014cd82d009e53cc3d974d66dc9f3985e0ca3566111b2fd11f97e232c7654d04b0363ad859;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e656e3dc47b0e9797bb8f93f148b74840ba9f9ec50775caeaf9230740c095a7181a31a17f75ae843f4ef074af7d3d68b9917af3538e4745fff66b4b7d6a26ec4a7d593853ed573234ad494d029009621182352a5b5e200a391d057;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a793622fb6e1b6520af3dc325671d7a0931d603122b9ec5cc9015516ff5ec039a80d5a2c6cec434bc11c8751c6a4895b35447d6e8c75b1e5344a1516cdd90de29a45ab47ed0c8ffdba366f54c7dd9e10e44f62453d283a5760ed68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd35e1c3865b3168175830ff14072d6fe67af03ea161bada2dff67b7872e9524f7a0a46595908911e152f2d3485592496122dbcadc5ed594e70276ed2f246928e96995999fd4091eb0156daa8b42c3c5be7e31ba4d3bc388d21a3a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca8de9eb75edaef7fc913d874fac974659338b6d67b52bf3aaf55683899f10ab9082e05d200ad2ae4c046217152ad25951036a18a6939a3649e22f510bf342636cec88847ed821c7f52068c4fd3e3815a5a2bcd66651edd9c231ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd134de35bc503ac9f0457feaddee01b66192b06e838015aea20f47b724f91de632b906975b2aa0c4840eb9910d664d09b122e3aaad0d75866d90604e341dbd1932606bcca86ab3af0c3872c537762315ae97f7cbb403b7450cde7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196c520f00aab616c7e5a08c4a3c85e442b01388b2a4829903903bac22a15cf9473391e8032b64a22d801e120b7aaee8fe4beddb4f38726fdfc0d7572d1cab7faa74b9ce57c24c30a92d0ae24e4e5961ac2acf8726ec8939f3f395a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196c4fcb754b9baa2d3e89cc9e80533e6af7bff3a92f943cf680f85237994ea8f6e09254aaf0a8354c53b40fd13d09b96c5b95a5650360bf79fb8d108ad58ef3a0d8c2f7774b05f38255720d41445295bc4b43961e3f69a4d79348c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174e8f1e4a66704684361034f4ca60e9d207829309b2846e77ea34ec2f455054a96eb653e27629599105d34da97940fd646fe7eee8045513736857e9ac96162200c7c0286a02faba4f6258959826072575b26d610ec5ff70d7c6a7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a636bec0b4a4ac53d5b91ecbca2ccf6c08eca24264371c1b7dd2f2b15d0ca05916d13b46274b9a7c44d4e5950aa5df14616a969a1d3fe53ff627a428be82ced9be988e3d86ebfbdbdb14baf2178df66a35be12237c0d61c34c06f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be61fae44b5a8cce1a3c07ec9b4349915028db3f862ddf630adb2e613f5ae586b80e64e6058e5b117975d90651737c2699bb84eda2875849d15251a0a92371afe62b9e7bdb0fb2637987a6fe1e4394602f9e0545ff4351f83aecf1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf63189d2cb16c9264d1d68e5133d39be1a5085186be0e9c69bc27ef8a7f87c381ac9f8faed1319f984e5a56a4660bb04ea737e2c393c45d41f52c890d7390fc46cdb0f00d4ac4c6b523c6be710a6bcf062446ab3658d128a99878f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174f9346b3a007406bcf6baf5de9ec1f10524c64221ca94ca5aaa5aabfdfa42f1717fd0453543b629105ce1de8d895e0ff075dc02161202bea4563a441afed7cba021d646749981bb9505c3d2f35c071ae3e87b3e43eb47b5c252ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19850d2207170caaa330fd0be26830e72e85830ae02f71f1fa2a8b85ace88f90d30fbfc30fe35a5ee0993da6042513b0b880fcd6cfe075af1cc657c27aa46f9217b4f787959adf00e2546bc65abc7f30ef5e50a8e6a8fe228265bd7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170554af3a9ecbfffb28dca89fb366b8d91df356d9b86f649ccaf96d462feb2d711662fce251f6d2f34d998b2c10277c4b5261f754ea73e27caaea0baa4b1b0e6bca28ba03786bb774508cdc22ccbd75a42e9f594418ebb36dfc76b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h890916c344d2890960b9916234b77f25611919e5e711cc598f4166e11a909e06b35db9e98f244416422fdd4b573375d9cd223701e38fcf19ab39e424977ad64800e98bb3699307c6ae39605839671dacf3c3b1e2ca8cad2d80a2c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0f265dfb74e26e6a5d922d68a96e56312486a65d1712fd3dd18e5746578d84b3e073d76017beab9eb58fde27acf313e661413f1c468e8746a3e07c595c9a87626afc5add3134ef2bbfa42f24335253323b1bb00b30c8c0a257f92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbee21673e96eea098391601b808182dc3e78008b8d8227bd3dca8081c585e69c3ed788705a914dff144054a91c19bbd2c1cf2ce18f55ae54a7824437e65c6a324dae582590affd0672c4fa74736ee07960f0beafa0f57c490b30ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d4e23f9ec19b5376c9063d0f0db6d7de7ea77a70491500d28a91a3cd1a814e3617a656f469159d26dc68134f902dc3196c9d9988d5600d20a48fda9b984fb6471105e3952f3442c46f84570e297b147c416a0727c7c827f38648c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb884b35ed1e1f9586ec1bb664cbfead3e250d7d9cb447603c15b26c8176cccfb5f5a326a99cc5b97e7d17467b20ef9995c6019b88a3ea9bd7ca9a1d93f21439eaaf5adea1a74408809329ee7f41a609a4ec40f905acba4a326985;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7d7784e0ebeb023d49157737d18b306d83aae54d5d8e95c419c92062568414a8406943039c55d15359ced52d71243c59821ed8e5c8beede85cb5494cbf96fc9d4a1ab64b2b1c89a547bcf398725050b3cd8c64474cc6348ef5c60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e6652898842059564fc9b4cb3e2060bb45134c8e01ac8fe76095ed4231acfd3605e98e5542c129b28f0cf34d694e44140b5aef2650db8875fcdd8dfafc2c1cf72621758830dbeeb88d1142f2e65dab2973a16b9f81c7136afe038;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27404f554ef476189110b529f45dfadd70c1cc3b0ad9ffad8639daf4894999a09e1035d118434bf82da28f78f639b857cacfda746a7db53fad78e482b2e69b7423a8f26e3f07cd882aee3f74914f411cbb87168596cf598fe06f4b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h579e7d543e55eb17f20f06bedabd8bc7c88d41afed65cf6c6e78d7bf002a2933b1492252cedba97090125043ad1051c46125f32107541d631ca53539b57b5d1a407a971b37853c12c31e06cbb6a6aaac55ecf4b736126f7c1f86f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1657de88f0317e20435068abad8001ddf68815c65e99f1d0525a03b42aaee7785551cc0920a8b5d75b45dfdc113b83fc266bdd0793b8b023a25a80293b53140fee5140b4d83c12aff17e13d5ee90c4d9ae2b500dd37cce945cc85d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13866a7071b3da117fd6c4c9fc322af7ce074a7678aa9d7dd00336d2a72c5e26347944f79e8f54587a38c23db17c60c75a769b9136fbecef3c8aa2c64bc19d021c89c3a2956c37d57643d621d800c267eeaeff06c0e250e08df2f58;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3924347814bac13e5f08fa88fa42ff0bc494b4f20f85bfd04a589fa0f2b797a6319aae501298edbc3492c09d581c5fcb5d8a3f9d99b19a90c44b006b186d48de1cc6aa0cd4dae1343db5c737b843b7e38f92394aa8a906577e481d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab74c434a60d4209d6f26b23f31b0de414d94daeea6db2b4424108198b38a5673bad9447f2aa9833e06bd0f07709d15f7a7143f0562a28e78cba5c6f4ae4251b52238e57af5184c09037f879415c2f5ebdc1459cc6f58fc4448b3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dea4550a8908a88b561f134bc83ce2babfd253bfb9a52d6fdb2b6f6631dc643a1b56f7c043b0fcf5aa646253e690bc50ae684880e1265c560d2208c09e828c304a548e4634552e50c9a9a50c194cde273e1328f4e205f323490d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ea1c6e6acc790856cdaf4415532cba09d7f7116b7868cfb4e9e3b71ee3bf482ebb253816ee03b5e20c7b70fe45da24cc870abdaf982f674bac2c8b2e82607ed9de703ae3329a834e81a83f5ac114c16c3612e6a83fcb64d28c7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53fe3919b9af4cfc2fb6df48dbc5fbcad022d69a4879422e316c4326411cd5ae1bb207397d46f1f769b7b9d5f2a898fb8f63f9908274cc7dbf5e62f9405f55e999909ab475e776ccf179e5df6c27c4c22f1fa2b3cd56ad23dd5723;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h486171f51923abdb83192270c0b212839cbdfbab5ce82b3aa675c33d7439aa659a9f131630b394e7c54cf2991f5a9f0c42b0d921d7820129dd71f1fa1ace38b2cc1d3b5d906b65af885d2165a96ee90f0ad524098d6df47d73ef2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15653415fe817c4b5e048d9f72e7074e8b65e32f4331db58608bd17531b49987c78396c811285912fda276c58d68cbe650eefff4a1389d8de7a83c70a0c50bd42a1ab1657070f5d7b67e8e4aa770d322cd96b96dd934eaa1eb5c716;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd0cdc4d2cd88da40e0a84de9b205a60bc21c9a74a97b5b596875100bbe97bde254d2df7113697d86da51ada1854297c815417498c6a449e9b3a90e4b0d7ddb2a5cdc8fbfad7f27dd9c25a7c222d9d862f80aa48b0e70ad22a798;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h871c3b75fed2d8e29982a3a86f878cfe3e0663b77f26c63c04b62b7db527e1506a081a883685089210dc79e2207545cf7001cdd047d359ab61f7aca53d7d767a650fad31b6f39e98bcda80f0a4a246fbd465de7f2ea8da12b0e34e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd3450fe882c9cd92dd43da445d2eac9c9a5d834198ae88255d158bda6541531700eca21f6f290941a4750e1e618968bae891b19b5f4eb928b2f5749d8e07dc90a617364ba37d228f64931e8f585b78d9fb3cb3d397a15c96bf2e65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f58869ea71d3cb253381749d0d49ddde02a8c2ec1159dcf178ed870d8100671b91f53fe0288edc3ea951b29f5af068dc0af033cc7c0737e1bcdccd6ce95285e18047bd81f5bc862b9bdd1c3dc342016c470acc8102c8266af77fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f43b2d172e6617e0e7e5762bb47c7181a26a92ac5c65a019a060241eca261c7b48a39c04146cd1c6daa82516bfb0fd630dda2812d04f9b8aef5f2faf55e829b01d3d58916648f053901a1fda2aad95d7fe5edd486eb7d5316a110;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32a2adb261fd65a2e1f74bbf2b3571b57a3ee4d37871613156546b651a775690758281781e5f11c786dc6bb05870f30059e5ebe9d890028b6e01e2ebf5f9559772ea99adca2bafde898ec35bf21192e2ac4f9b342fab2aa1ef45cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6be6bc610fbb4f28ec3a9b9b78ec13a7df382bd691d369c2b1c28b3c58dc38da00e6efed1a0d7d955dd159fe5c133c11b597e34cebd8b1b374e7b39edda27bc6cedc233e9d598953b6936f16d1e0e35ad6119038183b38da00c1f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3577c2baec995b70829be66d8ede9e9065eaa9b9f9a3acb99041b63059e33a520b35b981dbb533d89c6ff5135c5923daf21e167ffcf8f4ed53061a5a41689d957a5d7bb80c132f91c22c23c38c1e2a4e703d900e2af0ea451fc4aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94481abeb7ef8e28985a9cbbd34b3ed54b13aecd0e6f3aefd9993659a37d4e7f0dc46727a469bbcb99420f7d32b41dc530e3a791924f957166a4c74c1ec15564201eae14e79c14b36d1424552c1d7a210aee95f2954efd176515e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a9d8c60a2488a8ccd823f01121f2ce162bc3736f1176a22a14fa0b74fb6f7224630561a6e1666c68511e85afe4a7b1d5619d7431887fec46061b1f7a9e642843bfbfa075479f34c3ed95bf360b489a3e44bed5d6d87be8b1c799e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5cd27fd3fcad25aee8f1dfc859390ae8a9a8581fd31ab985168cf3be58d40b6e2dccbd68fc274ea8df29ca8c1d93d2e4fa3229178f3769c9dde065586a57503554b76bf8d71fb2d07213c4c9a57837d21db373cb56cfe8527a2a45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23c277694986dd06a811bffd323750347925095fb7130561afe10e093fa7cca538339ae5d6e0ecc74bafa472dff58e081089e80dfcb9fd3d3601f92ad46b31088003b422dc6dceb16807d2e2dd52c162bfce6e980e395f861fe5aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cc551f2c8b460d14707db5c27d0c3f4c603f798fc12acbcf682efa34e01c302e8d4c631b5741f12f9b55b18e1d04d1084362db4b03216ecd880b28051aa183ebcd003357313a92992b9d1d32bfdb9a55b479c4f8016b80f839168;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b20b020fe84684ebbb2756a619c7b44e30f2a006a13d1edca80718ef4c4184292444def74d0bb57206e3bd1765045b41537a367681bb86c6b7b3dd8c35327abf5bcd5e532db9d3d6d2292144760791c190582319470c6c6bd2eb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h800af0e1f3d10ea411ed8fd271d211f54f459c40ab259f676d90cb41c74efc568bec97d4be6c858a81a86a775e59a1283f65b0c33a22090e398d92f9098e81135f544b8b763101188fea25e78276ce0372f4aa42de99b5068e93f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1f89000cfc33f4d63353374130de4a988a2e88b5e580dcd2b76ca4c434feed46ca428e34c56e4c7c23535901b8426bcc1de99bea5b42be0544e05e602bfbd5a2466c6017b1fb0f646c86d2f97b46916fc7131a9722bed00d9b8fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h887bb4e9c6796ca41e2800f54080fd257958494ecb39ef13bfc42bf92223dc1beccd33fe61f2e24c251f16d5e4591be2fe3eb074b21700f35280aef5b2161508500f342efa8d8ad177898a5b256f7df0b3774697e054f7d7201cfc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2f7d99d1b8817bef28eb9b7997937e543b38952bfbc24d810c9d9e03dd3efa59529cc8c9d834a165185ad20c711c5e48846ffbdce0f2401449bd03768b3444e14f5abd31399c37b2ca37835051ab14da0686ae3bb6ad876f2b5c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37d2adf861679e9fb1283a651c44f51b2374c4c538c8f1d748aea50bb1fc4656a2913b82b13e5414e03add463df95c0e195879d0ae814ceec47c03aa357eeb74659c1d2e8db2c5599df1835274c34d882dea5e96298602b9914729;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha426ab964340c47ba55b3a281f0306d9f755fd5b1070e90dedf066db6f421b74ba7472338146e564228d171caa038afa1b47df00927e7f66f79110a51cc88c1f366bdc9e242d75a75233a1c8416380312e0717f61f191a6d35d4e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42d6b1ba2d1dc5015cae75e0fae989a7ff5ed197402bf70032a3575625f24c85bb4fe795a373afce52ee51fe9251b8c98275c8eacf8ed23cc2c3dc08c2e4d487f5ab98bd2536aaa36aba6be84f4c738aadc2feeff3ab2c19b774f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8095ff7a30a57c07efe5efdeb3331cb8cadac569112584b7cd58f737af18d9ddbce43100e04e1eb273cc023b1428a5e08c988301bb4ca380d8a353116c67820b045a40e3ab43dfc0d37013761a7ef03f050ae5027d7f35db160a35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2db6c65569b012aedc6601678a49d702bb4650363cb9e5b9b006e62efdabb9f51c9526657d114af6585d9e245f30ac2d684f37ab817fe7dcf1279fcfab8cbf76b426a2d36dea701ac57bac0333ff64ec4a3ae3e45bd910ccf967dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b23aaeaf17b8911869c42c9f91a281666df9ce006fffb1af3b5c2df3d2b9dcb62c2e2f0d3de531f3bbb3b0c09cc6273b596dfeaf97d3602bf1d6cc3e04f927c91de6e93ba929d3d58c8b3c2afebd47447fbac4a6520ec5f528ba1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5350e1024af0b51a05662c17bd9f2fa36e40157c1ff7ad41f67304571f51bf149c5d99668e9c396346290d462384058975ff93a64e8d744b60f062caf64e99521b249811406e0db1073d17d9e13744400d8090d0111709d3cbfe6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23d86c53bfc2131bb08fdb54847e681079966a128c11f85ec1bcc669e40c098efa11684bb0378b59247a8f723be3865669b614b4297d13e0ff3a492b0de1a02ad66074748c0df75bcca59417fa3f4370ea2acb037ff2b53d4252fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5bafc3dd7f463ddd327c0474a14e72ed3c6ba45b78acdc82af4c129450caf18169141476b4163c96f76e7eb3172d4eb488e38331538d3306480220d155a030d9a392b96f4cf9118d12f7bb487bb1175c39cd161513e9f4add1359;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e0bcb2fb8110e636d0eb2b1bda20f97bc0e65e2f0d4b013997c9033839239cad32ddb1afabe7b040eca120835e325efc4e0effef0b0004b6092ceb5991854524fd017ff339ab9957cf86f82a4b3a989b75961065472d34121c1b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14db3129c5d9ca089decdbc99ddd99802d92e961ff5cb35c9af8e7e48666ece80d19fd81f337bd0b8b2821868d950565011a6db0929b12083f481edf833b8bd930a738467ef5e760cc3a58a9b1df029bbac086f3bfb59757c53f3f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf46218d0bc0530d7295c31d034aa3bd65941700684753defdc1eca7b50980cc61c2e6d3015df63873d988f1d6938329cfaddbab0aa114539a617e7be5d73846f7451a1b04f0433aea9cb56998a46d843d5a60910c1aa15dfabee7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caefe82d368c0a4954da7ad39b81ef0d8870dc9441966c49a29844eff088628bd6e8f26881400bd4cbb519f2bbe1ceee221d02b07ec3180a3d843ce8cf99f308d390410c39e5e249f00e5657d9df1cefa34978326b7836f360b7d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbc012097850fa847c08e068c3ab0662cba3e817327e8aa3b2abeaef5157ab577994f236032b043c0c727a0a8a24ab60ad1c120ce379e7b36482ca61f8680d3a030ee25ab6c19384ab9e104823127c6efe8d353922edd83eeaad8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6109ab977e3d33911a0791cf196d6684f661d9a128fb7fcf13ed0798abd26c0f4d2556fa3dca5dea99e903bf13dcb1c9ac584ba6c4cce32faeaa683a3c7c0960c91a1d73b6ff1d99492074aad0cbc48ef213e8fb45399fbc16ae06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd73d0d2655b2d929e13cd7273029cba9e1da863ee0742ed292e7a203b6fb962860cf0ce490bfb9cd4cf07fe30aa8dcaebc5f2fe1e448ae48b1d994388b7bb02ef847680267da309c910636a480e603831126a037775d91c1aebb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187a3225a7d321ac2ad1c204af813d71ad0f8155e5de5cf2c18562a8e3505a2912f14d9aa8aafe63cf19bf98d5064855914309d13b01d349b9621e44854ef5aa5a8a63b80e29aebbf3fb3327761b0af3383148afcfd93c139d94112;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9b78f8d188cd498317451fa0934d778e076dedd72c3c158fa5b994e4153aa30c6a28e99b596717f4e4516342497c6a932b9960dd72981fb2be5b7fa5295a8b8fc6b0927470e2ee03812cf7f55b4ae410ea374d0e9fe64db79036f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41b6f456470f4f6f8850518a03eb9abcb344658dc5be5928b34e2e4c6022a9133a58a5d2029f06ee5fad24db828feecde6783fecdfc0f8fd4de040c9e5244fa460fc6436416b0b58ca396d6b964e267ea1052f055fe7545ea2f327;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5cb1caf7699a7c648a62bca6d33e87c4d22646c91efd56f2935e38d76cab5ef12035a16b3477e9dc52bfb11f94b0c5d49c4df457a516ecf7edc4cc5b8bb2be34bdcb24cc037f538b70cb217ad7b424ed16ac88317c4e45c5cbbee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ae7b27b0e306b8265d8fa09b255719629b7aa38ee3e6eebe01946f715f0e8a0deb2468aea46610cd99245b96a683af069c8c364a57d87d656b19f9eb3dfa930d9ff1a1946134f9fbcb871daed023f6d574d29b8477f6e39bb1153;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa30b4167f73f268e91ded23e1baf93cd8ea58f5db9187d4c972e7536f79a9c23c4dc62f809c970174f6bc3ecd6a0e943b5d0b80bee414db7e1c6708adc2dd152cbc85909ab6dd3131c8c01509c8f0430c2732762deeeef79750b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8ce62af5447bc871f8b668d8ff08cb01df3c876611ab8d01c46d1f749ad3435347146116ee4473770e75cf6db8c11eecb7f3710645fc4fc0402f3a6c538a6180de006a2c6280e302c164fb7329cd1e9116e26f71efc6e7ad43a41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78340bc582c8dc0460689d54b59aae99b6a040455df7cbb1ed25f176753652535bc5de00638b928b3f1884fc6de6c79aea75cc7767192e35770d3342ca383d46ac59dc2a4a9da384d12932a1525214150a0f49584336481d3baac9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h477524bb99629219d440c89db8742d3bc189262254189f6ace9c8bea5bbdf263f87636c994cfaea913b7a905231349f70cef7789fe2b3e8975c0f8ae8c236638f37ac21bc6bc0754e4629f11165cc1c67127031f5bccec80d6cea0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1552b4f8106f45fd28d9b5d50ffff9b70da9571b41593d8ec9ef74dc51a76f668747eb8ba9843bfde63882edb40468e3012dcd94ec1428a2da7b7b02ca29fb434d806239d1eb1a4679fcb0fde4ab0f6087d63708379f950bff6cae9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3163912f25fec3c54979f6f0e6d3c270445c999c6bd658702d3e487b92697e79858c22f3d151ce05ad8ca51dd81f851c01c33595437eaf4ea1c28a63b0369ea099bba6e434f32d6025aad0da20106a523bb21ac200a21ced04667;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4029d9349c9b91f64b2f38029e816808dd755d8b267f6b8c911364ec2d5e782c58c35410c5b9fad2acb90abea562902b93ad32bb44eb6353f3f8574a501b43b53c2016107a0a90ba773151c62e6046211e2fa090045f40ddca2cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d527081b637d75d849313bf035b8925ebd523f9b40983f19dd9f4f3615a68b6a17cd6b12f77e67673fae68f04b52380c95909dbf4685eb83f70f19e25025dd7df386951732490fd68c493928bfd33ea1d6ff1100ed361601c2bcc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ba2e6b8147ad858bddb0ca7e6ae235f1f97a77bad2e889218be80947026fb685f08fb972dc672e2df4513f33b4c8811edbeed0c42bef9a0787e93e7ab3230bb9f1f1908a4e457d835c3aebd9fc92b27584e9871e865db16fe16f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h680a1be3d6c72f5f78aa550f1e7c8ca584730f726dbf58bb427da4294a789057cf462182227c627ef8aff266801235e5f8441bf83a15633c276295c7b2a335ffbdafc3a9dd09a6daa7f357bf51f812914793d598083ba51f5f0346;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176515f7642c0c03e364c6c4ad9bdb08d7e3353599ccf53e7393791c5f10037adf89bbf3340e1a77e17b05809a6ff02dfca7f024a4bae5344cafd9be9718f5f0e7b5721a0859d3d058abe3e2933f646b561e316dad8826f650fc7a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17119b74826ab141619a46143d482a8a719eb07b760cfbf0fc5b8e96aa0eb55f574948314fae2a91405a73664333e81186669697a6fdeed4fb321d9cf99ed6435799b95ddda19ead6c8d886a2945ac8a8a1fdbdbff7428d739ab21b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129bde6c0f6d11524de5f97e0254e1f6d00eee67b7928be5fdfd217d5585ce7997409cdc1afd4fc4526de761798786d022806228e9c9ca698927b6894dfe995f466a607706a09fb8a66d863df21a4910418d1ae2e917a5f4d269c14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b396e381d968b40a9539e7d71830beeb79b3b4b468f60c317d0e1a113eec2997c66361238c2f0d075d8b3affee3e762e1144ae304601f342a1648c34533970937aebe2819a13759753d98ed51448da5a8c4fbbed716c8bed89863;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb91326f88f71cc6faaa064684360497d077a9042ec19bf516cee4c016bf0367fe8827cadb6fdcccb479044e09e60392dc0a4370d596b75ca225b35f474a053db610eb27743667d6bf434e2baa54e32476db5ef6aafd40eb94a6f67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h741f6bfb24e996431855abc60a691d2ebb90628bfffbea032d413b2288888f1e28be5b46b4770687e52556ff82bf2897481743ee584fbfa4cea68bec05e898ebc181a08e3d78f7f8d68f54343fb1c004e36cbfc423de45f717fbdd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9e6dde69f3d6031f88144ca14671cbe841519a75c9fc7cf8f83f1a765ca7ccee6f97552401623bebf402bd7a1060c348b4cf21ba763cf0b6865f49d9690e8b9b21fb979f697d9e5bc52ee0eea1535dc5896ce2b8ae3bfcca0ad79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13dc4ea14bacb9ae19c429421bbaf63517a3716a50ac75e9e9567d59a161f28a5f589e53153cb45eebc5b41f58e351435c6c7bda3ff4aa3abaf8a996dcdc1b1297c987a41932f13d353b1905c2228de472e4d5de74a99c97c9da574;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47f613c55808caa8cb5df259c0cf6997d193c7136607f8c92a79b0fc7906372b5c66611f272f575e694509f9078c82a2ed3c349f8dc03161e1b21be53ca69f655127512bd536332647239bac1d07e5d6a132d77838a69c997590cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdaa5187ab9fed4d828b6d13585e513889ceb85bd192b3b231a253b7edcfc4fd5fdeca91020bc6680cacc9bc3369429401d798e00d4420c9a634fe09272c069860bb951687ed7606923b90e0d5dff486a5748df6e33170ca27c6f35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f528f0138312369406e198addeb7d4371a1e4b6bc3e74e1125fa97245beaedd86040d42c3dbda81f8e31d92ca9c4440d8d2ddfde38a03de443069bb11d8f51842ab73a376552d871e83b1521baf6c291cc54b13d5a63f89f7e41d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1232377cbda1fba81a80c84662d4d25da433f4d2e9c1821b1e456ede71af2e4a231603dc5265a1027cb29a1eb2940bf7244069612075e69fdb44c8f7659cb73f3b158723bdd618835e5eb1675f33dbfe68f5e863588427b14d0c053;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efdb865d1ca1376e6c8aef1506aead6098508826b38bbc68691ffa62ac4ea724cbf24c227cc6e44104619ef5e36b6c6ba224b59ab4228657befa2d7164e7a76b74fa2a9a7babf796aca8a37dc6df15f80100f1d18234687a83eff6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd23d40cc7e0f0f9786d6f29a539b65f239051a0b56b9117a9b3a2d4b259cd6c4cac837a1f6f8d835ddc8dc03e457e0cb91d629b1b442a2919d22a8afc722d80d7337aeb054420eed0cd338f694b86b8a63a097681608eda4d523bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf93cb8fbcad5424e07770bd1f699969974d7d3ab4cdc68fa64125b7772c9238b72be77e9794fc026c6ec19c8355d3ed10c85cf740f0b63c8a1da0dea5d02e441a6c50b2d2526724ed1d945f5d3c20c60bf904ff10741dc675b6f56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7fb94beb4c24ca8f24e3d9a159e45d59a39a558cae03717881a3fcc710fb4418ac7f99da79c9edd54c006b8bd53ef4c0e8da500ee51edf4ea17ae15a1a3f5a77427ac02c45be957c5755198e77f69af3a68432aa95e924fb6f335e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbab2aa198c5c9f8f119a2ccaf05c340e47e104870c1aa1fc475a0052bb9288566a57594dcc6b35d0a18d4db2123592603851f0cdb45d2430fc2b9c814b4227649ad598e5a876779d86a87270f2fb4b066ec6fb6ddbf6864912fb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7bf255129b4ffdcc9c030c76038cd279ae4785f5e8a300f4437fcec31eb7c5e049d958a68ce142f29346e95787e32620010562f387282dd8b514d8abec2faa6ca4724865024a896bcc42b637e12efbbd7323285b24008ca619dc7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b172d85683301451e38918e7572a66cd15a44084bd6ac52591a68356f5a0662b63f362c855c005a9a0775d211eb76cebbae04be9a692017070c97e5c9f36a4578e3a59d0abfa91178c13943c92bed4d5617a7d2a35aaa5706ae5b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195c2499848e504c70d8159e1ac33011a19a066c61cba0c82403be01f3bc9d1d82a8791e7bab629a59e5965afb6ed28a9bb502491effa484c384c1863937bd059d6ec0ea9ae440110549821f94fee9c797842ab4f70c5a56025f451;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed838bfce5f1c379aece50fe3a4fe9322651ae8bc83f7aace37a381fb9ca2ae5c76a9a923c2f33ed8629a189fba740ab26dad3e92b7bad82d3e10a23f5a4b523c52e6da7d5a9e244fc0fc64d6aa8dcb5a2e6fb42cdf054705f5e6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1026ba8d18855e8a4c76fb687f27fa4790a627e4afd8866c30fb8f93449385c6aaa518faa322b1ae047e9c068066b069c1264d49f6302fafd042987c6ffc1f2894bfbd76588a083c58ef5da07a86e926d3e651b5ed7ccd84ab3bb46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d1ab06fc6dc5655c87835b3e93c7f7a03dedead28abe34df7602e0f1b30ce1e45d27f754f84202b8361503c8944516c677fb25b8cbed12deb0b6b51ebfc4bead293cd59ac08994ff9e535fc052abe3a5041a07462e34624721499;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1208069bb53c55d4421f1014aaad0c225f094db6fb2629720bef9df4c1bd93714b90133a9bcbea84446d870375e8786ec48ae9eb05e5b9e1cd7a3e6c43166ac9cebfdb3b0f52e140bbdd83d6aadf012bd7915543faf1ff8b5b5142a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd11782f37818b90cc3f767df24a3ee9b8b938a32e4004bac904c51c238d4af2d2fa53b915614734440920c1c261ef4600d9c3300941e0cb12bceaad18f634a8944963917524febebde380b24abf6fb4d4a74ddd5a09c9b536f28a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180b014276b156505c17ba5402172cc39ab319490b9b9acef3ce6cc8ae5ac65c159b86c8ab12c91ee3ab3c74d8657974dc51a2e650dfa5458734eb97b938e37c622705bbe8135ce920cf19e36858eb2ffd47493911a2b118c2e529;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61bffdb81fab7af6c3274e53ea4c96d3c6ab2e7b1b626ce6c6776377b826a5455a753ca89cd086f941802429bb5df2b030b03835f1ecf7f9a0e825d163bc47aeab9f7dfffe3c33eb1332e317e81a0226ed55f7aca5be8150701b25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h422490073c0ef2b830486e05e7c0da58df99acc42405b70da72b775e019f4a0b45b7b2b16bd037d223ba0c3eebed13ba65a84906b940404bcd5fd1b44e72567fec9a0370bf27d10ac986a893e6abee57f62fd8a6403f90e8021240;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3e293f361e6104d253a4d54db20205882544d55a56e5b814123a6bc6e0d50a111959751ca3cb36dfcc4f39ae5b22f36ddc86a3d08c50af2e6bd4e3f3863b8d1ace2c5129009045fe866a5873f678559b865f30e1278b89e07c2fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb1a9844d74b1e818048321d0be92f23a4bec29eefc97d8058ed39b22e31da93b4ae9506613bfc59c71cd19c4afb97e10f8d7c972c0b9cdda6a777f88a38c1af390ece9e99f8f3826337249aebfbdfd6264163f60a411275ad057f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a96f04c981576132e5300f6865e73f8db92d74b3ded9629449d67a0c72302b8860f8ba2a086bab396e6a8bae3cf37d385d4f2147ad76b53ede21b6120e8bcf55569974d09d91dfb172a666a6e3adc012ac9c2c0ed36bffd50822c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165b98d3c94759d49d34e2061b7f067c1939727c5565f2867d12fd814b2782f084b799879148e02b2fa5876cbee024d38cea880f6b5b0ffcbc93f2e7c2481ffe3646293ea9e182c430c62a0008258302b241a5c41cc8bff7a8dbb27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79333beb877261ebfe49bdb72e04f5af31de10ec11fbabd5306b3f3fea99b23c32b8051cf2ad10fb6e32320b8feb86c3d5b328669e3513ece1898c987ad736af603aefe62df8ef201f991216f0b20f49d4c32f508a7d3b674f5476;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c53c35d59b8d0b3d78edb4e449ec494c5c4dfbaabb1b1c8dafaaf7d34f4c95e39d2cc29298be88bc3817a9b88190ac87fcf3971e772da57647ca3c6445ab18d1491b091ce01aa1373d281a77dba591bd9b60e0cdaa98bff48c6af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h413e2cf531669c01cf7d93bce0cd08acdee43b8d674d833247273360be6cfc2b60b4725ed3963710254c8a68fff26151100b90074b47a2e4709b80836b7104fb5e850d190e35e28e2c660a31d503cff1985702d3e1c2b69e946f5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf257365f14bedc3d62e6080be44acdc2170f750726220dddd95c83adf089eadc7ac56350d4c66ec1ca6f79c5aa236dd05e28ffe19fc40a97c5b585a567253b7776d9616fb2b55a21dd10793664066cd1a4066fb143f25461315e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee0c9ad73423b9744f7dcfb1d70a927755cee62c55f74e1980312f44c42037838331885e1bcd0288c87a62f96aae077e78a98b5fb60d996592677cf62463c29dc437bb67b5d5b8fbb1688a0a61cedf1f5c440ab496795533c30ec7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb52499615abafd2140ed123d8a9eaecdeb8e8a90f29632c3b44392072c9824c84f0e4152972367d12836d3a03dfd474102b3eda970e6537540cd63b38709e241519ff7cdc8c9ee2d81a57636b77d82b10bfb89f01fe6fc5f44b9d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c15ff4fba31ed293b57352a044925ddaf00161f5c81072c6c7bd648c414440687e1a97ca6bd85cc34b77c413fd1493926d835e22d8d925a1086a5e1be971391ba38ef1621c1f80d8337c4ef308a0bd8c85d5de5ecd5d579f07b71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b7952c08145df0a3deacaf89ac240e817d804d2d2672129f8829c2c1ac52d7c8c59663f730ceadbd6de6f82ee2534698581ae9c6a82c816d83c7ca95da0fa903ea0b27af5edc2ebad6c16f805fb3a26bf562c9c34f93e299c58b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187d50902e92a894f16c9ce92ac25f28be02476a77a474172ee98b8aeb07ce3d69ac93710f544a1ab6fc468ce3ef70ada41cbf4f924d257fea3254b44914a37893b37c431401d8db50ca3b013be31b91e556b63eebdf8835c71eeed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ec5522a1aef99818e26ed1063e18ff85c86a50278b8616c947a2261710bf3036da4f5edfc0a2d356361239d182e66a47cdfd4bce4880ae257f0a05a7c8af6e31271ac5194eae6cc8db6ade2bc0c86ff9c6cc511fbeb546f9a63e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7260b3bca2c2adec5f4201dba1a16ee5f22f129392277c218c82f5c70fa08789fa97548100faf12eb271b1aed7971af03b551fc395968ba925c2a0424956e69966bb70659b36e4c5d496b7316c5fd8c7fb09358e1448f582c30e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdf17bbed2d904f5fa1146039865b11be9dded400dcff9e227131e3c3b99a76ad864c443dc848ecd74f8b39729aeb4bc1d841d2a839b4933b4b835c832c54f35b9ada69f1656be26e988b8d3d184a237d5d02d5323377bf206ddda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e6014c41afced060f37f3fb87914c355f6b5176f77b9577a40f02b8c5902666cf54129c9c22379d6aa896517c6940c71ec6abc2cc3df4e30b581667a23b955147c9008d7bd8c41b54651c04fdd54e79e90297d510c16eed69ef3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd3971fd2078339e4e79172acf8b175766ed78e5b874f0c500319935abbd64861ed8bf80efa7d0d8efa14270aacb4106cbf50a680771d9b923b7b09fce12779d319eaf2be620c2a3bd84cfda05142271374b400ff326ac95b6dffc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a474d58840713f56b223e68fa67e665fe327113326c09b8a09903bf4f2a2ea729330b060226f0e6249ab3974dd7abf1ef78932e292bc80d9eec48649c0803053dfbe9514b8c0a9c31c2fb51b3c807d456e9d21fc59581fb3de5a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d72a0ab9aefcc76121d5d5c5ab9efaf17f1590abb54c096a233c3a8595139a0da9c9b65805e74d35282d5a1d3f361ea8db696103b44324f22d7af5ba740a7e39c11bccc1a7cdf8220d99beb102a5fce7282a6de7cf88a30f8acbf5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdaf7a2d381584b02c18e15c472d77ab1eec37533e76491eb104272e06fba9c8fb2bfbf4a91de5a94998bc7a737be0d3a045980a3256e65bb5676e09c8fab30d05fd828201f759fb9b1fa3198ce73728d3c51458ff6564cc310478;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9b54a4af1219e91b72265364b00f35514678065bba35497c65ae89fd98db27d8d416350a47bac1dc4c72c7d0c97914c54f840bd3abf6711e641836ee33fbe274db62795c7470faaa6a9331090ef4d44474650b38090c262536db3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6088d9f9b9a4f5c1d7ee0331fc3b8c81b09b78a7394930353c7cefc93b67f0b409cbad966e8441b78debd323a39a5593481620f10874ccd74239f255e71ff908e00ffbfcf2afe7a97686e7481321797a1f677aa787362838fa9121;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1c9c97d1154a0ee56d9d3568933af5a9f6db363ce9abb5a737e27a49419b82307eba1b32a9c36b48356b12340e465498c5a03a485c527c3a54ea6b3ccebdbfe5fca6080d43d5fb346327ae5b56f08e19b0c510430afd7dbe229d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173d8787b4b86eef1167669c8d1e04db7ee26983c433b188cae74e62918e9299fa42c2ba04d85bb1a61fee92164d24100912f557bcf45d980d76c49a8dbb1157ccff9b1bed724d8ad63c8513ea406db1ec5e2c51d45414edd74be51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2439c4ed72e25de9fc0e74ee5e2811a66b7d2dc9e2cf3615f68bc43947a543655b2d599cd50c6fe34b27edc7e761ba4491e4eb30353cd6169ce9a53d689f40a4470f9868e27572e49f34dc108d13e8fa1d353fdca2aaa01f9fe36d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89b318b9373d2b37f0d22fc06bbcddb4e4996f5cf974b5c8f879de3b6551c69be348f4c3bfb68709aae6be8bff3ace28fbea871f31cbb33605d11ce813c6dd1f26b7bf5223dbf7c864903d12101727f32d4539823b303194099fb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f8bcf7ff58d987ae3c0a717f75755a91ff94c126cd0b4a11560e81c0b94c58672f83d27afe92094d85a77b0d33d3ecb9bf31e56bdd52649595fab13e4ab762ccf5a1a0f926fff317fbca6368e80014c3885b55e0e7778e215b335;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ed3deba1fa03ff2312b7599094d138e7526eaf96c218fa2e838e39d3495aa9500c874483e9d158a9243c3a30143bf0566639e362ae6241e0dad4b21932bfa5af2ae6739e57e42bfb36d8e737a83c50301d03cb0e3781d15330284;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1650249a240b9bca6a7ff8b84808e9b17d96a3764c38bf3c4df0c6be06558eee02f77425d2d34848eb1c37264f522f58dda89d2983f618914862df4460b6176f1a61adc4d4653b43096b0fd075093e2c9b5a4c764c3fc9a1696c77c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5835e3c7e91fba04cb209f83df0032b951da481288f01b5fb9649816e133c79ad22fde125a297dc0c229332db5d3094d13912de001f602e71da80297e550c7d0475c9efceeb175116de78e10574032c27a659556071a84569b8165;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea07e589c64c7271a497f017530c5820d1d8801b1ae7cfe6d4e79ecc9f4aaa202c453a6629ca407f2ddcc300287eead19c03cfebaec772d7dd6eb1abfb03cc04f905fe65a5261972ce309fd39c63b6e133a4edb429d8b303d4c064;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8aa682c461fccbf2cf2ecafaae549b2840c4fbc7236074875d065fa6cd99f7b10dadb1997eed1dd7885d0680e5864492a74584e2ce55c404ba17d860df80db8c5dc82290f4377a640eb2439c8062d5cc2264e23aee8a1518c6326b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ea5b727c67e2b41f61f67fdda94b9313e076ec9d6379ace54a253a59e087df196cca924bcdd6850ec83256fe7f30af055bd9e9e4436ff0e133eda0844e932d5d0714ee706a2be47b406840c04b13729f88543e7823299bbaa696e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2e681e1a507c837d445b5a28ee0bbf318934a21574772bc5e0fddee5aa0899f7e0527eb96597752508de597c69822d67d87f430547c74e853937f5e9e11ee597d3df31d6f02e757832f65f043b572f7437ffec6897941975dab25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7448582246d4e5ba3226f1f39944539bdb6f84128ddc3364e75cc484e941bacb8f785951cd144f1656ea34f9c71fe1d49c9f124528ebfacbc6357b41edf5d173c2a9f026859721e8cf19db8a0569935fcaa6b0d8e294867180ffb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f3f0ee94a67b1d7e908fdeebfa4365263030bf01525d9a632cf6c5439ef91782c885227cebe8140b4b5bd615b3c02c34bfdb531e71ed6d635848fa727499da99d1746d5da42af3e9d5eb738100f5ebbf7196fccc332355db116ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9fc387c2185f67508871cb791c3ad6de70c8d2a32e111c77c3964699cbcebd55eafce7d96e469a220a9be602f1d99ca822bc13930c91a516554a4304daa8de4a3ad6353556689dd6057c4b82320e111fe2b8a8c2dadcb5f77fd42e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3627e3cd0fbb65bdbaba303c4e3d33e176806b377d3c71e7f0e39a7bfaeb7dc5c040e20f708dd75671717088e95afaa4dccab8166e67af21551fc51645be7a751492b0d00600fb63748ec11439dd6affb78bda5c4849e5a10e5b6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad51b204e999d0c05bc835babbbfe5ead04e09d199ed2f0df270a38a344c2c9ab25e9dd46d8d30eb430ae8d3009a95403dd055a51f29f233daf76886def4f987625ecd5c7d655190aecbbe01b6050522f70a8d40b9e8d493cd43d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6f42680922b284db422451053332db807d4ac07fcbd9f2a1b72ebf62d2c30f400cfc3cdade67fa907202a4961f0a2cfc716d4dee17b00280834fd26a2a553401ecadb9ff7cf797915c15d47cd9c5076b4f01c9f7674dba23c44a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2748202a5dfde80b6c94ff77b26a327bc76d9eebf0cf0466529b1279b1addec7e80142bfd40e824097f99ef7ec1f54395fdc2767b346f2071abbe17ca7dd3ca432e5f8739533a467f51069a21421d2fb8d50286b83407e86b240f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9197d16150750136240e0ccc6f1fea798beebcf4abf8a18640b23f066cd7d9501666b2bd0e8b6a8c380673f7e6ad0d87d1acd22bcddaf4f2b05af4bceacba4c88464d7bcf9d943cf7bc71abb3af601a103d863347ef5c16ea3d8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108a6bc0e5a967f2d2821aac057b0cea5da26c159e334a15ffc3c7861a33f8e3450b02e15a38a5043ad8624e8aa64dae251e8acb56038b039047098fc4cde241a0513ddfd80dbd2698d36735dd9ab799cdcee362969d5beb74be1fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f8023bb7c3ac2315232e7c6f0a97079b66c6b8030e25defde85ceea3f4e28209e8521252e1ade17ae01487248669d8c8fdd4f56f190ec8d59822c7b1fb8181dfd4d8979ed557ea65397f1ef433a389808caa6b54e6fd1b9e77c3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173c49ec9028d0f2a8babf8a24898d3f417a396515fbdc141ddece1222118158bca8aa4c85367634a21e92148d30f73973b3dd0218c9b7683fc1b318a7616328a3f41f1f7c1a6caeb2a635c0eed6bb6df907353f5e4489032d8dfa2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2160bda9e2729506e67de85e5024820729f113a581c78ffad0c6408c02f9ed7d2359f96508c01821775d4c28a142277464684e90f12d8b767af2c8c89ec836f1097be5cf32a33c0c614e4d1c095ca160968107aa7dbff3676ed70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b79d14c1763f308f2a0c788dd3a6fb8dcd747a8c53cd6d1ea44a0a7440a1ce9886196ec87a2a66f9d29851313d645c87b1a0be3ca7618d741a05d344ce36a26c9c01d7bf319bc50b55100d03a63be3d037e2bc1f8f34ddd4b020;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h120c299a17bbcbd70dac0505407d8364832522ed9e871cc8c1fde8aaa158ee764a2d1c36e7edd139fe6943586c6fa316005b2978ff8056e335e6e86c192f132824904fe13988e5405f0abb5f5bb492ec5f3885ab54da8076469996e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa37cdce81cc76dfa56ed8ff114f2ba61b4aedf05e88ec9cb90d8142d53119b5406e8a8143139000adeb70f5dcf8e36a81c62093066ca1fc234b94694fe6edce97ecb14fecf0f563d6766a46511a60a68bf3b72e9b1ecdbe615c81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb8f7628f0a3b12aeee5cf6c03f09e5d9eddf489dfbec084f993420781781de12dcb8a67ae3a6b9f55cd0474bd26729bf27bd58ff6b07b9ab667f911c575d6aaa84a71db6d9e035518950fa38619c19dc9e8e8588bd8001d6bed20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a03cccc71d80c783d676f97a89c9c921f334d4ad408d7409a16508ab3a0b42d2686b01ae81f147e44d38c7994527e2b471d64be780699dbfcf80c6b547a9c701d2c6591833e8c95a4e4523e27dd0ec425f801d8de46be5506e1e0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10bffbfbe5fa3e357c6f509476131445990f662b23370596bd2def073463688f492f97ae52f974669ce5611529beca024acfe307085c6412c330f6c972e4cd56d8d8bcda530cc61c3d20e352db6a82b081c4c2ef3fedbc7c7e99f39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cfa01ee28bd61a74dd6394440983f9db6eb61911d1709fffae6bc7167938ed342245934c23995d37ef3ea733811aa5119ff9a25b7319e15738759498679ea5b6fd39c5199db44f12096f8ef8262885a80901d8b4396ace086428f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7a916bfddbe7deec982fdae38f6fc76d1750b7d1b3e5f53f8f0a43afb8474262280d7d2ea817e2ed55f3565d97f83fc98367c74d9566ae5e1e9398271bf719a615faf2b96766e3b34fef5837a39d6f09b615ad58ab707ff40320;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbf82008f022c0c43425d82a650a9860a889afac26ae005d850bf662d8ee4eeb60f1502dfa5be664185ac66c90a1ddbbc4b34ff31d65f100b7b141f18c4393c7ffc774266a541ccfc2303b45fe838a933e18e21f3843788b954202;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b93f405094d2eba87d2d8a70c5e6b7800fb3b06f01b748146c6f2dec6989c908ec537966f7103bb9dc35fd21daa146939dd70cdb1c48c4940cb01e2eef8ef056cac986ca5c2d98325d6ede62a6155364827ce6f943d02f600fde17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h747ae76a96c355c1be39c2db1c8fd5997b916a36a80a005220b1aa5324cd8f8b18b6f4f8910e1429510411cd6712dcc69b6e7840a5c17738ab3fb814007c5b447614422b8759da479e47db79b23e476e199757bf0552f90e9f1cef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1279e37d97dc148c7b6a78a74fe268bb5e411d71e9097137b4693aa4ef0258c3658052052c5becfbe5760e5d312cce328bfe1637902066f33e97f6ce14149f61fab31e09461cfd37630a43f2b5c0325fd35d2f7612d66891edd0117;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b8bbd65c9fc7313c7782a79e9c41ee52b4d6c8fe317b72c611ac9a843075ecfe103e625dab8b569e4dd60c3691a096f15be0c8b3a8d35468c26a2506ce777e21c282c9150cef2f6b045388ce2127e8b7777fc57c7a9459bf94d21;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1623c43608185f40434b68c154f91952f1e1b94dc6dd06af92eca807eec62849d3839ef71013f5d8b996374bfcf3232bf97d0c7ac8e60bf7d71e9cef21efde35e484ac4793e2c700eac58134028f1298937c26e1fb6e9e939a2ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc52685bca182f6a97ae2e80d3de946db67855e3c1f5763b6c3be70e8bf30c92c3979049429a75168f99f71ae848cf7303c3dbc98eaeb62e04b12b1988ad619c5e7e43c178b4c79d2eeaea901d90848ffe9ae5e49e1220bd72f29bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca4adbaf7cd1573d25078b0a9a4ebfb3c991bac0a48ac6a44db6977cc389afb59634017c62b91c8870ea3b76809ca4db60a4b5e68bee66d982e026eb393f433b692eb339c1b6c6040683f6cae8d755b85247c6b67724eb25fa0102;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb687917d333d9699779b583107fc15dbeefd4bf95c8535562cf91f25e297d558b6c26870d306bbe89da3804a481f050648253b0e90d18e9cb9815badf64d35ac94e48b8c71690b0ecb26905f8b39ccdf79827703dd7049557d1670;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1735a7f7dfa14620235d6b2f7403757efefe57e9f912a10539c3a795a1ddc849f0319619cbb5efc3ebc7a62795c159bb7fc5ca193927b2c747e61069bdf6b2838e2ede068766027b8c020f5f108d5dc1db771e9b2c7275cdb84050a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc83ef1fe7848020b92f44d5bb511f8222bd4cbf810a72465f75bb2cd4fdf0ec4b1c910bb78b6bfc29b355b13db12cff5d41b56a857621ab21cb27041f9baa71718221f659f159f1f47a4b6888601d035e787014b99984d7f0974c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd248817aaaa3541ff247007580bb5a967b5c9c76e5b7230aa43cfcfb1131a5d9c30c4787c42f1bfedeefe75ab1043fd894d7786e773fd4ac98dd8cb63b271e404651e78fe299479699e95aa5be2e8897d191aa074d1f04e1e5f1e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee4d5f66df9d865d5018c31a392eb6043fd96f7a7c42b96d3db48495980e51ccec1525659988e1f1592ce02325653b23454e2309f5b16bbe86820e0d2e8ba50a2155109fb384cd6359d28790e4ea81e933f7862b0986c56ff07e9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122eaa2e49409670387e57e82df7faf9357702afc4717a505e147a648734fe69832923faf5f4f419bed1b42cedda6c769597087231ac49240a6ae5880cc8b45cf7463a3760a5f443aa30e02dc742c4801a6ee81437e6c06f6db4a63;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113f080ae0575a292347b29e71633b2b9c572ccefc1611e69b7284d6f0850cd473e16525e8484f2346bf0d0c899bde28b50de29e8707db078fa2b7101cab6a254527aa6c37f9118112e12e92afdbfd9aebafcf8ae608fcf2e4d9684;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a2d9d593d13d8ed8d0d67e3750c3fe6c26687b8d468cffca7aa077456173654c196efee04b911009c8498acf7b1c6b3bf7ba21a4b3a801a6918e1f1ce8d02cd732d966c98e53b2c6fc99c6154c5d2def52bb64f4ed7aa69acaae4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcfbdf03dbb472f37c97e8c7b12c70a5f9ce57ca9abfd7f4f10ca24702c3fac3391fe58ca49d792c80e320d0b4c885e88cbad0a6529245cf0f09ecefab7516c6af4bc268c646130da8bf9d0f3375f9626d7fa0f8972ad9d868a1710;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea7232a73a68a8294ff6017fdf03eea86db0087f502965e3aaf38b314e5af9c789df20c8a5dcc717f7bd248f6fcd01353d3a8391fa4cea9c84e192247982c3ad1a7d349f2aa8d3850b5a46988d6bfc16c84841c5786f09bb774708;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fd3359498e4902a59c00503a1a71a661f053132a15443ee618cf6c0792729fee1b199adf50545b569d5858ed4efdc5db1254d88486f9aab6d3514ce58af99158c939aa730a46f44696dd5955347de6f37cbb096e43fe315f96fe8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1941d35a5543503a8affe11b610f523bea40993624abaa09fca175b853f2c9c66512921e092ceefaf66cc94a60fb0a37afacebccae93ab77c070c5cebc8c0df328f77b079823812c118183b40127e145988ef423b1d323d3d540918;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1151adcfde381578bd95ced044f70cafe2c69567bff6eedaa18904fd840e5a0c44e27b37cecc91ec0c5f54fc2f1d2f658f2af9fac6059ca99f6b2d1885720da5b792594c7f064590fedf55794f8ae2bf67f2bd5c5a6a3342d8ed6e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cfcb4c1b28d981104b82b7f6308b03827035a927c2a0dd16b1278798192f631f268516e79752d6aaf07927d75672c56f377652368d03a519e260dc7cca08f38fb5a64447c0078759d2238cb2b6b997389e5218c8d7557a8dfff45a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7ecc6a58a6e1d82c14ada8c6b5aea13837749922b1d1913635a9805de530d80377d1acaa05866f272d25020eab91c4783300b67e7520f2092e312cad034e5c4b94f984c4fc4ef5f9cd3311bda8c324680df8cc3deb6a107bf1257;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb71125ab3c4d3c4e1e9ba3ec34249c975f92832264e4e5b48d5585462f08271f68d72183ec5503c72f5a4e8577124c7876b8e510e7d95c722296f8056ba08476d89af21082f139994d3cde3480dc5f57f6e0f1697fea820e42e83c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180ac4c3602c0404b61335e6bbc6a5120193e3afa3515477fb1a2d948abdeaca806215262f6a59de5cfe40781f2b2ad87015197e5cd7f76ffc1fbabb3c4ac6c4fa2c09bd7317ca2cfdad33dbf46ce69c0e943cde1b42f9c3355df39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc094df7bd1ebcb4a606a6b15a0933aa4fab0dcd8ebe381d48a6e3dbeb856864bf6876d7a60803f593403e0b2eb583e7e841c31c08b837ffb6fea34d662bd44b3ddd634cfdf538e48b3243da8942be34be04c7cb2747dd1aa9f6cab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7dc432df59674ea574dd01f9d9f7c34cfdce4bcb57a2e435fedeaba0196670c9fc95e4522c7f112e67f50a8f112ce7d02c6d44d14ab43eded9c4d935dcc667d4ce595ce722aa512e4cfcb6b0d1312a184560d87f8bcd75055a759;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf3a134cf8e28b2a383a1bab1f07eb5fc1fee97268964fc3411d7641dc1e312f6fbd6b1f3b6215c204cfb417292e7d0a84523a7047be7e9b7927c340cf8e77f97d9139c0828449fc9817b4532b05836ff00d3df6cecfaf26c6a0e28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1078b65390f2766ef7a3ef087dc5ff3813e9fa344cc3aaa90ffdc479898a5d5dff113db0d3fb79b83e5bbd688b003cbfd651413b17116b3d8af5c81514717423d1e7af0238822565b89053a8cd29cab4b0d05759905bc91018ad9bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec4d905d6d474c5f590fe43b8297866a1770145be2947668ec3ffaac52eadf9d027d1782b243f7d2dd765f9189b3e79dee4177859af8abe77e4efc8fac9f3f7a906a9338fd8cbdb8b1b1480211a0d47ec6e4545c1e7e8711814541;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e4636ddbe42d67ce8cadd3cc45f86b880f710ce1e4a12c3ee4152d59a64939cf30d717d1ce6747e6058820b4207c15ed2c76d82b1cf31445b0103873358cf8de10b0d0a01d6ffda6b235a2691cd77b217877bc64718a2325cd718;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2fb7c942d17a3d285b462a6ee9f5f3540a0f5ee853755a8dafaa37c199923ae6be537b6667d2fa00f7e1add5a839974bd6205c8c43504d6f4c38635d84a9f02ba8ab8fa1f6c72a2f7babf9bf26eedff59969be348e8d05dbdde33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a6160a1c302ae92fceaceff36c66c33aee424402f6b2d752e4cf883eb77efd29e2930f86c73a02a884c25a433789fb57edc61a707acc2b8b26d11d1a71435010a9ad464c1ebb9e270ca7920b93d4f24d388e77959533ea7cf357f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a8efc7dc6d8af98581b8fd423d1ba006ee4f5b50ca8259f742b7f904ed60e354e4d90da945ac0187cda1f6c745a3576df69c626a167a743598e4982c2abf1e9e05d674624e961fa88e3707f60e95d02d699c47c998b93fd31fc1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9a502beccd50826bc709c6c9c12481d47fe78f626b009dad0b5ea484eb52d28d0c5e5cc38a5eb7b728dad2ca367b12b81c8d351a9a5905c2e68815795c8dd94651c0c68e17e0a757d7dab18a6f0d8c8f7a435eceb02eb955e6043;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9b44fbcd2f66e029f5e1b4d20a804e5847dedc6fe859ffa4f4cb09a6ee60285526341381c5c4fc742f1e7d3e8ff2ab881aa4fd92a8d6facea175b4b6e23c94999aac29e17d968e5baea266b96e7cc132c34b891f37c25e5fa8cbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1041dd5017ac71a615a915fb7af2ed226fcc1c501751db71a1dbcb117482d11a962c2a0367b1cb329e9dfa09b5e71694ed013b920800f26f3eab713f0b8ecf9186d0d80a6aaab0ad6ccc78bee61e688307e74d79ce61ec048fca9c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f1e2088e09c1df049a23af2824fe9411db3978c66a71c158e557f437da565197eef4ff35ba06c84bcc808294723b13b494d492c9b18d6cee471fba69b29431beecae3e1331d53384551103573eba5b901cbef24c6dfdb1367df6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae445b85c965d6f75f6ddb2906951750d72ec9ead7801490a150f56e62498cbd0afe3fc996584d155fad07ac6fcb2da7aa035138539c4945ec2d573661bae3c426c186a4bf61d739825b8edabfc1a25ff78fb0a59c21932f62fbe3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1787bee3037a7da5afc19cd9290bc8d9de77f0efd5e29a8467ab774abb56adf85118d3e69ed716d14b6f59c003a7cc382250df90f1353d71e7067fa41349dc5debea005ebe2d7bc70353f29d6304ed6d69007a62b1bed5b8e2617f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a1a057445c56cd1ae3e25f84e5fbcbe0de0827c7d314f7ba650008d6da36707f6caeeec71220c856d51a80b82e5c653af41c75c6a1b569b06e9076852c4dfee9ed3f7094aa2a0537cf7899011dc4d6edd376392708c0f056036f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6fe5f1fcafe9d55fd389ab60dd59e2c35618da509b03db3f5e6d8285558091ca600b38ca5d96b733c84f4b4b5ed7a0c988783623248fc304207f057d5b9e453881a2b8bcd024e25f8091ec26fdf87bfb441f6c67e0bd49a10edc1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1093f48d9088d17987219ab40839bbf93fb26e3f9cc462d35ded4c8262138faa1670ef767038a5a407a9fba3df9face3f9bf05e377319ae2c9c6213f4a652c56c106bbc5d00ff37739038f090ebfb071af5c8a83bc1e11b1ce2ccc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d3f1fa672a0df14573f9b6712de353e94345e9aa03b20108b03b40fd88ee1bcec46b448429c8d3eba9fc2b1c650d56c79e508079d4c1d546f087269c165ede1a306cf255c240f00bdc97af0d11b3f25ff2223512be4a3758526c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5817bb4cb2836eb1590138595237f4b2c039989e8d4abe7a26d69c36f5f4313101ca1b1a85f77e94e7d9ef31cf16dd838f080121df6b8e647e4c4be7c5ffc1aef89ed62f7278a54f401a70080c3036b4b6ed0a1261ba61e3fe4959;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9ee9be4e6e0a679220ccfedf143e9a9437f10e6ba5032730f6695867649b382e289e90e6d0fee3e4468a61e64278381e64cc6739e64cfd873437f5e4fcfdd577b4414f900a28cd7c1b916bbb8358f32e94b7c61237c07380c2893;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a498f05d985a59a19bb9ea2a6ca9a1d8c48f7c4c8de10af085286320f53a6c93385684363d4b3f39c5b94d33f1733340e474250a40fb0521831320c81b7cd978e6a5418220de6a3aad2936e33a71c891d9f2c57fa8a660ea13a00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25c531bff770dd836de193ab14ce893911e31e332ff88fc22d6938b1dc7d91499d2d6ce66ed204c70d5c82b0083285db0121ca50ec0179a2943ccabf9efdbc9c2bdf8b58b43cfd6ffb25037515dd568d977432e01bda545e60548e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188855c09b5cfd1f68d2fa825eaf909bbed4521b3d35dd42692cdec0981183a128107bd949b50ee8c1e5cf3fe126f18bd66140956ab09d52e72477d619f74f177dd64677f40e5cf22872b2080b9525cab9fedb535a5f098a4856eb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1131f8203fdc09d98fd2965ea2a0ac8199a4a13480e80070b54df614cd08029a5aa15119547d1a2ca71ce7da5d8d419807fffa462970769a50312433be2bf21094775348961266053b383e393ff824ca59803c1402f58db8b5937ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fbc5beff13efa1f48725609c5552bfa2fbf8a52d78d0c9c0e5805f52893086f706a93d6420a8b007e7e7cf932cb6b5614cc5a41950abdfa67dc68c954c40d0969b99640169f397f8b72227a5b119d59121c97c7921921d8acb296;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aab0a01545f4beb0875073ebf1d69e86b7ed3800b853878f5d5ed8028a3a1d729ca473466f069d425de3809d893b03b67024f6dff3fe1c71985de77e069cebe01fbfd6c620bf8d954603d2645e4dc5118f082b7a62b1a19002a494;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10de025e6e150eaba25b3b217a3c2ddc25d5b41e73b7e4c5a3c3dea92af3a0dc20e221abe1676f19eee48eb5e4851f866883fcb86d3fcbacd3fe7dec3a9acae3a5214e599ca992f7fd54351dcba428573cd14f5614810b11956f5a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bcdbabf4c57c8ff74c9d1c0c12314ae11093d31873a5dfd6531a22813b9c30c9c1d46c75653a829353a8384c7076e722b100a51bf9dcdbc6c83ac1d03dcc16b18ceb3dc0d2b753deea9fe2715fddbcf779cad7a8f14dff421fb18a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dda57137ee8ac250acf91773c98845f2c0cff54b966dbfd0a2b2fb0ae7444cc2ebae2e4c261810eb6b2a0358fc39db2ac56d6803c265ea11ec16cbba0fda260c685597efed08e723aa0951387b0ead65284a7c55c9df11c7af101c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f1f4283b3d167869c305a3306828b8c987c4ae87dacff69850a48b9597f8d51ec6ad33c550e162e5797fc806e35b514212c5f475866fa87fad0235ec865eb2e699804c08432a30142eea225f770850bf7f3a55832d07d69ea5ac5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffbd73b9a80a5a4faf75733e856c0b00d853da36fbb826f1bc184867ba88e4765b4dc45740cdae1828a17c75a1b08173598843b2b834e23c485d95c216ad6480f0376d743a3cbdc3bf56d6245b912eb9b80524c4592252ef3752ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1bd7f6b083bf064e4127e25222de63374102b2863876a09ada84def0c17935dc6ccb04642c1ecbe62ce52848a391f660e03077a84dcc22125706210b46370179045cbe4fe51478609fe69392f5b8e728cf44adf01b86a95932207;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c95518fa87555502111acbc7f51b0ebee05293f282424fff139d95c913e94bf8bca88f1178321ce6a600f65081b132188a9e8fc2aece5cb5ba2601c2f1ca506b925c8bb63c62019fb54ae3b94a6ed108fc3ebbcce347b2bbdcead;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b7d708457c399121f9a4034e5c5d1fe9fe6824c0b1e190b60673acff3b6569c00d6c0fb716aa3743b78f60100d586698df974e9ae806ed23dfaedfb3c516f191d0ff67bc78d73f6a575e784de5ed477d1e5cae4bedda82782972;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7bb7c36d2a1dea64e975fd09c8c76083ebdd0f1340939cec860ce9828eb175c74ac884c51ef178e05bfdc0c27f6c9923278fdc9063cde83b3875301ab378f160450d1eba338c3651dfcb394a4ce69ec53896a89b8553a280ba96dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a4043a387a89bd23d7771fe32126ffda66ee8c301913f44872e29a6cd5dedc2a17d3e080e4518985566447bed88023c277a6f4dea076b3c8229c5271b28bf9253d5ff0d86e2758e9f31b0ce0fa9a605a074bcd010718c38218188;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b31845f212fcd36cff4412d2108f7cfe731b51032ec130c65b55ebb34a112b9bb59de7f74809f13e53ba2ce03acc3da11a60a94360d362ed8a70bdb393917404c451366aceb29480cebac3fda919c911b25398d4595ff6bf45039;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b8151d0807393fcd2eedc993e42f8862b5cae565f327c15e18256fdca2789f08a232ebabc4812bd80006704ad7acb14ae8dfddc02b16c390f20face7f49989345d6ca4996f71513a79286805e8f1b9d4f78008d2e05ca0b2fb087;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ae15278cee7a682736ea24c01bd701908870f553f15d99c33759d01344802ea35a1b3328fa636ca9c63e9bec709ce88a79a2bc60ff1fc649fdf2ac5e4a300458350a2bd6b567032e76acac9f7cd9ad39a507b9b8433d013bc30f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9922fe8beba955509636dafe0b4b801b17ce8701fe29149f6994bba702fbf630c596ae98641b0752d24702d9c4744854318af26a226619119b3fd26f2f912d6ed82f41abb58713ed56a8c48dfa48a5627dd58188ae2f0a1c01611a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7ef2c4facaca98ff46dfc387757255ff5264ab30eb1f8218e5b6f8bf254d2d72ef756c9036ff446aaf0c0ef6dff2b1add471e425f0a7a115f5e8e138ed0a4598f46f1f13a058ce2c877a33e3788c555a21c53e360ca2ce729268d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb225c0cfecb025244a35ca625f2da9039f29124f2f8cba24f42ccea30497f3a4be8b67a20f332ba02bb1c5673aa430fb6616570fbe09c3267ec321ee0cb2f91fa4650ac5b47b71f30987964f641d627bd379d2211624df0adfbb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b3b6660f5b7ea24712c0df9fa74336702720f4bd095e00b61dd9d267b5d8d5dfcbe446cbd1c6cb804ee8e6450506c1e7588aa9b50d30587522eea5a852630990f2ac51f5cc2eeffd5726c5bb98a0812f8e12e8ee6b94abac96a51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc915f5e48b4343e2a85b1250f22fc7969f3bbabac03db7303d242a49c07f83d48917a95ee42742cc9f6c5a546066a5fcc9495c464fa49c3b8c0bda306bd224e5308901378ab2a122f382130a8a3950738161f8bb1f6f94458b955;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0a9ae35c86738ee20c0b9273097c1335a3632c1e23c2a503fd9cdd675782400058f2b5a3e3f534afe056f805998ccdb8acf6a7bad98bf2654ccc3bf0276477b6b381654e7b131c287834afa462e4c1d32b6616ea2d167aa5f23ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbde8e51da914b8b75c58777edef9b7985ddfbad15ebd84ea0753efffa6bd3826aca1b39facc53aaacabae1530cf8a7342c97335e91cd0dde46a64ca35d2baa7ce6e3a5021e180505faa4895595b076da4277861a90e14e0272589c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91c0c118c875e7f3c650d3b329b25e42424027e277d90a5552bc1b39459926344a68a56e774b8682d47577e60dc01a8150d75711f6bdee735fdb1a5968297457864296abfb1ba0f5c690e8e4e27bf47e9f9b7cd97b2ab15315151;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e697ca6efa7133ed2d4e96a1b4478d8c11b6f945cc6a9d6b0a63f931b96d6a7778d55e448b023bceacbdf848f061e431b63471819cbb4405b016d8b291e7d80bb8f45487ffdfa67bbdc9d99cdedb96dcbedef583d1c75aa2c29519;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c5c9ae4e193dcdcd778daa0ff7b54d49acfb6697b1bc6fd450b1969b452ea52d33512cf5584cb17dadc38f9ce67eb81582d9760224a027aac84d0c547b755cd579a2bffb003075853c71b6dc5f6d7784f73a555e3bd8120f98319;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea3b959b45a12f99a546d99c86d0b5333be598bd3c1e85f059538bc2de5a9e73ec4ed74a748c255283d5a93cbe6c32b8ee9bae0113798f73918bb79e8d1aa884a6c3fdbb8316dd7f82b15b196051a05f0952e48eb5e285806593bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f403721d0fd4e9b7432711e23affd14714026a10beb1c4db6faedad4e68dc476a626e2562dcb0f0dac6fa5d57f65783c2378234ee2d7ee7778543ab5ea76aa596382e0728be2db4a2118000844fcf4aed16ed3f1a808c3612172d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h60784d0b481a0950c30dbb66995be93cc132efa275a9bf96e997723e9817f73ed03fd0f00c8e193f75dad85cc52e37c7f2b7dcd1e6a3acd2e6964241ff7ef74e2752da48c177f0a8659e1664124a6ee984e097f391f4241e416b69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3742ca2b4a851770c091b318fa5cf10e72e057f45611374b922d19628f0c60edd43a9dfa1d649a66a7a8e8bd6ae10c07f5dfa8b29f18409523f815aec002140cbe92c333ae83309feb4957a92e0cbf82fc8da7b90e9158f7a1e61c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fcb0e64ab8b1cb4ceca11619024d225d2547d0afc173c252068f30aa2d72da87a7f37bc3404653a8e2b4541494087f09b177182f0874b2961bf284fdba9a21eb74c648734093d1d3bd6cd87611525c2ba06e02a73e02ef673bb5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf67ce1b62bad9c176d9bea41f6e541cb04f0ae9c118cdc2f624fba0c0493350ae7240f9b5ce82688fc20f0ecb0a941b340c96c5e595fdf9c070c459ee90e10d7384f53250aa6103f796f2c97de0bba88137c332a988e37dd006e49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d057ce98bedb45aceadf0e14fab849a1b9d36d6e12a19b70ef53e5b5d169c7b5970be96309f0588b18887c91312f1f2c1b952d62d2dbab959379bdd73fc40ef3c6f520d36546dd615fa315178a2baf738c29e4ad985bfe96e5a29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28a894ce67ba0946f5edc1985992c36d2d001f4b286e94f1cb6be167f9c99359d0de2a19e2a21d567ce65bff40f3b692d4a701d40036c68d0630e5e5c76a5cd76fd44f3a596745015194acbdd06c699c7f92277ce032af7815f3b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14adfea007340f620e805ff1cf40cf99a1641e4cf88c25482de80fc5e12464b785d74331404604e8b32ddd7a6662910abdf3caf198760447939f1d2e92ef30130cc5136ccf9e96cbb3e48c8318ed556d44ad80af3c48fa5f6d255de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13166951380586aff9b2bf61e508c1c4ff8a4ab194b36288597b4f7cdf6ade619f7f0f7866a0bac4a9524e8ffc35dd69b77cf48cefd151271b34dc22682f484d52bbf6f9b880c28d896238c8c72f6fe46e4f26661d6d2af7aa56ef8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d2f0b7150ee0e49f45ad9e192a169bd4acd492a4d9e306bbae7d277c53ef066bbf7b3767cbdce6991ce4cad2afa0242907924847c492b054d766e42fedad5b63f93964260aa8b09f93f43c41f4d874399e2203d4a1c00c4022052;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h770724796a4474e3216bf6f3c463709993e106594f5c4e295a687e7fc9eaf73a400e9fa01a1feb98e2512de1dd54046ed01b861d7a734e0adfccd83973b6a8b9e1c4943a12193270e89991aca3ba4db1707ab884abe92ea20c8135;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa83c4288f78bb2e8f587115120283d319a7a244cfa1ddb9e84fa7ca6cc3c658496420fe26f5308e6389de59e15e182fe62de76ce4a29e6ae342b05153f39d7fbb465d94b84ac541ab8a09fb5c011b4c52e5e355bd9d8308d3642;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h363efcc3d952c7480b078cc679cd43724d01663892bbb094a0f62d31713b43f14dbf601cdfa71ea93e6618b08f2741dacfc0a6c66f7e479b6010e62b7b88bd069fe963f55d874698ac07c41132bfeb3d55ac93613f5a7b1398448;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f30673ebcbd5d3a92b45baea94e94452c5485ca4c89c6c86ceb61965491e7c7483d1c518faa6d9b6e8f6c8b085122de2303f359c8b73e64ae5c7344acbe7f2b3d5f29bd860e8f0325cb3250f665fb755b3a8f87b65e6ca9ef9b37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e96526dcb41495ad9aa9884746e4f054d6082810bdbb14c430be991a0bec9be7f064f11f117cd7c0a67b6c659a7661d62a5fc829bec35a7418bff8eb93ff2ae31b10f570fb8c221694ce8c30c9a69a9b11bf97ae80c303074850;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb62c9508dcb202d2d57e0a0a32f56d13574a4e6aa1573093c5aa3c1ef7993e58f1fb887ed89d1221af1e8c6b308ca41575cc7204874defd2101df71245733779ae18221bf9e03224f2e81195976d7f8152509e079c981ef9f91c64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea1ec68cfaa76cbe0f7d84735ac16e0d8f5b91c413628dc01bbfa7af65e18c84752e72b429956f2b74a5fc350397cdf4dbac7eaf79890aeb6372782bf505f31d78947ad045cc73579badf443866ad07a4f458c9991506a8694ba8c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143cd3ffa162a7b32fb14698ae646a4b5bad34d39ba3e1f3e7742cf06949db838a1b440861b4cb347e49f36dfb1a51aa345308dba9281877e4cda010b41fe6d3d64680b52e5b20f17d1b1affdd6c6a63c1c2134eb159d77a099a5c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107ef182b8409673a6b0d8eb9a850199778e76da35e2ca5e461789a1a6e830da10c1bfdbb8508a7b17c159748030affa611e9333dd7ef87ae1c916073f41af3b13a24bfb416b43ca0feb4dc98888dec96196cfc49a2c1ec483ec289;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146f96040a495b582fb5793a09a5b45956fa47dc0b9d6bfc974c061bd423bddfa8bd5303da39c607fb01eb41f3ccaf8a1d38afca9fa99e6709b193b70ff883ba7b63ca125efcf9cc07e434359c676ac0605e81c799f90d5b16131b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1580730fccd9b69bd00170137d7b484a6b55cbcd6106e96127fcb24a8d6579c810fd1d3dc70853736e2d1184a06a2f980b64bbcd44805031928fb656830c0f3682523a369c32c24bddcb33b07dae0b8bf49f4392cc4c73453ccab9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5eba1a15916f6f17ce927c6846925728142acd38636619c3a2192424b503633dd8ed8ca3e3d175c14db9c4657fceaf043efe5febd1f72a348880dc7dc0a0b0c7616eebfa3b129e39f2b47176362b39a141d3940332de46ed31f68e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1600f65fcbf3313460abee93ac6fe3678c0a591d41197507b0ce34d01fff238847762723541abec8d1649ae169d2b3979b9bf11541524ff06ed77a5e0706a6a6b5b3695a39f51464f4ca6edc52b69a19f1799fdf967c75e334f5d2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5262bc882cdcbd97bc123b7811903f0171e6cde24ab10a531f64e604c74e641eac50dac7ef0d719659cb84887d17377c16a057cc545eec3374234b079a0948c2449d0ece518cd0bd8593bf646e48305a84f298f71243ec51bf5ffe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a581f512f764e1c4664462e45a9661a0b8654e67636d8b7eb0b7e343834c5889e421524b8526c5ccce4e6b2d80cce9d2b245582949eea6b215853734cb279a2533967283e8e7835a41e36a7128a80208878d7cb2e5a2560876df3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf35a5243135f36711c22fe4070c49275bd93736a9e857721b3a9dda3306c01bd002f9e7ec62922f0f382bae533f094956e1f1df296d8c7d519799b4acfb2a0f41e2ea52bc577166798ed25ea7fbb86bc241ff617b7490404a8e852;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f34e48d55780055a063eca206ed657e7952ffb3d9d46c08967d428aed2453e9c8961dc70193cde6b82b170587edfeb2e94600dd042083275f01a4041cc3a895f6f209129fc1af3bda48fde267a745023bb6192f4ac8d3a45535329;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h363493f291d2ed36780bb1ec8e840f7120dd7b67d14bf9c2e46b82464e6874abdde797aa9153b3a8b3e7ebb186e39772cbe0030c248afb87f88e8b11005e8034950779c180af768c380b2a4cfb478f4894f79c6993d4c50c24198b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d58ebe8cfa6a1f3d241de6606c79dbca7c0c68bb5e3e486e7534b0d9f2524e61512861976e110c139aa628958bbeea783db37f81751981f5d9c52fc1abafe496e11ef0896329a90c5726cf3a837eb41518268829076cae7dd3a66c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e9a76dc5e7c9191bbf003def5e6b88664e1e43c1c44dace83fc10a59e1ce5f6697ec25c7345f35897b1dc989af5d46f321b1fddb0a2b742b7dd80c29a8a4bb5fcfab1c14601f025e36bc596ba7fe71568227ddd57d351bba199b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78818c79d403f62c3aaa61354fed2ddf2c29c981dc4cefe69004cbc3746b03504445f46f5d3cf14e24fdd8807c5ac3e1d120c57a135f6a775991a9f0e729427f5b0f48316a03b2e8dc059c7e2915c793c2f213c99066839e63bafe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12057fe87e08edf2bf8e846fb7afc56e712a9661a76bd0664b66c1a4e1fb7b4e41c93466fbaa8b0623e25d2b8536e25ad4391923a81b97445ea724f3e7d4fa4b3f0028df2a2cec929235c77ae293bfeaef5bef7706577d2b808950;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13fa2b77e307ff06f6b648e1feb2f9906ae813092e473befb75456f6b82b3944d3bc4947f2cc4bf8330ec94d11656f3970a36cd157cad317428856d964226855b64b423db9ef093313a0e7b1a07679dfe40526d4e0bbc51ce4aa46f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8a56e6366dd79d1927d981c1720e2b9f2ca9358cd5e1e55ec887402f5ff745afa1a77421cf50ab742cddc89301eda4c3932caf0232778ec5b069bcf9552c0b55b96128f929b57ef312eea5cc8969b4f879db994d213c5729dd4be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e58fc7e716cb83a977624c83ac24ff4797ac763943f151e2bc26a302d308b12c18f8036302315e3781401730f8474f6665510aaa8edb237d471c71f19ac251e2addc3e23af20b4591a7a8e209cc23b6ec1c3b0f2e7195936e76393;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h243ac968fff7f5157f8f0f9c7d1d3edc1eb05dd2fa1fd3f8dfc515e5b2b9fa041aa32471399eb3cd7889f0ca944204b39ce6ae4f99054bbc9ddd1c4013229fe9bca64c8504805c726dbe00556cb83f13f87c992e1509f57e84df9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd7ac75bc609eed12542d4350c28c0acb653480dbce3ee78e7b3ba304eaf97413dfddca9ab80fd0d42a66f25741e9e4f460f882d491faa7e157349efdd6407c6ced952ed685436addb67a6bc00705beab8a3276b95adc9f162114c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf14f987862754c0b840803046d9b3df47738487d94f972cb04fcb04b4967b735b203ee76ba3ab7aed9a66d6e4903ce985b7bf5b3436aa7e416a80025a24491e359c97a1d4577f313331ff4f3150fa87763ae2b0e66f25b2c6813d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h641f91a71a3e5d15cab135035885d1435e04e9f58a207df92b762629e22641340599ef753ffa2c89b40c16414bae24ec4527102fcb45bebbe77f71c91114cd38914c46fc0d0f3ab8ae0868b8591d44d7f26224cd3d6982db175d57;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae18cde6f795f8269008bd24f2e856b8eadbcfb0c71714b61947d1705d3de7f19134ee61d2056a6a9ffcfff0ca67a6e509508a4b7490dba9576dbb266eaa8a11b3229edb8781b3e637ababb292802515908c80cb5f41d27d39dbf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa8c1e2fbcd57e9aaba7c6006ba0fe860aea43d23368a8e5974de5e668ea5ff85fee1f83bb97578f45b865437c2c08f44b4a957dca14e0ce7deb54ba48d1b7b0a107e9c678ca08aeb60cac3a4a67e391f2813788adae41bb408d90;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a793d01a8416fc0748ac095ba36f3778874d7d66416802e7b2a8db591547d8242a8708cded17a821ee3b01515b434c9dd554e5de8615e5d44ea9686aa98276caf6848e155287adf7c6b45e766ba1a15fc3a146ce0c09dd971dda8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h863868bee5b84e1b2e8bb2f782ef05d437c2c1d32d0d0f7b076441f867f18c74a9d0b757134b59553d6c899b0142f3ea967bdb964a5c805d21bb0c39c2b4a0c0d71ce3a5951cace9d57233ddafadbad7b8b8b9ea31d649d9540c23;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1379235393d777c1adf2f31276db2a9a8d94f6d1cdbccf738f2a1709d434aeddb87ccfdf136172c37aa84042403392f64401de432a7748b46764580834f77f78468a7573f49eaa6b5045e5e3361bc002ff7d004527d81b0e2b9c07c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166efa07a1a960ee164582092971e5b3abfe2cde673474018bbde38c14360cff9f3d92b0b64bc0ad09026bbbe2d45f51a892fb4b74fffd84b4a1b21bf8d28f4ce686c25baea65d75543355f7604c872491007e8615978e23912da81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1732a5b33de52898daf8d67069738bf85f2bbe9d69a8ae5a39113a9b90a376d37446e97a99805d7c0de70e5256c46f84536b726679e544246af4b0ca956b2b15f74870950d05cd1f01b7269f5ed798552d00c76f794c21c89fd5b32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75b568858800b8ae28dc18498664856f7cf3cf05a6189f7add72b7f3431ff7302e7817e66a28bb6a343632382955f32d4ceff36f1f2c2ae9a7a8cc2393933d95dc4d63deb223f755f89cc9cf55a9c764725f059525a3e8f816f68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1d1a05184f99b52a1293c8a9dd0020fb84cff89b9c38ce9d1451758e2700ffd1ab742153eb9f448b91c4ffb27cd41f1f31726bcbbcb6ccc972ce96d1052ed03ca9cdbea524a3e596033168ee8a77408bbc328a5ea2a618d638da5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d08d73b79dcf49014168b367c47c85bf77b042d46298c105dc0d65b28d280fbaaa36162e859f1d2d5cf8b5da9de068995a37ef3694987b40fc592080ec6ad4593ab65a8d25bad6f38a77b7285e20649f5e7f874b305b1c3ecf411;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133e15e86cbdeb9d8da736ade88f5896632cb7a6f074e478afd93274100b8b6209c7643b23aaa681edb99683c60de4948773675dc4cfbbb413811bfac34f69385292810390ee5680de35cb9bceccaa9c68bd31a4220bb94552f05d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9fee9167aa866cb2d4ef450759a7b6aab0423d6d2650fa4c0748ecd3adaee592757ca5ff6418381e19fc2226359b3f54504e465cf0d5d89d0243a082645a90693948ea90478dfc04ceec9178bc8cb39d4169260e0fc356e5a9ba7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f3c96551bc35f6649faa9d1bf140d4ba463962210b5767317193a35ab68349f785321028758fad38e51c8b50ac652c8fdd3618baf8393430230915dd6896fb2b1881e1a7c1c71f2d32f0ef13e799f64ac74f1bd4afb4687533cdf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ead00bdc80ce5f88ad59c9f2f246b2bd0b2e35d2b2b3f1b0199302dccf936711f8e6ab25b9a1b35c02e770cf24c58f73c36bb3176cb250e3483fc9599db683cf96a6c33a27ceeeaca39a1ba225181ebec1503a27752499ab00fe2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h756534c8a470468b42756f8d5f0596a7801b7cf876406fc9218f5473cd756ba39c26e0050dbf14061e2b4db2d711e2c55fc88fbc90db91201d048cc16260db4c6566df45f7a3f15c2529cb734d08e98f5ab023980df05133e7aa40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c844bd77ecde463e1ef4178ce953f862ce88a59b5c19298882cdcff1682bf55f858a322e54f1993934537c1e4331bddd7bf8bb3db4d1657c838c26808b192c09cf167063971665a061e11ee830e209c8bf2cc0bbdcbb5b7b018b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50f3b14d224a24578db7c1e351ebd43d9356d5ade38f8ba0510f4b6c6d4df49eafae0237e121f743d026888355860d0707789c84a8565f1963434b11be9c0da780e24a6d34d96b4b15e759c1f881c6ce243ca4b7861cedfcd44c5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b25970324f86335db36040ea357a17ed254f4a1a6820f224d35b62202954d5166358346520cbb0581c3ca50529ad1fd52c3a2279ce2f62ba0ceedc4a548ac9c22ca7824d9f50056b25110d56239a6df94227a6e9c1139ff9e3945;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ff3093201ae1b9877dd3b9431f72a8af8cd82e5bbcc1f933cfdba7cbd8cf6d32fb57251f8e95e822274b0d2cccd317d093420cab66883214a8ee55668015d7cd5210a61a5658d89fc95ce3a45d86986131c953ba8125795d186;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47b6709149f1f1ac075a81d9960f3fa0a53cf41dbf9581fca2014ed7517204e03efb197a447b7e65e21abeb81bd90039d6380f753cdca7a34356d82a8cbf6f531debd0335bbe19708d5e1b26d73e0059537e131fb73c87c5146081;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1685f93c79630cd8e5400dcb2f22e550cf7b9dc00c0218f5425cbfb31e59f4ace89f1ecd835700464dd3492b3d9a50c34003be8184a0078a0db1d21ef7b8ec1d40cf335412f184ed635714c0010123e1ccd5cd052f72132f29bdd7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5fb6a57b7d6666453a92653c5d3c2374bb4a59081a1b2064df789e0f0de203035509ab89346de23b9595887d053c681890d4f513e204aae8b976c61fe04a3590b8eed3022de45ff2ab87a39896f7fbe587b8b4a963ff7d769c749;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44fba15f12025ad36da554125eb51245e67767918b71dd958881b621a2468bd46fff280997ead1309019e4021af8bb994c3afd1fbf865496b5f7fe20ded3aec3a1c78d358b2d257f1a7f4a6bf50f668c0a5a3e599fa8a439378fce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f31a5624383fae3eaf0c643203dfbdf26227df2a44b6505592b6405b9fbe8297a60508b936f6fc4673f35158cacb7738186cda66e82da1271d5b30cd0e23fc546995b8bc90457f49aed30807c48c97d7e953804f23b39671ebd47a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd0a2627e69b3df1e169b8e72aea2b8df5b7796a3d63c873a40441811d70b55a8937b670cd6cf90d4d9d56894294ee0e6932a7444bef9897adc383aae1f05316281a4288c5afc71e847ada50ad963ab0847f0eda9e32f2e9464360;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ee0608c996290a781cb047782b5c04cc10706dd27186b7f466b455ac8f70a05587eb0ae907f7e2d2e52d13112a03586ccc33d0db55501bfbc205be71481fa2f463e129b0bcd6d8a99c31f58f04a66fff3ffef58b85ce7831f9425;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ede36fb69b10999cad8cd52574984e31bb3dad33044e3e51986e329a6d1406fcba1f38a9394eeed4b8b05896c9ea34887c60c43e8b7596fdfe043ed267dc01d20ce472c7321bae42d203e7bb7e5caad287ac31f1b09d8a3625b66c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91c99f4780f8bf0495a90162a21e9710bc51df942e5101f6ec318290ba632e62edccc395e4a9783ce59ecb2ae88639b230835b7fe38a2cd9c2854f1b5154e4ed5732756479a81784daecbbfb1670cdc0f257733f45bef3c35aeaa2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1c413165bbfd38c0ba6412bf96d398584da1506a966ec410ea4de511966e1bfbc4e54a76853b87953d4fe19789239ec79097c6ea37bd6dcae75b9fb2a46da2e8b1fef99edb53c7eed45591f3cfa04cbf7af1a91d925a2852f3e83;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4295335ff6b08a09e20cd359db67bf3f78d4acac73bfefa322aa279ab4e85a1777b3c38472440eefabbe97e5fd870744d26f50c97c874dc066a4553ed63c193e80474f37b015eb9666d2c6fad33c6254da1c7d8f4931caf333acc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd53eca2624d51e720be1534928f2220e9300120cac6f5cea754b0632a5919443e7d1f2837f145d6938a0bf7935c8c7d8ee6cd27178d35088bdd5b909a31bd85810f165656dadb3bb14e65bb2772d9be62d73465b3081e9b029434a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43401472fe097bd1ecf5399fe52b46364cbdcc24f496126d65acd520902e3e912a4191d6067b0bd6ecf3fbf1690c864fa3f5293fbbb9204c7a5a51517ad6f8942001958b742a03314699b530113303dc6d4475ea97a5cd3d41d6d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1816774f99c7a74ec3035a865457a41a0eb267391f76298a4a81531af5a00a5e5f06b1abb2cbb5f52f9fb27de0937151cbe1d5fc973f9fbc3aaa4cffc593e9ad32621425741f0db3c7735d735b567c4b979a735d73cb1ed0203c87;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f406b3e4e978d9996de9a790c92885957ba6b0c0a1af2faf798b53568182baac561afd67c6aebad5cbda860f827b5ed2457eac761a07aa29eb145e888a53776d8b68483268ca041ac9900259f826e32cc7b915056f95ece86d86c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f9804bcdba04afb4431f0d6e00bef53567d6add8765ca6e1b584af440781a58a1010de5fa37e0e5a9993917b5a9eb3c53ca7226933da18e912d88ce821c2c00f1cd5e5eff56fe68df328dfe053bb0ead9255a2ab5d8062610dc94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9b4043a1a07d7f12fa123888e5dd4e1215815b110960f511be30b53e2cb1df1f378deffa27d8b77cac2f1384cb0f5c3641875f8ba0df209a006a8efb8ceff6db1aae56fa06955460fa2b0e4f44cff263d40891b4b1e37311319dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8ef36c825e32503f39e43a3d29b478faae831b7afcaf73d57cfdb10d80bdc2f82c275023199a281f3f22853c39e10c9b35cdd47d057cdcdd05cdb38712cdbee9a0287fc8222fc33a64f799b688ccdfbf2f4f2948ad04040c62b8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180b88b9e53010d4fc538e0c12f02d4a0694948bf5082e146ce0196d3ae5bfa7791c3a8ebdf1c19e6bfb7bedaa7f2bef26f7bffbfdd0af199bd5da77cfac0111997140562697b689d5a948136f291180c580fe29529fb2c1de5cca0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83354943f292bd961d96c736ca2a3d3bccdf6772295a708bb8e0855da872d4873c717aeba3a28d48e5d5722e891539f0a9467b8c650fc98a36d673da170fa0e2a36d8f196a700cffbfb5e3dba5cce2966805c2333e34a9bd1ba5dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h679df2098c9ec0c93f894069f30402cace2d724361dab6d1a20e2fdab793c5fe4a15ed8b8a476f9a379398d9ac6468a9c992bd44c28c5bfcbfe0156d593cb53b6930d801cd86d48e9aa60ff9674760ff9d82ae327cfde0082fa10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4998381aa72fba21b929968aa2e0da8eddc7f8be2dc100f535f56c17ee30bc43e3f3d0325b105032a084de29fc3efacbe5d1346e9bee8bc6d5d6dc860a2704c4c07495b2ee0466e08acf435e4f9a883ba2269a35c6cac9366a244;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ba1381dacbc13fcda8f6f1c6bfa89bfe9e2892b0bb140d3c9b64637559b4c873483fcfcb9635b1d526b56d665965a9396cf1c2d3bc05a81693eccbb291379142c1bcbaecf902ee3bf286bb6e0205a37dd9894185b93e189d7a468;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f9a7f2699f0a0c235fa3ad123eca820517183a930b1ce348543a3308f48c0abac9f42100b67d40d4d38bad51d46b4fafbc8d07e237cd83ae4a48103e0ffffe4565cab09ee82df31ca446ebd46c8db594c8a451c15e3ebe115498b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd8c93247d55a067b9b06d67270e18e597a3780fc4a20d5daad927378b97e74f6ab1f91018a2132954020d2665c4b1fa0f2beed7bcd329df05795451ab165b7998b0b4c654560902d79095bf24f4fd4c9ed0b465d8cb3bc95f8458;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168e581b3e573f8f730b4d3f0553b59b9a23b4b7233ecee60e63d84b44e154a882dfb91394786f89108044e4fc4dcc2a84daa6add6fa206db0a7607ffb54e00469b1fef2c13826be5c15ec532f575fcc6f8191a89560753ef580ba7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf70553f4a15325f3c5e55378195971713af5090fc90587df2dc6ab9b5b0413c145c3698db60fe43a1ba19ba8b3196ff4a095572b19d84d16c75f52c0a4d90ff20e433624189edf4a22b952bd7014a7c7cb7e31f50bce8636ddfdf7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6712045b2df9e81d50997db154ad5174eb6471d0a1175076c54bf39ba1ceea3c5b1cfc306b0a51098a98ad86694330312d5e641add1042d9b1dd34064ded05cf06a1420edcfea2b296030d52604b09b98c7523474ee1dbefd6d971;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1ef4060b56ee63a8582d7b5bc303aa1d2506fd07a41da41b67abcd277f7fa862aa750f033ed02d1a0b5e48258b2a3913d880b4ced7938d3003f442313e1dcf99d378786b1616e26c7c09d9b8f35551fdc62e7e68869b0c9df5ec7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1230aea63f3f993efe3d8a58864053c9382d1c9cdcea5f6d1db6fc16cd22245083f194d99960d02e7f4443a486ce252dc8960575731f9d78e04541d365d0acd149dbcbf1003948e98fd110adad4b8eefebd014b949865194e234b2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd69c2d779a7aab65a4dc0a81a795f4e0130a719b3a701640391bc3f8e9c7f702c079e3dd05f3000253c0db05d5ce6a62bfcc7c21add70b8bea61d1eeafc54b99e184fba72d6cfaad58d7eec204e6048f1c64ae1f66cf823d06eab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a8c0420af611cf4b7f6200e26db0fc33a96ccc17b459e64eac41237da4e1040f1be24207591d43344235416f4adca5d7b0cdbb03b48ce30378039c10a4eec388a94867155f9dfd2395fe2819b03c8a43c693e413dceda32399074a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15deaeb203e8903fb726f84550638f569831879988d1cfeed98a1e9c2a2159f28b87d4b3bc35eb1ea2ac52b78ec36c3299dba199838ac74aa84562d38de138f3effad1130aab3eea17f8ce44f74513fe7d9dd6502f618a15d815bee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fb33d954cef305f8cce6483b07f1ed1410c4958daf9b3d521ef35d47500a743de7006d84de7ab3160c25171df0b001433fd5d7f7000ec94ba41f931c5b4d9308ce05f9f074d3d3e3c6edfbf6dd3664c0b80574f41a6f55b475da6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71fb5a4001ebb7a9be1cad44bee84bbda5e69503c789443254811c831d7f4f715a6df1da61c6c9b54c88d1223690315c2436bfc3aa8993f2a887bf83258f82157bee938dc7102289ded91ae27c104a4bdb79e2eff0458236c41ec6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114264fc621b6c80c6aa83526bba2bf92f6f1e93311e1e1af81deca46bc6aabeadbb8cf7ba34249fc8c1af746aebf602a28200fe20dca797e2b711d39d77141ca6aa8cc77d0e9f751b16ed881026e42443fe5cd41adb4c3e234227d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc417059ab8b41f08ae805f6a0c8a481464e942419cf7e4e17b41192207af507184e186c8f9202c43f4541f1ad3cfedb588c28216ece6f15b3af41e52cb17444604c154f93a2d249313cc14b32079b9ec6d367353a3ec020cd961f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4808030315518e824de2ec781200cefddbb9111920e9e94251c7c53d621e4f90711c74984eea109a25a9bc54204c2a49a9083ff54b465f6e23ad5f4d7d18989146d9290d50523f18a46039458b11415b1c3db1bd509ef20fa4c280;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d71f7cd9eb008650e5f3db978d4146912a4a9c28bb63d6db5eeb3019e993661277d51363bb0c6920623a34ae98a2a13ca17be42ca1097aa4ed43160ca27b4ce679319281e79fd66e06be077b30fd39b5bf5a05d0a3a05f4777f34a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbae8d34fdf81cc405ce54807f0f899f35ed898e1548de659c75627c15aa585857e4e515e2722be2215d1dd6e9266b7a1682c01b4db5024ea9b07070b300cf192c0ef2b574a680ff898149f1933f6e6572f2db61a63a345ef98ec7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147b299b5f59fb799d9da193a9b412b42771b468c5c8f6a765eb86ef2a2f2a51f082c19108b40bdccb8ea65f8b2f6a79cf7465ef5c12367d133abd0116709506872bbb5ab6b4fffe80ecfa07d0a3ba6d712ae78eeab7806710340e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136d1f541132767c962793685f0287927a61a22a8bde4a3eca6f51e65462f3adac9aeca4c6756dc4b442e657ce7b17da0e919bb47e295e718976a4854eae8911413545c15a3fe71ebc720cd425a5abe00b44d2c5518d7267e02f9b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da90819f55b8aec527a22881874fa59ca77c2e982d45a2b0bfb59e584b1ca3767526e63a42bf31793a2839e586a14389f8679ed5f278a48d111c2bf1240253906dbc0f8a7ed8b75f3a4fa4f5e88b1cad0e2579d6f6514f7405a603;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afb11ad34bd426fb21842995dd25c4ecbc6fcf0c49758dc5795f1b4ec77d0abfd3709b6820a30c1cd3201c5e5b0a957ff7e8073f457240fed413ffddf284bf0fba3ec41f38b4e28bb38bc167be215f21d4649b59a07ef0fd963507;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18629290c6c0b7bc1ac57a194f8cc8d694e90f83852df2744bcd6d59a8a89941cd9258961b6af531abd29d9d1df8cf191fadded021fa4631bae7f91aa44b1bb8fe1493876a1368ab70fbe2b712a73c03c16fad06091f97c9d54a127;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a3e42877652436eb4e5a4fb2d5fdfffa3da6bc4935c78f52e5a5d35d414574169a7c15bedbb736e0f2a0c090a344732c67616369e269b16777e837377aa972fed6a94c98b48545b77073ac1e5e2fda772125453f0b082efb8ccc0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc542db14cd600e99084d83bbf4577dd2865a2ea61556f90ccd8e544933a6e5995038c29487d4e584895d4bc197c4e49966ecb5423a19f238f2f1410fdd8a8d28006991b9c01a20c829c2163a6b2be9d3da077f9956005fc4cd8417;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd92b6aabc9bb0f47d1ad9d1711e700c79dfc6ae66187e01fdf70e7bb7ffeca263e3d1c365dde9cd8a3b8157ff01e10c07a15a088de7ea062bb458382fb275478db7b22b1b72d821424f466615fdf55ed9e8e7285975ca1fca24162;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0b5e5a4f0f3e20944a2012794c0eec2a7898253511b0a9ff4c08d710c9de4ea4c9ac495de052e5b96246c5bc68514408c06b4da265c11bd169070d1e67d3ad220e7fac70c5e77ca8170d7691f4912f5b70eba5942ce2621569148;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7cdc04627008704217b35124de1e0add584a386bac91ae0c03158464b6eca6bda9b4338d810080d77e7b50c6b53ac5ba07583447a90c12cb199b5c9ca2f7428b3a5ef6d1a7350c168e5f52654eb9edcb781c1dcfa30f1c4b8ee86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3382ef1ba19bf049bfa5a06ef37c34c8b3835f4b334a3cb3b7374a9904ca389411d9af2ac4d95f9462782ff63f92a823279ca93f6b4ddcbe6d86038e7efa3ab8a7cbdd0e3d36b5d1be478cb9381e6f12093ec1425156a24307cd40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcaf72ce438a33e1791a1135cf1e764a8f91000e48b86ff638e68c62bc464cac365aabef4b402a2993c90ff6a526e1b3ed74137144f6c85875ed4b4008ef247cd7f9bd24c5e764206688d48ad785f6b6bbdcab41792aecb119206cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5f04216fde15decae0c8ff7aac8fa888ecdfdcd65d524f0d59376449465a98f7133c33ed8da02ba037ae7f4f8e75d4ef48719c39277d46493b58421b530baa6afad72f488d30f0a5952cdcbea1f083e8dc9a509a6f0e41273eee4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8eba909a82fa48e4d268be95266dc76e6045c5dbfe56c91f3a7b476860a0b4d68c943892f22e3ca6e6b07aca6e1dd8608e29bf70c4407184bba8d996758569d3f97cdc5df6fbf615580d90fa2bcc1c8ec0f9b59aaea1df26032c8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e05ce25774c5634592947591ae6ec51dc1f38fc05d6550e9a8b828b41f6f97b603fbcf7b9c3881bdba7a633ef3113c9bac2f70f9ff1a9874a98062c76ada7d95e4f24d408b7a20ec42456eed2c547a424d3ffa3795f79fb59a2df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8b6ceb07003efeaa9e6bf4a4a46cb6bdccf9b76305cbd182944150d62a2544260d58a47546c31487c6067d41ac8db9ec746329c0f4e28cf7d1e4d05f4cbe803980566717ddca7eefe3617b62bd14a052e0867a831e742d7d2a305;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10139062702b8c764ade23578b5ac2b35e126c094ba4da53d325d41b0ae65f05196bf752e63ce9ab45de47979de61fd9803be340bfef0c5d2f7b0c20f40595d67e6ca2072ea761966fd71bd9a27bdddc6cefeec19b5df98c14fae8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1792652f2aeb5f345363d63cdfb26376915ede8481708302803198b7dd355de443c0693efa9106c3b36c12ac5f0d7025a7a4ea6bc5c84492a3f704254630b11a67017b34647459d4295c2203bdf799fac4bcc06f9a73f1c63472073;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10154f1d115c59c4d631e1edcf909bd916fb039d19d3dd64ee709c552fc43228da9f64898b3ed6c3fae7e1e740b3e75975f905deccdbed32b002ed6ed1f75c10cc7d370975230657038ed46860cae774081de8187d86c4af73b7f99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7939ba4bcaf97c47b5617329b132d44b4e0eede3816a4a748ac25d2433b3cc541afe2149bf22bb687c7c7c61d9cb9e524955c4de273f7f22f0f3d34e562d839107a2bb330fbcbcd146d3c2515638c8e583e04d437345354dbb9af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e17a32fb899b15c4140d5186acbe84811dc2772b4e6437b51f54d37c86b69218b0441a414ffb08b54290659e92dee7d0e0d211286abb39e9fdf0768ce57a08776b2d3c95be8be0658d3c206cf4a8866940d64583b75a0286f810e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb3cf387aa43bd43b6d20389636fdae06c880674e3b1ce2ed5464f8ee84bca4c3ef14cc151263076fcd9596aab83eabc058243224e4ee014cb427cebc811d34e1dfee83e208f9e0cab52565867c3643c73911f1445e55b5790cbd4;
        #1
        $finish();
    end
endmodule
