module testbench();
    reg [30:0] src0;
    reg [30:0] src1;
    reg [30:0] src2;
    reg [30:0] src3;
    reg [30:0] src4;
    reg [30:0] src5;
    reg [30:0] src6;
    reg [30:0] src7;
    reg [30:0] src8;
    reg [30:0] src9;
    reg [30:0] src10;
    reg [30:0] src11;
    reg [30:0] src12;
    reg [30:0] src13;
    reg [30:0] src14;
    reg [30:0] src15;
    reg [30:0] src16;
    reg [30:0] src17;
    reg [30:0] src18;
    reg [30:0] src19;
    reg [30:0] src20;
    reg [30:0] src21;
    reg [30:0] src22;
    reg [30:0] src23;
    reg [30:0] src24;
    reg [30:0] src25;
    reg [30:0] src26;
    reg [30:0] src27;
    reg [30:0] src28;
    reg [30:0] src29;
    reg [30:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2722063b0cadc769860ad1675421256ed51eae6cf11e2848a9e2ad3585027b56cdd4204d65449b56cae230e260da0c05af7e64e36da7d5b7f6e8ca870d7276447dfda015ad7fc5bd1c4eab9ee53649667d815d44da4f485dbf49e4ad27dcc14dc83f678d5af0c7120b9b747039849920eea1ab684a7ad16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha95cfe4268568de73706769b7b5746ba0d636bda6e897a90e2ff24d37aafa7cc2cd86eef850626bf54c6c077e0f8df8661f2ca11345983801021ecf70777d308e1b5a3f5539a9c11ae651de0e87709e007a8f3f20425e349ea4c3bd9005c68f266b87658e2cbffce81dfeb962a91843fb269e518a2f6c6a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1590845e87f777fb34b1141cd73fddd7758967220df3454616a153c264ed4336d8a4227e1ab236f528013a3dce9d1351987c911c96e13111e92342aa3ba66144443a648d7e6de787b712c936882bbad08333962076b54dbb6296e1e347e9546fb81863d12e4c3194fbd09cff73c851de426517eedfea524c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9b3a665858d9b009d35894b40a8598347c1cd2adddd62ff224f6c15d1a1ad645c54887e46c0e314ad43812226bdea5a1e857bb656510f99943833798e7e36b16e34da39f5539352fc2d0935db32eebd61cfe654c7fb73fe09af65ae2415e85e20eda99f4efacb739dcfa7cdee766fcc1d55176889faed43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h55e2c3351b3278598df370248b341fc76ccec293da6a478a498acbe4f913ec945306437e194ece9f137ff77845ddb7d93060a8286fddb57bbcf6bd1e838a5b150ba3aa95f917d1c20ed15bb753003aa3be943a76070dc16b2dcf141e154746a43a7aba28cc72ab3b7d92469cf4174def83946ee0461b7250;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a14a1842458d7dd103a36c787f40367fa4b9f0d86a5c3b9e33f1f2ddb9071db65f21844fc2f2ea1b450fa5f4a25f867f6162892128ad564944edfe53f4779628f7fc1eedf2a89b5ca8f4b9a86d7db1e60bf6d5ecd9519018466137683268be0e90de9ef438300e7d68cf0d59daa5bcd265935d072d18a01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15197fd4253465e97ceb8b2a8342f0fe315ece8a35d98a852d52426afa4523216a71ada8e0b017edf117660c24fe15d2c48e32edc41cf705de52fd0e20966e502268f531ffe9f3c0ff8978aeb501c584cc79fbe6a0f7ecf4856517182b459a26ca3d12b5cc895fadfa2db59f59df68f5076d2785f707af305;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da4251b2f01951faec6ec10db8246b66b848bf6993fe285d196e05b317c19bcc12e6b33e3535f1d70acac8572cfae9a6ea6a1cffb6077569531298e4db7cd5ee2e31ce5d599269c133961effd6db7ccc01caccfb953b726d6f7cf78e0d2264a5584b2ae55e2792edabbd5048627fdb3b7a30ac8a44b36107;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb8e1e06d798c066f6d2859dfc19ce781280b9001645308180df8c1a67b4cd4e076ad8e8237e0973dbaae8ac95d7ab6c04a48110aec57d94d96609278487fd76948c919bee0bce20fd511312259f8655b7a00ffe5a2fdff1c41f843be84fb56a3e6d3bc5aaa2da3f18289797b134a6f83f5f5c5d0a3fce41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b41bdaea98eadd3582f354a0bd24b8d807dd85e98f70ff211deeb531fd5e26e252d3585797b8afd39058717f4744b4817390217b3bcf3920f6965bd58a2fab92a4be36eb8d5188ce82c0f81e0a61470113c7a361a5bbd5da60ee9406481d7bbb74bf55d36108ead4cc7d6b7a80fcefdd48cd9e596d414def;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he126d21eb56b572546d6fa32d6abfd8fb2241d9a4e7dce637a15f08d87d1a4a250826f814a0b8d4b33bed17e76a2f30b40eec3e26b615f1ba0543f81ce980b1e61ff61918cfd82e0f412b90d31e7ce94c8d0e416bbc7682e5a5c3da3f25906a270f8b53e865d507c9713bf0adcf874279f5070af730b148a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7670b4ed739edbbcdfda198f6301786d3890bbb94a48702dc626858074bf3e7e167485fa2307bdd82388007fa1c4765d0c2e66376d99447a175b9fc3afb43611d2db8f3c95d441471a87ea7ec18ea655a2af7cb63e47fcd805b9a8f1b3376fd3bab4c7f4f83f8b43d925892b827f5ed1895c2e5016485280;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1daa96594eda2eba6caf787db8fe91981e29fcaec8ff58a9ff383eeeb9285ca89b8f96c30a8b4388e616c4ed244a4ad6e7b204946f4359935ca28233b98287e1efa888b20eab75a2d9cc42c84b81431dba25196b7df9ee192d01c722033552904921bf2ba9b1347e656044acc1a11d7aa50cb427bfc05f1de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7f17f210cd83c0cfdd8456e2e674319aec6340485e67fdec84ccbd28004e4849aa558774b6c5b678ebad683704c3b1d04f99f783337df871e37cdc7b8e80659fdc18a4ffede2287e24972f424e822cdd68e3044e1f3b84b51bf5ffa56943145b958ec7b9614a7d9b207e15e4e3fa7b1e93f14967c991a8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22f73e23c56f1b0f430975931f5e61af64eff3c024f643f46f10670ca307462639f0c83e427134ebe42c6cb22d16296966e6cdf18ab8108d11c035ad27c2282cef850e86348aa13260f1dcc1315e9e53b6b7175ea0bcf97fb0c9aaa245740cb044b787969bfa0cf3313df711ba833bae2681d690ee3baf6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae6a8d601c26721308a34109738748a3e17913233dc850aadad78e9bac544485e151945781f0081d31b25538ed693bb5a249f68cd09ab19fb19273bdb331ea4129163bc7f2e6855df93f7ab4cb539016bd65fef5ad5be421af584f547e45c90bcbe25458639244043c2d6e67db187d37ce768352a16f3135;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d8fe54eb52da1d30357ce8816e3153929caafa26b53a5cc6f9bb0a5e083da6e87e0d060e79e695c588122bd0b653dcf26d3e7c76b859782aed33a415f8f17c2e2945c8a3c6c7b966ae8a07599a9217806568c38b15fe7a9915d1c3eb000b68ffffccc4a3dbc64b3a54338f25c1a995ec478738bcdabf26f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1140fdd1e14e0165ee313aad6f4ecc9b8f698e08b8d35956b830d1e474806e99224d94447b9a647d5de642ad0892629026d0560d45dd987dfa76c2f98cc4b4fc77c9374386303f54cec1e1f128eefc28de4a3f789ea7897eeb61d9d90ba60f70b602b98fd6cb876950074e2f3cb221b416e406a3e25ef15c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8df33f09926b112def190ac1413a4c5489ca641693909cb7d0066fdc74a6da55f891a5287df3a5825b2a55acb61537b6ede1703da4dafc52515717790c9305fdc2d2d1913f86638114e86919dece97ec3c14f173015270b7233e904ddf8c6bee1b7314711072078ffe065ba559afc84184f46b61cd06c75d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c1c1e832879ff979f9a347da7c4bee8b42351d441ff1807724ab23a5c5359c226b98a702a0beabd241e5f2ac52e89c6929ea55a9394b956f1df96518bff365c8271cd27505052d535e1b1c3b5d1db54bfbb03ff5129ab4321dcefb08875906485b8c1f1d8c896fb2faa9349dfb6f1abd8689ffb2212dcb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197f8b45c7b37170bae62ce2a0ccea44f9c5154703dc42f49179a081fb6ddf2d0c92abe806158a651903d2bf02e2b824b0ff1e07e98cd1fa9dcae8386525ff8e82ffd440d4d8789b2680e35e2030956592d65be793c0cd5ae9e1eaedbc362b251a9503641f65485b25b4a4b1b3accd8444c17bf301b7a53b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h649ac93dc3f792b649ab2f48c77e833ba0766c3cf32fe0c75b8b371326dd1bfaa602a74dea9b337513fced369b67e5630967821247ebd8577c87cfb0ed9ee1d1bc89e0b395adba3ad7c127b836ce499ba33f9cebec488ddb4806a8e0e3b8ca1873eeea9542d090e6e5b27226edecdabe7fb20abc3f4d20c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6496aa021a4a22aa01b4140c51505d30e513f714cf5bab697ed298ceab819493f700b0962c9195bb38b95ded2597c26175770f8a73f3d8670aaa76fb499040718979140c0a5d10c8f167cc3c2ce4bed23619edd343f1bfdc8c996146ea79bf1a3faf8e33613f3f6273dc40708f683896e72a0e4c03c28c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90d4f984c79e52e0e363aa84ca94edf7fcdd9dcfd56dbea5b090f737ad50128f5f2d603b38dd89076f74de93a45d5297e0a7a4c7d0d8a360ec2ba9d6061b60a62ec47808310f34c38de37302f89864f67f1e7c1789cbb5d4df18015b4edaf53c7340ee47a3894150527ffcaaddd17793ef910baea898800f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae849d480f669596cb3f389b8bf9b469b9faaa72061494092c5d2f60b2f362287dff1688bb8307e5d321be2f5a81f10e32fbf61c7c42f5959479d2db065f8f56fa6025cac381bc10719c39b61b7617f202509e695b5ddc02a63b051bb6d5ad6f8190e9b5a1bd1cb62887b32e2aef2c4abbf4ab26b27905cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5a4b100dd6ac2c8e9d6fd0ed36b37e0ba4a5b36c35d4c4fe5860d1b8fb1c766ea1776193a5fb1beab07194d61f58cda45082be8239f9372d398ebba87459a1e65ad23d84a3332ebc53d4ebcc782bb146f3f9125d105f269dcf9b400e1c8377f938a6291534a5462789755ec580e363b33eb1e74d4897ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183d1a4aaaa72d8f5572e3e0b852829dd48ef55ec8c69c0f44f28c570cf6977309ceaaa1b5843669233908d9ae16c3b0d0017b889de6d8f831f2c54160227e629f75de2c528121ea8a70ed270ccf716b129279a840902cb955e9bf3976feafc50e8f08a7972cc9d9fd6dedb4ee3c29a9da0b2d257c4a719f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a1ce7648fcc34689df17ffccb689fb1b459d8af56c0d478f20b6ad6cbf4e6a7ddd526704766a899c87850c6d014c3a62733a0124bb77daf52573d2519caf9b48a314d6076d0c7c0bc42b72aa46d551277e7566e4c1fa003f4ba623b4f1c0e7b0254b313162e677cbcaa5b1411339eb77c23cb3c085e055e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6efb1de89a368423b7a1af3910baa3cfc0426ff2e8f169cc6da79fdf70975c22e46e058eb20366d50d7b947d43fbbfff27b0a56448cfb187e9900f9b0b7fa75947e5998b5cd9d1655c8bc02e54fe13e568deeff84c5a3bc57c86d7dc27bcdf0780310db24c78a7557bd005c3dad7e5987efdd1ef08693de7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h280be38909aa59bbbe6f055fd0fb154b05bc098d38a58b4020eb32dffe38d90671114203afa3369293371c01ef6a80207c82c4a1918f7e9d3b377a7b401b5a9adba69295dd43752c4fc33b14414796a99adf7813c20cc9982453c5c77be7ce7c8926075b0ad2d8710820c4ac9c576162e9cebdacf17e434d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c996a50d90156a082b4f6a619f4b75f962ca31790dac8a0752277e65efc3d1a6f9219b7b8431b78559b4d3c07f8398ba1bdb7f361c893340c8b59e9fb9ccb745cfe22eb9dfa8df1074e079ec758d066304f54f8b4fb8caef02fab1ee35a17b75b4dc811ab2013d5ae7bfc760fa09747a01f0eb4824fcc144;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f20a0fb20d2b8c6417007ff1b6f8165b6251a294598199b505c5baafb8fe5bba7acc78e49187d6f9368eb47efa0d14a3e04ee33dfe266fbc2233af98379f5473062f082994c5bb3f8830b53c566ddcb7cc8a9818857e415ac2401e7de78084ce5625e77fe5f14b307f9ceb432c7752346b12853f5852eadb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16fdb974ee86620c6184dc2fb62997ead209969bba9efc70c9fec12c6538428fb2cd99b850de58887db79b62bdb00ace3cf27944c58d5ab5cc6613e5e219c0b64cfc85ea4f58f37399e1751e2bcff36788f105cb01cbb2ab214d82f064a21355bcf2e57a6b867e16b941fbbbd2c189408d969581b83f635fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0fc45d3626fa3508a2ba3c34fec2e04d4a1bb30f91af49c02e3f84b8fc4a00c7c8ee8e21609dedfd1a6d6b3dd08ed8188f72ad162ca4e6e73b99b95b891f10655d6b69d47d397607347cdd03a0789f191e3f6ebc0eb58d0424513762cc82ac55cc8970fc6154a8cfc5d7210c9a99a4573dd1fc4f92c7839;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118f250573c0d955028113ae12113d425e6221d142c351938fb4cee17d1036f334dddc0b8e84d21b673d7b8d75af1fd0f3794efcce97a64f2d6392c116893a232c15b02bc26abecb64d5e22426d082bb59e5f30ec720774666fd20ab284bbc6453017c6208c38e133d126d627bb5e4020dc2468465b697ec2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h947adfb6f8b6306298c6c3b8a0e85aaf0b575bca50736589e9ab0d24f53cb089f2444d5e464f76443947ae549b70f5cd2363a398893274056c1d936b1b596787a90683069838266f88ac39467ac40592531a96ef01e546bab15e06f588ebcb5538cfa95e26f360618ef7269e673d6e7cbefe5e9758094193;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71ae4b760d4bbf71e0835dbfeeed98beeaeb48b0900e0eba2de327a4c5eb2a1eed30922516ec129446cff5248823095cabe4df925cbd5b5b96e70a271c6968ed5c98569e2ef64c0a5626a87c6c3913d147575645341c2738666d737d7bc926d0dff8ef46ad325e786252b3f6ebb7ed0c5596c15a4ecf530f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196343141f9af00fccbf3fe8b321f58886ca37295263cc9b04ffa702d92675495b056c947a2bcb70b1b794ece88d51f0b7174c640c05771e60d560559825b2e88ca3d11c6a3c2c4362129e4e4190fd56daebbba945ac8d759cb06cde5e0d948f97cccdca3150f919b6ca04f89740a1ffa0589e4fa8085feae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a121f33c94b68e7995d6728b23dfc15b26dfa047a9cbadd9fa157c377246fa1063d938cd17ad7381d5565742c0e2b96dfcd71d3669f8dda039514012960e22aab24c86ca6f995eb46572080d6e690d5fd8fe49136c59ef2a09a2af6aa1fa7c763231bdcdd501062b5338cd1887892a26575e268651e42e99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h502b60cdb865de6ad01e1730117dc08212c11629de09ad4a5fcf2675ac95367bbbc0b4ff255cef32e30a62e76446237c855a05edd133762a47e0408ae73db4424035e6e86d27b5dc6b778f161377585d5dee2bbb9a9e524e0bb5ccc470e16ec7bce3fbfd3f4f66a6a46643624a3cdceb5a063b20d61f6bc9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12326046b62d7f88bd824abf799751a88520fbc447a78166bf0ed1777b1951c442abaae594ad3e58dfcb27e05217c5f3e326e3a75973cb95125cd0464b733be8c66ade09c063ecf2348b7e6f7678ec95acbc14e961e38527013e9e6ae09d783250b834fdec8bd989682815630421ee6c3c0189a2bab87bf81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h770e961cfb559ea8899c3ea2029f9e118c647981c42b1c26da96d795c9bd570c5d2b8f63d47f6c21e832a176b90b044745425467178f7b79aa13678c38f614c7d5382ef44c6406351ed09a70b286d9470c8e01f07c13927f3c8d8883d0d2cf62be613761e9dd7a8980f7f29b24246e1fc7ee146fa8bf9423;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10afcdf9fa38ee62068930307b57d5b76ecacd4454fbf40c30c6992b9344640747655b58f643e3599f365c9c3e554fb57e539a0c40399e218a4d579c6735231ad5fa59a7127a0968e216e30eb9b679f7c079c87cd64d5fbba605b0766586fdc1690bc88ed47617e59d9956e86ca098addd65350aec437393a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8520d603267feb9695bf5a86b119bce75bc7a298d42072916c388e9ff9d007eb6ca04dedd07afb59f57d31eced5d274bd5db9abd9fd874281be12ea47a6f856f6f717e678c4d1dd23cc741db3bf054c481ed7199da28d90c8a079628fc7e31bd98529f247e05148d2e531b8b24f5b2c5de7b46b487079fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1116a738f89c1c7a06d3200e11a117ed865deb868aff96fd3142ffd793fe59cb07f47feaddbee9f23cf40c13a63b710fe3dc1cb9dca993173afbad9ed353f7b6815e79bb37d0924f1a4facae3327831bedbe9f36cbdb827fe92aeb9ee622f57cadbef0cf3bba4fde69d91af1b1776e99c84e362cd9984690c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198e45400e7f80ffdef595622869b951baed651decd3a95da797536854d76f733b744bdddd29d44e1ed00f7be79a99b6ed12d7703a0a2f61d00faf5fe029834aeb7504f6ab68ef6a8e4f37a40c27d660bec33edce8ff085a8c3113154688f6d8cc39ffb2b9d7f2a45b448ca6f4f3a3b41ee1cc5a3bdf53f71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e95beb7efa8d1e2148f12227e68dc94460a9f0603d683e1a03df7328d16135f5e32d3379f2a13b907c29e416a04301713c57d94549ad830747338c50f65ac65352bb7a08238b5c419ea830a752104158459d8e57951b05a1f43bced4e8dc4b7db9f6ce1a2f55b32f956264ccdd07466048bd7c0d595bee7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11872efe4901c10b5ac5c83ede4c1bc10463e5694453ca97f596841248af1bfee7ffd0d406f60e716b866cd89e942ae011a8c89b8823d0ac4e16348e567fafa762b08de47edd270f57797d968f6b24f60687a83be5eb1e1d765eb0d01765c45997d7c5ee72ba0c44bf0bf853808bba399efa842ad34cd919d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14734ff540b72df9d2233b6a022b42fdb8568dafcb794a063e0d710f95088cb7b7ddcad3435a39028de7359edf8cb3916b9137d1b4d8c86fe9114e8cafc937d5295ce99079fe0f45e21e3d468af0df49b98b4298ac8c15aa28a9e88781b1ea3dafb351df8a8a3324b368c5c9db9514cb384faebad7a73ed79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d456c356f636bddc8055ecc0703bf4ac9e22d726f1cbf571cd3cbdf2470a845676ce64b740f636a120da60f01ddd3d700b5eb556cb95929614f9e3bf5f5bfbdce6dc282510638b26fbe77b6e7526d6a875e41cb2a7cc3168dfd78da194e1afe2b7a5ecb0001b37505b7cdc23d1d664a0240904e402ba3e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136f37ebd37c3f60c9008b787f1efcd18f0d669a4a9a11b93d2166d5b296ec0e80d73bdb233611c51c2ea5883822e6494567c42cad4639dfe43a3ced7ea81c39e612403b6dcc4bbecf2f5cbade3a44babafb2e5f99b7699b9adf5881d1d43bdaec9aa007bcf3a251773deb873da4472776ca9607a4227ad4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193e90065430b16e27f1b8f52c4826809ac5e0aa6f3165629f3fa2f9d0455a5d7bba48dfadeaf40b1b98cb1864fe5a10cb6aa1ab3ed9efc7a110036661a2a886690f40e507538047d447c073494071c21f14fbbf95a094b9ffa5d1c4aca0823ea5789ea530fdfbbe41fe7bb1c4546a8272b71224424f7cf9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149b977d2cd56fc15d82d0ae95612b87d5fbae24dff89c87c7f44ea50e5908e643bbf1afbc90f03c1bbd749e6e2c4134fbb3b30a63f42bb0d1e8be8cc0729ce90c6fae897510b4e8fd3e1e7cd3d39d417650cf1fc0fd9e225ddf71f07e88610d893ee278d50cc87bbe1e2c273d310552263954f9c786f40d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1031bade20423523e8df54df7d5503f5ec38dfe7eabc59e3b5a5bb6d46b6e40ddf9892f89ed5632d8cb0f6561a45ffaa8bc6b55cd24dbba98dc9d34f90df011d30f92b02831f1ac552e483120ced50841cfaaf6bf11a0fe65503ac3e545fcc762eaa0d3f837a9a12ca128b15988a48d3a014052c7a2fa5651;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147998c92f1be122417708479ccdbc78934cc5aae5e4bddc09a4b9e9fa66395cfc53629dd32a3f3d968e3ae6395535eda5eb5b65c2dad28ef441663f9635a3d78fcf9253fe61a08948d15c77db942b27f786397368a61506871be9d7262b019cc4325d57079556ff08b8ce6e188b8d915cabe8ddf8ed7d3b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h835be0ea66a13959268dbbeb16e061d36d1eb3489f26f8f38f9093279287285a28696259f8372460730b3e8d8b921faef6200e915f9d6d8dd0d2ae05748546341d8866a82c7643f2e9da005a0bd672aaab86203bc380ac08faf80c4e168142adf8161cb83c0e579ff529743b19f98a1db267bc232e59c2f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176393da227a9478451febb234b90a9a0a6832db1d769dfa967c1fa1cdbb3175994e4fac9f1801a428446afe6d942a15088ab8fa80c6b328634e9867de3bc2726d3b2294087d7a7d4cbdea9676d4b9f87a8bf2d825f0d574204c5cef503e4db2a1de266b6366a0b2a7170e292b975346f8094ce75a611074a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c17ba34a4cc71a78d431080b2c09ad664966efa4d9510f55128b28866d5a380e92075909cc3b018f8e7741195b36dbb44953e425f20a0f3adb9496a4766bf3329cfeb20b95123200f582bfe459d9abb1d5236a1d5bbe76922f62168c613e276b942c1cb38bfafa41f3446970f25f6657045e766a5cedf8c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd754669b7be687da91d0826cae1216d6783178209f3119a1f78230886bcba8d2051984a2dd596d0df28672864bf147d56a269fc37349c2938db71293f633214e4de2102940a5d9c55d18a74944d9f8082cc08daaa7cd68b793a0a412de2979e10bc3ff53af439bd6e7fba7b85d7dcf16434e358129fc8ff7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b5918506a023641ab17437acc875bd2f688df7cdb411aa7f7b57d0c12b34f9820934132ed70e1637fca20e5683b9850f16d97c9768e43067c8f2dc3d8bb5a5fb3fabb11fd0b673abd8cc7817d5c6d604bef7370e3c1b73bda9363b82592f2544219f67ac26c3670290f2d6f123f8a9d4f6f184a02526913;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88ee1d91e1a547b8d71dd1f8622341545d3ed231c455d1f37e7c9eb126ff46085d5f2dd09488c3c95fa87484d0ce0c8d40f1ba0fc83b6372f21c35685d2dade7d131082d14aa8c545400e486e984c3b4f5b6ef29760e9bf749e85fd8f96781c5d52510cf80fbef55b03a584706d4ba8ea42c2e5c71dbb80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa3b54c256f9ee8d501291bac1823177e6b9eca161ca04dc128adb3deaff09529dfecb411686beaa7d121b3f15bf5085585be19ccd61e32c467e2405d85451b4a90691690c48f8b4d34b858ef7d39898c8df965ce515fc478c8f9c8054895f8b644c27c8a0cae2cc826c117067096bc5c8058a297da92166;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13324370ca061d20d3002a4bbf899879dbe7bdd449943eb7475934a8ebae957fdff441c94e4d81b23b1cde3818d8ce340d5fd5bd7946b9e40a5fa079bae0db4378bb856a116c247439ad03b9f68979ce511cc189a954370b4177af56a357f52f889a7dd1ce0cfdef6e8dfecbc80d8d82c7e5b4fc688898a82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba0942a06e6177cbb3d06af6caf8936801c08a3eb388b45a05deb7b0a40567b7fa20c87600d90e14522f629e61e21cb81a7aa8a46343e24c8917e29fb77257b886bc8f06d48a6e339c9d8831b1d6c041e7e6a9ad533e17b167c632f4b480d41cff8aaa3dfa5237a073300f7ed504fbf0fc3b5ad79eee04e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30a3121a798d607326149a89b1582c6e981cc0d1f55768df5647fc58eb262ea2d73842e85b27e0bc7472aa63a9b756e440cda7a16ce211954f538fe3b46f579ec1fd1104b398f94b227ee99af33274f6afc1022ba70a3e30b6da45bde4c15858e6a45ae084cab13475aaa2262bd52643861729d077fce961;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7b074222d1c5c8cbb934c577d68692656b8dc2945d4688b8919b37c25e3b35cac853465caccd143ac65588aef70ec1254f79268188eab9371925d3dcfd606953d583da52fe4619771c44e37c87d2da9d57ba9839cf7782d6ffc7cdbe2415fbc34f4345cf391653d8513d2166202cf2fe22ad21554c533ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9fdfb78b4f098d8930fbc3f45e3e283cfc852e347e4dfe5ba30eeb5520923dfc74cb79440043e4457cf79e6940bc4f79d3f1f31e24cf218c467f3db8aa9d07969f1c1188eedea4c438936c675c190a8cd96e7b25fcb2d19a25dc50bcfa3f41f43db1e131294967ec65c3ff11f5065c1a742435d8d21b8d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1665f64da7a9b4191a9e8b46196bb655876e5116b52ceb0f27b40a6ab69025fafb243d769d53fba0d51e79d37b1678e82eff259eae18c8bd806ac3840100d210e3c053f6ebccbd96e83d2f0965dc2b844ea18dbd807bcc82bbcc224bb7705f03e6652b26fcd454b3cd7875a547d399d1a01bb8fac092c4510;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51a57b2ed45f10c23b239011f49b3dfc326d7125aa3781350eb3d0005dd849b54f49bb7d20c6edc2d5a754c06cc206cfa040e8b6e4392a4d7d6b1c62d7546f2fda73657ddf797c0bdad54e290d58fad2022e37351bb37f1ed0ac9adee41b40b82689a1a9fa06c13436110ef3fc4b11f2da8f21e91f1be99a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13630665974a0a5d8f172b2c900b3a0ddbc500fd393ae3220f9114722912861965a650f1cafade1b1082c815a1291d261f648b757bde021e10a9ac835d46bf225042449c9acf7f6d8f75b504da1ca970c2ee278d1be160081f52ab03d855d69dc31f3a8be645c23d065e7883690ef27b6570aa0c248396eeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcb3882bef1ac6874458085a896b45dc188835f3ac3d16d34172a0d4c73260717d6c40fc7f34c969b51058f95540e82412dfb3ddb0de07eae9bd977ee8c72ee058690df7f3542d3401a8fb411fe950a60ee4894336d98c6eb8c109246c8d829462262b26a8d86f347143d267a3098015967fc69123ddc13e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfc2a54f70c462fa7bbc184fbf8be21dd89c1cecbe232d020d18b4d287c0b88159b72dde5b10b56d60083204d6716ce08c3bea7daf1f31159c80621a33a77c3783180a42b2d36d28fc5ff0a85cacf20ac4a9836060e0bf141e2a857af8776a1f9646584376050f823a17bd89e73942d909bcf7dc820b4956;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3e10e0e2eec3a93c7961abeef29d648d2ec85d32bf384342db17c647afc4569bee2e6f02b331ea749b1ea260553d73a23dfd4f40bb48f9f2ba3c2e7d67718ccb56604e87f4a2ef5805bcfbf344c19c08e8d52c8d31f4227cea6e128f429366d03e10d84e15a35d9da86d9af73adf9b47116819e14f38a7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14905b47b8e1aa1e47b9af47fc051a16718f7467594a971a3d10af31320fa9ed8cf1a6c3d7611f9673d53713acac61c116f00b2852196cab3ac38c604fcea42bff1b3d639c42ebae5d050dd2b3dd6d21bfcfd623a570ceb8bcbf0c9fa9fbad1e622d46723e66ebd3fe821372f119571c23a36b60309f3b9d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19df457a9ec515de9b66ec373d4ade69a73405ae2126dda11d1a7d01042df66611b7d1edc36e168e36b0646e7bf2e83e61f9e644b9c953c89785bd1358f62fd6a191b3c80048677bf42f2501886d70cc3b7f8f2967a5ace2e6a7b2243e71d1f22317a9ed4d83ff4460d0ad708c95073416be934fe908c6a06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d53fc61c21adc2b5c470322ab1ae921ddf5c9551e26a3a5747b1285b3b1f69245da9b398d39e6e8ff0738240aa21bb361ca639dbeed583ca2c935560889b21e7a9cf64ab16bfbe95585a41956d3bb316a1989d26c57612f70701604b64b9db8daa61238cd114b6fe49867072aa8a2a284ccd8f4be68f560e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb33bcb583a109db9109cc2969ac803985e9ee4d3e400bea8d715bc1162c860dea81ea4b1de2f8acf47e30f7c412e36f174e6d751e7a775f1e780df1d8fa5c88b2445beb1e87b1a1fa8e5c7baafd64a334c48e4ca8d5f9fb35d7f9ebf0c8112a82bd1cca86746ffa04503ef111dee1de1cc7c6f1496fd00c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b99d9549dbc5166c6b32c6c9c88ecb874f9ab4185b2ccd0ec70d6ad46b6bf6d12d8ce26052c9b2f56a2a3a9582a2a560e3efc9878c00a9787a8e086548e9bee9900160d54a259ca32db8cb337492513c88587ae18199e73ab37055564fbf00785253a5e9ee42fade2ae9b6c07661692b1538391971a37b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed309440f5c49d371bf3ecb2c23b5540f84ae8ca3be41f294d4c672d97c57b9108fa3c344987094ddd8595e3256c1c402d8e6541ef35d53148fa81d8cf52ce573d544359f1f7718672b49607a28f244c0afe9bbae663ba3d9517e404c16a320866dcc6cf6fa0c8d96f4e42cb7836d94a80063b227b9eb40f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1542f9a7b781c0496e4b38b50226c01359cd9f7f44b0d66544f3ea0cce90df63b49592a0e95cbb26bd72eb76688d51ebc53f979ed3110ad39f798ef336e00ac531b1791427471692c4a62e425e06668d52cd9a71eab586fd8f6d9469b1da9f46ee4eb303649b2332530cb7d992a626b751ea172d63acd95e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be7b2677f5fd7b2fb4e57958da2556b1e1f88103d47f1f2f2f82add6fa3acb28a46cd10d70ec1698f7295945b8b73bfc44a1331318aeab4d43e1094911abfecc7e01b17562cc66b94530faa1833a555dc02b39803d730b1b87c9be4f22af5cffd7c925f629139c2282cb3abd29a5b3044f3d27a9e9ff8ec1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hffa969aad863136849c5ec19fc867b4a28aa28511198c5f5706fc0f7f609a1401a3192021eab443d8171fe5dc924305ee38692c5a6e4983013ed87fea015fbc3b8f319dd555570c5c3941b9071e013d13ccc17ac76ab30faf7fc8ce6485eadcbc8b86dc34c31f91bae31eadbabc41434ea8ac7dfa7ecd9a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17950fed09d6b04efe9c6dbaad3e1c1b27fc184092f322e498855f4345eee5c692507f948778e34eed2867e912abd3a299da1685f25de1d93d9b55e839790c5eacd5addd7f7d73ba3ddfbc0f76ae38ce152bca53f9bc3ec0c6fdc76746a7beddb35049bdb771aead0afb2605e663cd534b514151d0fc34b1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c69abcc5d5583744a8f1831a0c2371fc64a75b1d00fae495b8e944d88793bcd283aeeab23120febbff7293f8d57f10d9aaae7c9e7b67063a5f9534e5aec2d9eaf201f21cead9a52420fc295c7fa3e1273f8fea2cd5209d3c433b7a7ebef9b5e6c1c5bb97c5fed6f2ac8842784da9884b5cc4302cb75a085b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196cf22a9e60fd6488b6d56756dddeebe3a781393a821ae0305688b3b2a38b5af6098eddaff7ebeafb58f50b04533c8f1bfff782edc1c99b616ed1145d878ec7d5ce2851b0df8f38de8af6554cc0c10c51cbd55731f12143830d4e0aec474af0a8929435df671e85547da5ceb90840a416ff96820fa6f1d0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77fb23b895d1e75ddbee5d0c329d62297dfe9cc42ff79b145e1328dfd6757a8216c3fcbf5a68768461c5ec44f0f0d4a6d46265b1ed87ac64c201c4a8e0cd6a8c99e8ca384e8474d989eac41f907870b748f06c5e0b9bd72b7d50764ab04fe045688428ffd8abc978d3991608d2d03be0cae1a6e0d4c0dd87;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56a9d37ab5b142f861529c97fb59933c1f659a3d6f800b5b8cb3120e5ac5bb5adc85441443384e0db7a66110763b3ecca2d988a7ef9a7ed7b1ef61e1b06e0b287bdbf74ac06bc05f5b3fb6f089edb55af6a820a878ecef09af85c52b6ec6a36b3666a62f9b41944b78c20b4849f472613bc30c048ac55fa2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4deaf17ddf3d700e82e8879a1dcf1a86c7a6d87e2bc065558c1465ff8a16e79f0e6d69f16e9fdcc211790952a80314ac1b00639ffdf54548a56b5100fa9ff682826211ffe6c831d57525357425eaf980e66a620c3341361c376a66d7c9cdd34cee84029348e41b4aac3008d942989cac88cff05abef2eaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e680868773cddd3a5003afaf5d7220c7289e3b4b5f73d46ab450e523529d6209651c5546fe092291b01d49994dbbb0080047bf2ef352d07bf5ab14f23d02c5dcebb34f5dcba61ebd33e5638ac37c5913094d420b1a96c7d45cc72d1e51a4a3fde4797457cccb09d84236cb605caaa755a2d3fc7a5e8c6e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h488fc61c7d505bf87aece88f2f5c442360012fb9bb3e762960657bea3e9fa89f9ca2b84b5c439cdba1945030c037c62c269cf7e2c0a2a09f9bf70f34666f36387b46b5f0c1654bf539fd58865e0625fd06ec4a71e8b8c3da2b32b166a2cbde8ec47385654ff990f5493a25393d0266854f04ef28799ce643;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habf798e9fcb947032809f0b1b80bd9dfb4895c5066bc8c7079067669f03296d8ad704accaad08cf14631438ba12439d49a79cac04b65ba966b63ddfb3459e16f736a38ef70fbcddafae2c9208bd5afefd8cd571794287aaca6257c58f124ab67fdc35a50d07fa5b9c5bd97be3b1888a35c8d84bde5fa4732;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b2ff4617f498e2ccacbc10613a0fdb541029caa73bea949860ab0ed2fc33e6fcce54b5f0dbb006e9f385ddff2978114893a63c2d74c60af225188583870ebd0206a71837332b6789dd8520e0f92620b75ef62104aa7594a2bac42ad4c59bc606f81f51d5bea33da02bbfd601f230b330186f1f22dea33b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16df5bb951bb3918775ea41b2ce693d9d5e130859b79bf80ac402512b16757b64b1fcf86cc17b15deab472a9758b2d002fa207f74e1c34562bcaaa9d7fc36662a31b86bca992e7c474e0b3d22b9fcdb257e01d1b83002439a22c64ea89c0a325a16f98349469fc8a24ee793341a6ad1a922aefe62c5930e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc09a200cde289eda70fa8303c63c7ca3b5cb930c3558fea3e27491af1dd46c5e1932e266b887453da1ba6acc482b3b201cdc9467ee407f2663134c65c51dc209cb828ce52d0958750f26d7f0cf6332c371d64ce32ebc3f9693c9abf8b80c54759f1719df0396bf7c9fe2c1af80d9ae2e68b07c7664c884a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a4bba8bbeff0e99e2842a0e72eb738898f73b914c4db4ff078ef10c5592f806b0f375d68c5f2f42504ac7e6035caddd1c78a8463bf61a34410b3184f543576adfe95042154ab0fc75ed18263b3e87e78ab64fd26c144d5a8a8aa81ff16eca21d5474ec93e73462c56a3a951308c476b365d87dd99fa7cdc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5f427891f249d567cc6fb287c13ad143151a3e14989523c8e7e0e2f4d4e667323b5b2421023e6083c393e38ef40426f5fc3120e7526eeb3851f180598e7e4736f6da85351f17fc9f2cec1fb6808597531b9dd3532f3564797522385b77e7466c9f140b32cfd606d91023a6db1d2023597aff53a9c87a90b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4505606aa69df3800b822d02af3d9de9b109c50ca7ecd9f3a9186587218f3dabd1d2ffebb1c5100710fdf1cd5b3dcdfda8bab88e4d831777ac9d31c291a70b3182adbbad10867287731e7a34ce7e6f3094c566bc08b044c65f6670e5f9aaa0c9caae2d96eba84c5ac553c6911daae1852bdac4d4fb725b46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc47d17a2c3d4df287216e5262a336619927f6cc66342485e656d21c8e24a3b6990eec42d97199f085a049ebdeeac01517dbb171467a6f96dc75e9b659b8183b364a15e9d1bc671b17eb582ec01a8c4c91cf8055b68c4dfcfab5169b5766b1b766b8679f91a53834b61f79368de133cd54daa2d959eccc285;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haba0dfa93bf8ccb6945f2e92d9ab656bdf7276666a6bb0c0031f77d77f79a255ae6fec5debdd17af19cb05a1b537301e6ed55e55c170e40237a34c52d011510fcb375c7abeed29b1005bdade8674226e549d43922c24fe4933824eae960c71e101b5ac4b4149bec320753de80483b3db8f622e2a75fc9e47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e80b0b82db0db8a14f7a796c74af63d2fc6039f0b8012edf6d3c288f8284925c8f8e115d68fa7e13ccd6bd85d906b9578650f8c857a57a7d4d62b7b048170a67380de679ed4f64b2a86fab13706fab32b5c9e15e2fce51966e7b9bfdd85b978bf346e30840f0beed102f03bcb2b91212254f4001df500b30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f6475cd89aa7f972a5d6598925063495a744e1950d41ad02495b4e73c291c31ffe449f201b2bb718bb3c3ddd23915ea276edf1cb5bf15111d97a2490c06d7ae0a86f4137c50df6164080588e94feef0ef9d2045eb57fed45174b5786d882a0c8cc79be516d2b10933ebaf46e186995e6d7b33b296d1e26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10455ba74f394497f33c95a1d0348e5f5769d1177b8f718f48bfb6d8598b24c455e024d1a28698f7140156ff32120504c39c58cf26ae68d64693247f675e2f94dcd2b856b55eab9ff45fbb6b174ac828c5b50de100b129a9c811fd668c846b63103b3994d473de82fb8160decd54a0beef787d19c6e3e9afd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1940ef7c4bcefecf0a82b7f3a280753ecd8f1eef31dcd5ca1f00dabd4081fc89e02f74f8ceb043692ae1660ff9d7148c9c46e2511433de66d7ae9b4deaeadb8577b1cc6a1fb0ff464d56199e4ea22a4211fcdb1ebeb6408e9734128bc58c7dc80173918d38da4ab1182da4e4f4fc63ab8f9b44045b49c78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2dc13f5d2fe3fe8a1ce838fdcb145c21ef7af3413b7d3f121dd243ad24381ca4106d2188d82cba03c7af24588935bacdb5915399b06b38a0742d2eececad8d6e7a94cef3852c8fcbe74e88c06491ec83678c515e427ad10e9b0be8ceeaafcc354799df68a647a5752f8eb8bc4f955ed3cc44825812a66154;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e5b729161f7fd2f88ec009578b3ec4036bdc120ebba58dd6b4889b691e9196ae246e080bb15c59d039e36d4c6b8e11b37447d33c2b7e4b317d0f7fce34ee2d0531613bbd8f48024b447667c2ee735677ae8ba531dbe7b79f37822d85333515ba0cd43ba78b043adc353591c1c0622eb685890a0f4243584;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h206bd6d5986274eb4e1e082bed84ab3d4072a991acc751e421846b6cca3c6e41f9f6190321aab4020d728c30cb0ec36c7987e54ea1b2b2b870f88b4f4580523c6aeb7af075d03f79af2bd98b232a97c8176026c5ca50be1052437c45792c78a7b6bd566922d2928e47500bfeff1e2606c0bf4a8a3ecfa076;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106485c6b9a31c819779b446a1e9c9214d5a03e72e8c237b601c6976f5d183d9779d3cf4d0b79093087a32d805b89c0c364c3fd56410dba4ae4d946c5f7c490c7ba9f41c6ae2c4b29f279464fbdf8e7c53edaece438cdf8102a4e9d4af0d423a9813cd9b6eca6ec2b36f79d120f436f4f2a6afa03b02f945e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacf8d4e05776f6a5164cdf2a8ba56e14d2a1154de6eb58a27f4f907c5a54ca1171646b5b899199761c18dc07eb6963ef246dc16468b0e4b283eeb839c0f9a5a3a9197c96d61d336fde21ec19d027a9113e46c8236f34b08e40190093f6cd539ca91b4bf20cdf6d4cf24bac157cf592c96a61434af8d3dd99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a111c96595530d07ad71df1529bdc387695a9eab990dba1d3c8f1ad614586a75e64bc2820abc2988f432faa45ab48e3db9cea5250f43b30ea37459f47361b27ef456986956b5124bda395d83802d19aa56abd823c59be1dd3221b8bae47ef8c43e4a616813c02bba6d0287a1914d5fa66db4766ed6351eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9a3505d9e2a4266ac95979d6d02b195145636295386d9bfe0cad1c56a87774d4aef4c1a3e603385d122c1f60f67ba0b8977c9c06a21962dac4f67e29813cc5732902bb6502d8fc9af7e249ade60f1d52ff73e38430d3720bb43df5340935bb113eee1070a7e592d4ae5c3f3cf00e672c34e7d43242c654;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h578ca49c1edfb1c669addebd24da4c5c36f6c31fc0d7c9707e0a0fb7f2a0f663128deef0b840eb20296fadb65b696897c3d62686099ea03070d2ea210cd1eab2fd698097cac5c0862d69a69aff6f35b00b09bf8df91355c8ba707eba39a95f371f65dad80216f749a938452a136a36895821767fb430560c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105ec2da4c27bd58d4ab03104d20847d26018f5e3bd73acc1d1c7047dbacdcbdc4ec9c21ccca0aee777ea7ac4f70481b6fc1ca42526a48707444eb0de2627c2727aabd9429e37468c2932933970601c4476d47628f05c5ef06fee8849288d8511c5e412497b17bf66243e6dd14027dc0700308fff2aef71b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e660ca23cf96b77808f9a2814a1a1157a026c079c2b83f113dbd1e2ec4199c9cb65b0435ecdcbc0d9b31ed96ebaafd0dc12ff87266e301e6042b6ebd70db5afc47572e8c57fddebd9d24b8890de9bfc25ff4c62bbc6b793390688aba6abab4cfff063c0ade9743a4258bb34c182878d03b0310eaf747132;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha52c05c43e68241d6577babb9899d832e107cd1faf4d363e494dfa91a77e119f3ce6995a4797e339045637316246dda4cb3325c849956c392135c49069cde98d2089f50f673003d122e9943a518a1cfbbe425dc754c54100a57c2a2438d8f578e876cd22272775ef7073f1ab64596774d59f6f0f96e27f85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147bd4f0b7f9cc2f7b7bf599da0ba44d2ff9882c10429ed30ea726b838fa22ca59a0b86cdf8da9804e387db418e41c9262db87232edf695ded616a7741d0929261c5e2a963920c98e78ed0159effd38e825684beff41989373a8857477e7bfa2283337f0c6e0b63e15b5b564f8bb7866110aad71b455aa91a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19948037cee2acdeaf4fad054167af08a3677fd18ba899782f05e09cc5dc410bac5264b0012a0bc2104a2e62177c3fa5c42fcde36962a73c3bf71baa9ffef4c8ca752bee7bdda932411532d61fb36b0434b3b592fe6af52767470170c26fb8c10268853f6485e9aae2aa38110124ec1b32b7d34db61f7c597;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e0a808ad19ebade6d9248d693b66fb8b3bc57aae9356cb72e80b8ade8bbb9bf4a73eef3faa23e05077a85cc8e1bed2ca03c23352dc3da7d35aa5116f42895168c253871c2c463c26eaf7a9a8210550c1340c93d38d84acd7f2212708231f5f7e6bec3f97b1a6df695710c56fc41cfc6f95947cb191f9f64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173a912aedc3010929613bacdf694768a4064c28ea585dbd19417ed4ba353bb476370e232f3f5005b945a75320730c575774b0ac43d84958b8b623407086f9dcb6e2be187ef6daabc4645f86b6721bed3a187183a52a0ed0ff626b13e125710fe207442a4e153c46dbfd3c4325a82591f60af4455e7375ba7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5738af67774b42642b1e57cc618938d5e2a8baaaa2ac6c92e0681502dba770a2f947205f2867703a1f691b64506e258fcfd230420b8fb866419a70248da852acabfc278e24398e85f31f4af8cfe12a2886cd7c529e106a64150a3e6608dee502f9a4b04fab6f138d6be71dca0f74552263cfa91b75c4c5f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13453a09d0aaf16a63a58fddbf33649ada497672ffde688f201bade5082666c09bfc41ad1f2d5c0099e796934b6acebf9684cb462cf01a2ca593a33bd984c0dfeb586162ea4a75c81a630cb3caa8f0ea958330cebdd808ffb704428b5ad7495f44cbd154ffd73d15cde34e5f4c96de100c3eaafdec5f8a329;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1370800f0b5b97f5adf4d170ad1421cfbda0d46cedd0dbea92581c7b833e9818302c75fe4b983246ad9796755a87b9cd349daf22a0d170eb233e04b8aab16241b4d90b081df3ab47de61464d584de98a03222aeda7811e541342c4e5aa03e323c56c39658dd217490ef27317cae9a813bbf2d6f05afea317f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79789c55381a54e8cf318afc6352129fb097a4382b6d261b1b7d3499b508354cabdc5ddfc81f797538fc3696bfca8830fca7298a2ffc1174c257075b9510ff5c9ddb66e13d470fe72a57a0d91c2354ce749d29b315d1591efda80ba961fb063cfb02cc7d9b17ce894dbc10c3f108ece07c3696f7e6687d97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1306380313e91c0504053727057bd1a145642e399e35d1cf627cddc1d38bcf54a570d785c95a3b8fce1b1964882a95e7111ec3af4c12090a26c90f61add4c10e8cc77e5e2188c9e0a4dccf2f36cde0fd1c4969e96a280a24c492288fe35330c08540d06c032b0ccd36d569ff81c7c9fd9d7a9c4c772e3c794;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e62007db18490b199335121e27e01d05ced4bf61651228dcb9129809d44ba9b5e861c77144e7ba94d9985cf2e512694b4fc0c580766043d2e9dd1ef391c2a4880cf9b73df0657cfff74f44cc151eea27c2c3c38ba7eb54f29b3ed183ddbd4b0c9cc8f58bfaf682811ccb71f70ae68ab4824bf4e6ea28b388;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2ebe1cb13c20bcab10304548f068e2b85f0668c4e947bfb7867dab1bb5633e38fef6c099ca788aa693be420e94a59f269631c8936397650885bdec66e28d384132808b456553d0600930989fd8f8084793ff92a2c8d9299b504f3ece802d42e1c4b6822163899384ac25999a901268839f742c8d2e036a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c5bf961db551a80f58d85944810efe07c75f8833636c2ba4b134af0d59be92af53c3b303ae180d68d8f3093ccdd963871901f3ffa89aa373ccc5800921014f533d56efc4f6d1621eb0faecb0c1ced587f3296a2e35cced7d3b2ff4ea14060e6ec57639ca25d3e2f227317de08a1021a3ce4b511704fa0d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc50e23fd48328d4da176f043fe3b5fc64de434d236fe326a404c5634b6ae614e18e7ebca4d6ff155cf015ad6213e1f989a0fcb76046b36abfdadc3c5bbce50086011148d477a06b21d379a865aacfc1a89f196ba997c7ecf08259189f1fc2467bc89c4492812ec7066f9078a1741bb6fdf39b661231baa4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1507b07497d24ed4b8c5e985eb21be5639502db678c7ae287974ac88dc9000de8606474aac2b0b1222ea2b338eabc593bfb5670b764abefa010134b182b80bd4c8b902c8f0a5bdf0bfb42a86b1333d63dfa6c75070764424c9a447f5cc77f5d2da2751892feee21ab9c4b4c748edd0f837d3bd20dd4c3cc2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103f903c5a682172f7566b2b1fec2a3f90205aa43e2f2ce737fda6f456e1944cf769432ec8336a1d2e138208887d8ea4e23821bd61ba81a7d2ffd31a09262b470dc01639b9877a79ad68481876c053cb4d89d7d5ae6ffb83e16f00233327ab624c9dc611777dc9437c1a1592dcccc9089142273ac3c7d2753;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fea0a4d19347a6de53ac96aa3f836ad6518aac764f6c0bba2d9b1ea094a664d06ed23ae4c2ddcc1c904980110a8d9e9d18441bf9aff97ddca9b532f6ca6ecb77545adbf53c30d2333f30ac0fca187f4345c908a4715dbb3c78e4b5782e305aecee952f53f68b56215b06063d0511277a2c476dc328a74e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199e053fcd691193488fe01f63d1179807e58f67c8c7f48212d0c0dad68d33a7a67f127777c41e5365270f7ce65471ccd7a57b684500adc948b4fe0eeb4af741efa6aa1206798e41952e1a8fc57b6ebee9e10edda22666f82d621431a93aca2ae3e890fba2034c0dafd0170455bab328c03f54b6238aa244f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha049f65a03d928c7d0e6bf3b8f61ab41c098c71eed2e1c0a910ae2474d557e4cc771b7c3b51e7e058838368fd0ed41ad32115e11c19c1df0ce112ed0c6e83049917f623e8b6b1902cbcd0b2f78b8af79230d311fc4c9b4cbc90f0ffb131e917257e7df4a0faa716122febd9741248bdc8d57ddfdbcac1ea6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4075f62036b32a0203b5afcf22975ec6145872b906cb71bd90fd67bdb3714ea910fb21e3ab78a7921e9fe1be60ef11521e64a4c92c98a24c3b3d6b343ce6edc5d22a6b2c3c2db9988749996e03984e6818914eb129d7843b66364938971508373b2d401d58d835e35630c7cf6d0442eab2e94813307506da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a50a16cdfa50fe1f6abf088b1e04614e40b6f5d64f2eff83a0494319b497c1370ff46dd0fadef85f4cc3955c7975fa83c84760989416cc37e5d2527dc331457bd13a1e023b991dffb22097c6a31745eb201dc1b329c6602d2f4e4ea996b11fa7a7347e01afe235811a8f1c5764fe5df03268ad4f3963ab71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d6792f22517a7ba02b41f83b18665d038cb6086085c4083346b5e9109a3dec21da0cfa626f1c34001dcb006f14a8b8642284340a71c6e6e70579b1a464f108f72d31f9533f7889fa2f087eaee71b5fb76856879bd02bb879ae9c34a60d48c4504d1101ff5fc4979e1468b988d52dcf1765fa2b0b5d7f5c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7071c25be97597ce6aad12b80a96bec89f629de8e1157973139dc42c92a1451ada9244aa03d6a3084f11d4c31f112ef38b707d893ab84ade5336e9f07a460f7c355a13bae49096711ec83f918144609a8fe4ef24f688e10da493f273a33207007e46e94072011354b6a91261cdf02bef1fbd969da693d63a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1061635ef297afc088c6d7cf01317e157fe8f45483fae52147085a40f13a84533faf129ebceb0a1b1652a77ff4ad5eef020aa696a357a555edaa8c818f971cd23710523901f3d34a7081d4f49dab530f4648ea8566c90025f924fd6d341436c42f21dce3e37a6149f7bd6edbd1f34b7266581bef85a054230;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5907dc9dffeba6ffda3a0ac54d41fa3812ea43304dcbd471d4041f222b0bf3c0447560b990dc1636ef12a85e87d1b6a07bfb98416342b39225a419d3ca7afd0947268b7855556adb68370d26fa0e0e17b9c52c1e8ed9c00b8861e9889493b49339f6e4b83ff18031b2d341f9207329d488c981b09c6fd65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e68488dd98d09fa68e8817d56d00bbce04d15c2be8918167bbf092a1167b91f39458309c4a4bb32cdcc70a782681cca9d5fc2ca6d21303963d1cb27848167efd216223984e467a5e2138e0769091dc23afdeda0b6072c144770eb2ea4d7284888b8916ab1e6f615163b94ff551a13bdabf7376f0dab59a41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90cc9ed3f23531da16212b5713bf9b6231df1c878abb6c9c65a329c826da00e8b1ca4b60af83f50f78b557b0d42be7b26436702906b9c9416d244c5561407d46b4656c7fcecc02bbec0ae703a80df27042bb07e69c19e6afe395a6d288884c7e0a49ecd2cd4af731ba9401bb66703b52fb030f37ae9528a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf24066e159535d231578b0a11f3d9a29e5ecd652425acaebc06a6883aa731950551d21f377cd7324be48b5cf87d1234849a31771dc9c9497e41316880ea74b918e6d09cf0d12f29dadf8a370df3ecb83937a7e0860c9c9e2eb28cfcf22119d6ee396bce345da4a858e5d538805b90dfb8984ca87ed5d207;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e0ac45f1cb6872c5fab9d9eddb348c7f4b85f4c12d297c83f99d849c0d41227477275ab2c7122185e4b971478126800130fa4ee5fe10caf11733898aff7575926a3457475bf01d5f433b2139b5fba4c630087b0b14d338da2235951bbbfe0523f96009fae2436bcf28cfaebc9f3afa79d26dea9b08dbd74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfdcb3880fb802467427147aa5bf2e991a2a5f1f7fd07ba35be1f6e03910c7dbabd628ea5ed4abb7d95d7703cf9d396cc6ee7ea79a4e556e306859ed127800b7fc5b92fce5638e10513e7eaa0a4d441b6f696a9d42158197f40534e093b1b3cd32737ce2f2c99e44969153fd9b1f683fce6305dd42d790088;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ea11c8d5be1631eee9acb453da706c77091c74236077a705bfa403ee3b00be19b70d360ee8c33318e0aedb6a3f30768ed63e911867e0990cf13020d386eee6f3d332695139052693203ebd05e333196babbf4968f69aa6d16ccc66591f044f093f533d8858216d68c46d14a2784e0e00606472489e83ca8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b57fb7d54cf593e5c1df9444748e3e57a92dcd3c1ebf449b050b671201dbdd95c5837caf6e33d473b8d52941dde49caa6a839c08838f60a4244ae1b613db8009c42ee235d22d36b20b0ee4e38727919f3ffcace72cff81051896756ee6e6604ae3d7842c4f4b9309cef00abd9fc1e506861c3f94b7b44f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h992d09012b604e809cec65352ecce4b0a4b99a340bca3e334ffb259f3eb8b32bdd842dfb9821efd10d0355affca20fc3864d843c53675c9f3a4458354de650f3f2af677879ebcf1aad2205116e57ca77d4a8a17a39265a3b6b467ce58e5b1998cfa2aaad7316ae4431db25de2e845f50141f286acadceb61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8efa8afcb3ec527728bc357d45e0c9d2d4b80df78efefb4c66c2e99e7ee61e3e54dc0b3c0c1baabffdfbdb7e9d55bd3c79d9595fbf71ac6f868a146deb2bece42e0b1c35bf69b5f5018ef418a246ae28a4ce80a8c33fe1b818732a0ba079115fc885975e4635c750d89c6d3238e8c33603f25a53f7e53df7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h290fa3b617e5157830e85e6854f0cae9d597616ef955a45e29f478ded54605aea393237c785f8de720d2c45fbbbf5b409b5699ddd2a507231eb3939ddafc99c211153e11cafee04a866307a48d9c615676942e9cfd824e54b5df0ad7d5a0bac3d6d776a702169c342f19db373eb6d213bef6523f77d7a242;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81466581085805cdbf5e3b3807051f1e31220d9bdf3c33aada4cc08b4ba6e289d3c807f9f93490a16bdb15e79de1dfbbb0cc6c77bf5aa6d520c59b6430c5bd906d82da03d7962912a6d7f75bf2635fe99d39820198e452ea0d2db6e814b44504cad7e2416c303adb0ced727af8c96370018aca1aaacb0b79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dedf5e9f6e263a26769f9f12fb907dfb0d0b446a61646271918634ac07adaf6f5b628da521a1393f3b97bdc78591ba9622a81b9980014754f20a213990805335da8e882899624c3ceefc8f8e370451111d08e354d12b3bf2aecb96e8f37e4e1387fe428ec9f2aee21759932ec76a8a2dbe3e329b35cc1cd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b1723e2e92a98570054a8ea978053bfaaf74c09f6a96289426990838a7aafddad805467a35b6a96bae58bc7b18476f173dbe07058a1ca494af0f4d3ca9be8a4a4899350b641603119a3ef1049b57cc9185803fd9d2e8a234941146b4a17648487cf33f0eb452c80575f7ee22b3c55255496f11d6eaa0a2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148911d0f6569a76ce2200cd08c1506269ab53e20b083cee96694ddddfae858d069596a849b9e969214b836589c326a6e122fa20e1d9ab2ecfd88dec957e246f99dbe675acf2ad12c4c6bcaf5581cbe9ac82060601a89bafb0635a1172557231c144ee4f20ac4814fa7e62514afb65163d02f29d8237ad6ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b89be885c94a2ddbcbd5b46d00dabb9a60c58bbea7ed8aca4fde42724af178c9f55bd020da5c9d5803b0189906d94bb6b4aa3c9b5a68d207f3ee0ebb6ca73e206359a891269a91f1b3e1dba45afd9ac2f3cbbbe55c34198d7020e549451a9339dcc89561ce74062afd8f945be7e8a8b2e43522a70b82063;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bf5bdafe3dc5079e17d30e315470615254a4a16235784679b6802f7747c8e62e25983b8a15a7317f731b44850ae65e0fde06dea1de4f5e4d075a36624f23a5f7843c94701693a7decda3bc43e71532eec5e4033dada8690af3a67579914766eced3124759036a5aa21c04d090e3bec2269ddb801fd414a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h902273cfd11d3de787bc5cb9292c341011909584702522cb9e537406b3b7f3843e6a3205e93da1e3af76d7d35287991b0a912b5c5e9a86c0cf39eed1f88169b871e2f66b862aa302fba098ed51aa6b60ea854e78c875609d33f5ba2b37412622e15582b547eb9752a4d7e4285f5e0b4193e4d8d83b88fd0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h215abf4b303f9654cd9014732ae262c6d0865bbcf8e0c17cc13b75a22220d0e2d6d04b99849f9d9fcadf28950f94121c4267c5c9503095a3629c74b1c814768fc7d597984fc2d3e4eeb332f9c8c51acbf69980f9b184cf6cd1e429363b91b2422dd1d55aeac2bbd971e215cc7099a56df39a8e10db39f0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b2e6e3fbfcb4668b789357636d634c1731c43e7fbbdff1a46b30ca08b0a8ff4575e44c05d4118e5fbd9494d3e5d24f58e556c35de1b9bb16a829c2d82ff7a507198e31364e204c219717858016918ef5733bdf4211e079ede6560450d8d1c82ebc1627afd6220c738a51325a26699195a78a0b863ce5334;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc19e9a2d41be7309bde3783a98f5fdd59e81b93dbfe80abe05967fd263600b98c8e7631a3a34866c3306819bb074f50532b5dab015376c5e320235ba7c0e40f0b8a17ee3097b026d7b0bc570cdf0b0b9a581d5fa96c0e9a4a6193f973ae27b8c9a4ec1f382f1ee9177d8833a2f636d935843c7bb3e09dae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8db002403d48d2e69142981a72711203e5876ba28d2e9acd040ee88f746770ec72098acdfae3e4e21e91dd9d83c43dc209c000c00d2719b8c237360c404d1d5cb9c635a49dc3cd58d6b38d6939719192e69def2dbcf3513777768d532fafd17aa390fc424decc1f7439c3a7fac50c427ab08d868f54e29a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacdfcd2309f6a61d5fb3539e269ee73e4a69fecc3e5121d2233f2b938237b3683da24810f47a73cf5b0b6f9586e7977df72828bf72ac5c9e6fa6e0b5426b8dc532b40d4a6db65c226394871bab05cc10e790c3b8d33162bd9be24056bc92a8fe77f08b23befb24c61d0cd866cba0fb9fcdf762dfdea43fa9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d3d20ac257ba3b0e8b2230552270323e9f62608d15fc57ec2065c607c54c31ba06afd997adcc374deb9a33650268e52c0b7aa42af383b43ad5ca85bce34ddaa5364ab440795a08524365349aa5ca901c8a012473edbef7854adb906a9c5c680e2cd25ac5f5e0e0d1858b32d945e46953c82fb58917b0740;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he322bbbbb3d1d33f5f3d99fff55baf8ba378d065ce43a02cee204aed671fffb2cb5cb224d666372f6f22f6710b7d6ce9844198b9de1b1825e1be08893adf63a07d8c0cddb925bf51a02ec2ec02141e0eedb6ac796b84f2f734affc8c4a59e5dd491da69fa2a5e95765bfed0a4583b691521293ccf2effb00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a36758e12c8978695b92742d0d51cc443192eb9c1d2d0f299c6e5e5d9d5448495a4de0a79711af3d0c810bb667ccf8daca7fa376e2427a8a4fb66da46c2f6b339b01470697377bb78760c4e346934a3a58fd1a5ddfa340f4b52f0cacc59163c8046c0203816f64c00e6a6b30d4ba57c4bb6ed2bc0f31f7d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af1516958306c54b58834306406c72faf7f42924e85c9c82e26a1538b0dcd4f8d0efc1655d84088464277c66766f46ef6444fcdeacb8c38852c8567bda588a916f7c2653d41d3ed15b45c2dbeffe28c9d8300675233453450b22b7e4d82bfe2c9bbbb20eb5b56498395f445026a939b9f828cf59efd83aad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd79bc2b9e61587a2adf3f3994fdf8fb4d2d07b3bfe69ad194e13e731bd5d812bcabdf335f227ca2490c231faf28404b375ebb7fa44d416208d7ab275028aadbf2c823c5a528e4e44f906edc0dd4ce8038624be326f8df93ef9374d014e017cdf1592c4df52e5204ba0bd57b589f55b8542e59a7420005a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d5d706f57e19195de0b260c3dd3df951cc258941fda9a0e13dabbb5c099e91adb459262faf38b4123200aace4f5c31f729f9ade2c2305a8a3c7ec48e5cac4c55075289341b4d031c7c2d645cf77870804552156b2e9ff60a28393603b2b4943d6e9a535c79ee7ef6362070007c7b3549abc8082bcd61666;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1560ec3c19b2bac1a59ddd290d14b3cec73dde6b9c7e2c05a2b8af97b2e81d2dafb4fbe1e45d3173a899a74f2d635bef58d3fe6c2cfaf91f9dbf287ef268bc4a09d44de0ea50435c3dae543462c5504f34a05aa8f2656f01d59127e37aa068a1e53f1c126e51d43243a0a00863d2136053c68c9fe23555d73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d7787ad0f04b6e895baba170c2403af2fc3c4e70fa0956709f2cddee4de60c7242802acbe68d5e4529ffbadff6163bba39004c3a9e1ee58b42f5f9bad32005f01fa2a39696ff20aacf3a31bc6e28429f132a7ba684f326955a41fd197a0e9f68e7cf91d036a73b82404a0efc23bdcab64073b5008014f91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd981ed26a0c46a9019ffc2b987efb488d6d2967c17aa461eeaa29959ffa77fc9f6a4a86e7928b58254ae119d06f09599e8593a34733fd838b826f994d23d1c3a4ecfaef8466e0c89aab04aa9f39e109dfc2fc941ccfc59253b8a834239825585f49d6647af1a4a94759dd4d97f3342ba07900d71910325;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fb130a66ffe2ecab79b002d6e1b84c241dc25b621b3d8b494677ee077183c0b7da796d95dcb0677dae8190018994c4b0024740234ac5458a3e8c620d02f8610efeb491df599335d792f858ed9009b99c48a09ef558fcd12505d721e0359ad277b8d21cbbaf80f25913f24a2fffb1ce30ccd78142419670d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1811ecff0a43ea06efb62c9eee4d577c994231ac2e106741d6574e2638a5032a57598f07f7b329c822ef2d83557e1737886f65b4a4dd87c72d63233bde17054e18da5a0ba637046a1e04ba74760a5513b841ff635fbd5e0752944f4b81a9e30db823cdca55172f0a02087edaba7b95a03fb47ff2dc65b2514;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32c5d8aa2b0e381ab373d412a22b9f5e557e4ff62c61e9b4e8c33ac27c6ac2c413c6c61e2c81299e6ca7e756d6ed4f33b8f86463de42cfa597a20d26e3585adef67e58b5b4b00aedd244b8f99e371bec46bf126f5ebc4869dd16685f65ffdb200e775838b49a61f99f6e4aa1981cc0b92b44158f57c134c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2ab9d0b7248e68be663e7fa1396eb25e407b11faceb93b217b685c82306f85b49d4a4c1ec59e478dd5316e0fbd9cc76c92c2da422c09debecfb77931a6a92adbe2a654906b1e4f464dcee4d00e40ba4ebe503a214c64c8355b544f1c903d3e7a6bfa5fd197402a99085955dc7d5d2868358a03a6a734cc2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136d944f95f22a8002df3a1f818f306b208b5e00fce776732267910f1f32d1df1ac194943eff42cdf25fe4a9a54bcc0b2b0f148a2b593b849baf9731289ff6362729a52601f5b5694a9044a215a1941c05f4c2e7763afb110d3b0c259c9e322b613f3841246495cb535493326e39c50189c817021cfccc3e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b6c52da903b983b7ebd2ca0673c1be8b78f595cfbf47113a4bca689f24fc3253f858860958d298c087d25e94b8cc307c3cf7a06cde8112caceeb1e57faee54aa721040d538df9bfe9030532e925e7f80ca9bdacc71c9248852267b912d3e0e33b314d34e01f9f7c4091caff4101e62894eaecc7521d3212;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h858eb28b32f757222e2b57da73a4dd2436ac960189a6bcc6d8260fc3110dd3e34e01c5d43697e958af239df5b0be740f6c1367974b106508982721c0e11d514d0762b3cdd9233e6cb0a026b4afa9085d08231880838ffc5fc604aace43fb077a6d20ac7e4c36c552f00621d5833801fbb26502c770cd4621;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d923917347ebafe0a75b3a045ba55274a503093b14646c5fd0bdca980b3a814fb412a18edf1811f40099c2943390ebdd498f5f25526664af0caf22260312cd6e4035e10466b1e60fb788e0f63be8e4baab669211153549411c241a40ce3a2a9f825b06b82e38d02c89f13ad22ede9b4d22e5f173d454e15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7b4a9a9dc6e3a4fa0520fb9fd3d0ab6fce4dc4d51ac54dac79eec8563d3fa40602af9e8f68170c43142cde42d65cb55275a21795731158b6d0398f8c718c8423c0acbbda45863869f04e99d255c84f5cb6e02e68082c1faa4ebeecb15392397f47d3acef04ea56a540e49185c99d50eaeea452881084f52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9892f8e181be1e459c5a07b82d6738823181acb1eab665b1c26f641d3ba96efb333b39360ab1941eb590fc5449b537935b88d747e4da8e165c7ba7bc571b4d619cadddb99ef67ef6ea82d42de8800fcaa1fc81596564305a0489e6706d15fb8cfd4cc919426e40fe9d10179feea2f16976278db2e776d0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5380e2d77aaf4322e03e14327ecf3b0a3ff643c65de1d1b0b2b273473040666d6aaf7b3926a0261b8214208106741786d0faeb45bb659c91eba3186dc517e820118369989a849dbbf3d42e034d59a75dfff703b86f4a01c4861c93a0104a3ec1a7b1a00b37b0a76bf111fe87fb708f67bd8be3f9411f5a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be922b11a89f4d2d5e370449a5acf27c34d6f8a67a446531421424123f546d561ef2c00d1be05e66d62148b5a6ed9c8f11039379d9d514331a51a1ab5e41f6d8c068d70c6849a7fa9322ba95660643777e4d744c9f49a98ddc07b1f360e6447e2823976236996c7d6f94f2dd2f70731ad224a39bf866ef2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h223ed7bc1512824df137343755d7d2430391478b8a0af07d57232a72cafa2e999043e8b1fc17dae6ac8f7ea7150f567c3c1c32f89868a5374ec823d22965dc465b034e766cd4eac2ebff43f40b0725a0b947216db3b0110dace340d24e0332f07221d8657f7904e180992482fe1794d5d3108fa3a702aa8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1401d9c7f65b62366ab05ba905dfe597093f5030aa6507d3130364e7685bfdde22f76610f392ba9be1ce9fe420cf8ed6bc43458139e761cb1a529cbd44a241c0c600020cc8780e4d730d4ec6256d37625e4c83beb5aa28a3e03e90e686e240da03dc6f9240b28ffe86309783dd481838edffca7356e6beabc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78247bff8ca5313a1638bb1fbbae00137655c131ab3cbfa3ba9c9d5a6ec45f851d17b8481cd8dc111cba8f729dd0df7fd53bfbd067dc1d4fb0167f86298f391b841958555fed8fef12a5e7cf5bd9180b90c0f1093f2c713f6a0e1cd1448d5ed20a9c329eed96bbc9aa7f492c579b38be4a906165d1b1f121;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3322bf5a3a3d29619b3f647d4e8e38ba2219319e649d1842437fd9cfcb1215b25f95077dd33b7eed174be23b126129084fe7cf8ffe9a631d36341b9c931c4c095228f77e1aa65c8b4d7c13657c720b25004cd5e8afed958a76d2fedf1624984c4b2f80a2e4853c12062d8bc5d33e6ee29a10f3ae0de69e8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff0f8265e6fa2ae4e9d5bfd326d51a3d78db58a13b4aba38071a1436cc780860f1c39d8149633544501544ac2a36d25780018cd7945316a9009433ba95d32e6beb08141232ddba990f7b845c2a729dc03e447e1366fdd19ab4d495dda9ac05f1e33b067478408ddabc74aee597ad7b96bf8da86a4e73e37e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba3d7997b91df673f919162e63e00d5d9ee1f8bee71b9644afb563db210745fb0f29cd9b75effa577692f0cbb3327fad530027f55e212b4d15eb2ae9eaac88624159e9fcb2a8661bcdeb512a7bc09377b4418fd93d4ee25108a4dbc0d0dd1d961167e896cf0c00f64bfe12cca581abe6b5403e2bf9240aa3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fe0ee953934b8b760732468475d81b6f4f351d7970f20133af62b79481d949e4db4df3d50c9d998776e5d32f95c76842398b34728b3e1ccab3fa9461344d88c0c238c54b3b96d950aacede557dc37caf0f20d68278ba080a8ae9c167c5ae74ee685bcd5397117d199e976a13e88143c0373c913267f9358;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4ac75c9b7161e5fbf9e03a9283c263978d1c963d0a9c5e44c00e156a7c24c001bbfc3beffd8da3f7d703b34d6a843d0c45bfc131f72cb048f926ee33966e7fd4190816799f4982f92c1849fc333ea9e7f93d86ff14eccbd800de3c0eb5495b2b4cade812a6f3c8aff4a3aeee243302e82f2b6b353974cf7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e9dd6abb30c4a377ed0517b5d3464d7a71e95985e68b92105f19b1d28008309044ba96ade14e7b41666320e777a60561221360f464dc1f19f74d5a8aa0652fc4da03303d84455e9cff19cd82b94be247781b00fb0339fe6e19e2bea48b61d483b24e8883647260e533343e2c13d98106de31056db9e045e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd04e77a7659bfc8ac44ff59ffd54d843f2bdbf0350e1d85b1d380dcf0e7f41e6634a02e8dad7f5fc4a253401c682ffa9087f6597ead794e9a596cdeb908c64e64367ae943f1a92f06bc611a1416b21c6c6c73ce83396f1a81f661bf58a2a14332f044e098e056e1d229c960be6732d8d8a130daeb79a7d7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ca5194e2e10b9a660c9ae8c0ac3f4c8dc444e8eb1441edfd3f0eb91e7c4e0a0a21f0b856271747604f5bb04146bc7aa12dee32e7d752455ab70d49c3029fb8ca61259338e8ef420aafdcf93c73a01bb247b3c708a0036e5baa2628f5b7a4a951f13285222a29c0583232a7c96e2e99efea01630212ff2f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ce7a458f2c92c5b85f09391af22ce00500819d7c6e19e4487e9db0e2c6ce25f25f44ad196dd7b5a709ba0ef35540918007871cff0f7ba3010d63e4999e8c68006c2c0cca44c58f35c2d211523974db851b93028c369892d69db95f36fc21fee5de82ca9fba9801d3bcfb9921fe93000e85c53d33570cd17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d74c25184edcf72c012d78790d683bb8417518f791e239d0b3d9405c1f51ef21a1af2bb5176028aa507d635cd4088964596eda8ef9e76b6533b2f6313bf5fea336e6f319de9f666f7293cfa01589c983de28c1e5edece401746cd030433e0ae4519809882dd904a037ef15772134d31548637ca7003ce837;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d3c950c98fcfbe4d4959ba3cfee6475709896e77ba2dccdff9360ece281afff999aa9855dd193c20afb1df279382636246e626cc004aeba459473a2ee41a78bb1b4046f660d2b87bc881a36f0328a4bd559181bbf3d7eff13c26779f726fdf2e41b18bbced2509af5723fc34a27df761c8e3dd4dec3d98a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142c3bbd61b1f450285d2f03911c29508def518576346dafdd5ff9e22c87a663b3f48d125a6df89f3b76ee4e3af9916539723aad3d766028f2fa6a878434ceed052573b32221abacdf82c67f49e9ef97eabec61c631c681cb7960951f12e78efbd81a5200b182d67b86bdd3d0a8389bb3781e2f56f5ef2147;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1688f1377a7d8408caf441d850a99519c6c827c8ad653d43f01754b71143da44c2da2f3fc3a18023b026016e44be3e6c2f8e19237147936b84074ace35726f1b440972cecb9eaf1fd02d69968b92b311b5d062d62d3d1c407a8807646ad671c80a9e566447013cf3ad62355a31e827ab91c1bb3615ce9d39a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1e4584d68d1b62c21b0696aa6f33c81f18b7c68623205d94964e476d47e8f4f4dbcd82f16383c285089f02d77a80260d182962511e3ffd6643ac1f9be708c80cc0d6991793ab95b073858033b089ba9fbafe8f2d276071ca6a0306c63b78154978e36319f2f03fd531bd4bd24e9d661f858a8bfa9c31727;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a80300bb948d3ba4a1fa1d251352b9c8ebdf534da8aec8e43ce1457135717bc6244fcba187a433c044fc0943c4da08e5cf7aafaec85cf8048e2e8ca79b2a2a044ddf8c76210f30127874389ab18bb1ebdbf5b6560a3e27df5547e881a9719f773dfad9f8bce493b2c2dff3dc31b603c66d72f935040f40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68cbcc48e0f55eb843598a546aaf22ba0169150c80bf523251c0155e9ee1a4b8df81a37530647bb7fe1f341a84f47d9c686a4cd4be4383b2711924959cf76dd44e8423e93b82c7c5cbd64267a7591b52a18fe443c2132df31563d083b8e4ceb5b044bedb30f8d9394bed0c5726239fac257efc4074b21af4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b5836a8edabf9054292cf065cb165e8c14802fba2660861ebe5bd6d787a337a5a4abc61c878c4433e04b1873c5900756bf0a1e040d401e7ac558c031c69b54da218fc774822326dd8b5f7c275c6ed00deff97d35a3a584da9909e480af672784b93ae64f47140de1e70eadbcac7714121417bab54fd93fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b09ec2444219dd93f8d8d0b38d61a2a1ab5cc22c3a7d6215aa174ab7e0e0d43edcb5658ce8a7c52530d150244668a2e4d6f5f82133e233afc5cf5c518f36beccbc5596fbba77800da2f50e72818738b7e486292c9694a2db161b23b2e66178809bb7260f58bd34edc39ed7221a47e900336d49da7c278178;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131565c90edd3554afeec883b2421e5c0bdbe24421e1b30ce34f24518abeeaf17b4e93e3545c69624068b66eb19aaafac554c9cbdabbbe769676b12931ae25db923ef3bae2fddff625a66cf1000926f48f0c7776a8302c16b9ebc24536cefe8e1a1f9c575257dd2003271455b265b2f4234b4d3363512cf2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5460738886592b214f0f06d9e2d5c0bd5664c70ec8c5aa7312fd758cfda56bf98eb9b47b01e652b14f22c8c7390ddf250902e9f29508596961a3155f58b27c4ec20e55f2b4df312eca6b4895da6dbef5ef7d4d26ff7e6538d2b50a11f9e972b934514e25c3bbcc36de4ebb2aa4338c8dcf038d365ea7d6aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35a4f873f28aa80d94dd1e9e8a0683113991fc2236f44adbe8ce955897322c40e121a2c3e7ca96e7b63389389f24496e32391669bf844e5ad10d69d97738a0eacca071e5a09918150742e6f8a2e5e6c16d6f6117d84f730c1450a85fee0d23ad00ec7f24b90ee69ece4a302d8f3aa6699676e3596d2320fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h944139202e0db36b4ff99b8555091c065ed13e15a029840792860567a29785a959dadb301ff6dc03d9b5ccd9176f74d064ac5f0de4a8ffbabb0d01eef642d01493fcc649f6271443c51f0a572b92fef79390f877e4124d2a881883cc5e771a9fea2c890f6bf971ea4f959620f45234b2210791b6d099eec2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1489ea166d1972dd39c6f22b1a8775014c60e692ddd287bdee283b1d92b51891669d9f0100970a0c8452972fbee27b1b66d3194465f996adac31ea54200753ce757a129c67a17eb2c8220a740951961b8a1050f5c49dadb5be9b3a2a9b103b4ed2275e9f550ac4183404f4463732ddeb86bc13a879067e61a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7ea00c1aaf5321846bafe0d633c630ba646ec30c8813798e4c4145a0e5737eddb4a244d4243b5e3c220b5810854d183564844b84f8fa77f648e1c07e58cb2ca8b18d6f4bea6d2ec7f1cf5acde4218ee485a5e093678d3ee473266d9eacbcf40e6e9919bed145cab9af6c947c346f59a3230f866a03c1757;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157651e246f2ceb110ebf05c160d3530a09a7159b84be914885376902bc6b2a9fd9977cabe774c5ef3a452372be9c8219f1c0376ebd684a86399a297712fdfbc17e9da28cd3a5d5e7bdbc8f83aaee3ef09d53be7eee8d6216fe1c282c1395b81c4100c72d206d7f3e84a43e6555a998926d6d673f5e5bcd0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f6efd9088a08913032ce49a15cea444b49bedbb559e9b66818045750a5d65c47014def3c97bb6fc75650a271843fc4e704d5032a3d7628cd6894e9353dc068321b719c0091db58275efbca28297a697365aff157366604baeb2d7a7102846f136299a58baaf41e38de043366048cc17776470247e3e2ec5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7db173dcaed6368e2d4bfbb62a20bce289fd769655b42c40fcafb2e0ccf85ffc16ceb1b2c0fa5cdde649dc3cca2a9eaba03d7178cc876e05ea6b337bc760f5580c0a1513d18034ede62ce29dcd0a4ac00694261f080f00325f362674863c61ec62c85dddfae93b6acf4fced3ed66423243867f6953e6ce10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ecdf5f3a4be8f8c882dd41faba84da80e1162233fe16eef17321a5112421579409e306221a587d6aeca96d75e54e497447188f230f842524d317b3f6420cbf5ce8a906e99bf06be12c81add2478cc883099bab119effa3e1e75461b425ccaaa4cfb4c13ced07d575b785d183f919930a619fffb2d99d290;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ebc0d6dd618e027fa701869d1ddb2b9d0a7d7ffe5ce46c9a5f5484d9aab755a5861ca475bed1d548374fe355752720970ad3d600441ec52cfba11789d8fe75268a58d803949d54860304e4dd84aacf790d12be7d7293e02c8055a4bb78e4182f678e3d57ef018f9c333006f9ef62286b2e816fa398da2bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18472a4d09e1561322af94921adb12811356256e6c4202a3e19090cfe3636822f01531c29913ce46595777df3fe0dfbcaafe6815dd7cf56361ded019f41de1199ddd7cc72f54e59f2caf0caf4c6d15593791687a319b0f454fca3fa345fc389ee02b2343db429fcebe4123cac8ddc2b2eb89c5aadb9a79952;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee6937f5b18d5e43fd66c3e5623abfac6ab0611892edf8aa6b14dd59d42d50b5d2479062119bca7be637416f00d28ee18602d9560114cf03dd08e1c24b770edd71d67b08f9e4d107e20676c36a33a946f5e763426fabe3e9512394be36678d57629d6a03267f9437adc4da729e0fd211570b879c3a830f09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16434fa93ba91383ef86726a28e75ac75370965b055071641555d9369ebf3f47b7be21a76504332d9b5eaecbb157cce6dcbcdad68c5750f8255ea6430f0025b7ed0b8af524134f484f727536dcc21668a6c908786ff75d659e21c6f385c2ae39c65a04236887072c31fa2671e7b52c8478c804d7974aff567;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cdcd48ebf53cec45026e7a96a171648ba862fe5d6eca6103d492be7a9bf53524eebf9a956f8ec763178d71ae60d73041383c59eb7f3487aa39a697fa54f8be372e52065ff18740f6528edf6ffa9bc4b2be36361df9713cc1431a4c6821c59532605f0c776e895b7c79b8c55515a45f508756c20290efb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2d55b8d96736690a1a4696313887c3c0113bd763e20882496221a52bf45b4fc586489fdf341b67f7dca54a0cc9919c53ac312c98045447fa1da82536237b413782789132b66d03ab948a9875368b93f97b6331e7bc1423bc87d69aeab86575b50b97da4ed0c8534be6576c5a6c2a696ddb49eb810b80cbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb064593361a4dbfaa87abbbaef2083e409cde845ae1841e8a48ced36c38a27290ecae0ca41d632a9ee09db2bb7504ecd158bad396a782d403f14fc1970adb29c5df335caa7ca91bda24294f5eba027f4e241a81359698ad43783385d88c86d8c55d569acd63157e103fea85376fc817024381c2e7c17b2b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf38a08e25af667b1ede9f8397eb36bd6b630a8791fa8c22ce003f104035b1825576957d318d000a2762a69b6bc659c88ac7873356b9fecb04b6d6f9d8c9bf37bb62a96b6807a030a4509f0249b08ace87e1c72e9e65bb6ec263375720e0cc76ccba022c9ddc90c24c8c30b6640ea6f35c884a4248f0ef136;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e26a70de193eb65afd1e22b0a8fbcfc79b0cec053b522b05e1424972b2237c4438def9727de8649814ddaa608d2cc2f16a3cb68f6f75b582541b2d91314e7cda1c8a912257552ed5b4ea497e443a3e3645c2c9c51b18e71ed726445427b78918050d499fd8f8ffd34808cecd76a070dcf91f94e87160024;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4fe6cf77be3696071d02ead63b6a5d1d6b58f85afa7cd26a76eb680fc6673447ae41b9f34cce01585411d6c41c600a840889e19bee5db2a6e30163a64889ef7e7f260736c76d4dfe4ae0d571229e4e7d7d808681bb7e905134bfe4b11520e8d556f23f75e88556045f62ca1ebf9cd77133142e717c43822;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha47a173135d918e57766c6b876b3de3659e42c6ec9fd234f5d06ca199c6db72673fa0f51d049ad94ca2f89b529d904313f5d596e2088e8a6aead79e5563b8de071ec1eabb746747d20269547fe49dfd989e897178cbc4788ea6146254de4d3592ac2594d75a5a36c85ab37bdccd3bb1f4cb31259064e2963;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94a98161a2b42cae9b39c3bedba87f7cb7779345be9e76a922be7ab0b7dbdbe243cc48818fea24f3a156b11fde58792b3fec9e7cfd19134b7cb06451ac9cfbf9f3a2396b38dfc38abf21a68b040fed513ad9e393f5efa5c684f46bec1fe4a92a9f04d2b3b034996c56bb3d52ff5d4d0f1d41f4b96442e2f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136f49afabd7165d1172dd12809768583875455f99218f06b8341179b22a197584e65593b018fcb2841187b476b3cddd28cf79274b52df4370c280bc8cfaac11ca12e928562c41c6d3da0899a07fa7dc83c2660454cfbb351bef0ca99c2ceeb95025446c8ce33c1a4ee6c88e98c91e4572313664b21f877af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafaecc9e5ea519c3e248ab5a0d5e593a1c71355099fef577e390b6522e9c57c39330c1f4ff46ebe4ef0b0921b9e2fcf5a1d793f74d7e43047350ee1fdaebc8f890e693cce2ed3aebd19d3621ea7e6c8a3c0f3255b17845c19da67a05d597628296ea35e02295de253298af5d10d0201153c66b4af4939699;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5afb76ec76d2f69da4431a62a1d65795170e37eb06aa14cc98dd31f6eecf94836c8584ef0d25f2502d0c7167594bcd1d6349750bf1f0b607fb2f8e6af6395714a501b3ba5e9d882e003a498c951b944b722d1da30c95e778692a0d0cff5b4ddda0576157da47ad36967cfc447c846930b549e49cb914316;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1beb22e36898030aa09c37e0114222db65ce9bf500374cd80d7345f55d63d7355896c4994e740c4b839840ff8aac46138546c78584469d951ad290782d10f8e0fbfd5ac9f39fecd26e277852fa2e56dba733d9b7aeaebcc8faecf2036ebd3d382dda325aae90b3fec15b8deb1b623bf667580ab325327a1bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e52f02a0db5664b46077a30c0bd1805516585758aa6550e67c83ca0d9da609fafb4964a83cd3622e7d730ccdfad11e08d5f299979ab9fc07e89afb8b16c164bd0e0c3c6d74cdece30728e26baaf6850e08c26fe547a5847982b755fd0bb0ff9bb6b2b10a86d5ac79f234e9977212989e3ef455c6856feea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d63a06063bd8df022d6e0579530dc7fc1399c7db187fb784f01874f284759c41f113931ec0f19b3489e0f4ce167ac4e9c9c490e47c91705aec022e92b714557d0657561087df5725288a11a93a335583e702149d6133ec83e2fa7121f865223fd509730717815b5c46e642b09490cfc68b2f1a0ee2e4c33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16650e2101562bec3c6d52980e6ee03b5d9bef940918babddffb3455240f4095d57ba678dafae4843266218761cb44eb7f5689da262678b2c5b14ec7ed18f5872ad67193ccb2d134ab6aa66aed2dbb9bbef23aa7f3f95b6c79675b37f4c1fda9b7701d15d7f91a87282695c4364cc6e044ef945460e3e0afa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h378070f035ab6d937593e7ac060390f039234bf836327162c2e13aea195a461ab24eb86772d88708ab5aa05dafb008461375f12cc5468e4c8412b82c9c9fb7760f14da7cb6d0e3690460c0cce6962d042156c60b566171b2588f7d8ef5da7d1daf4516c64da4499cb2921b17d5d82dd2916851552cc8c6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cea95ac7f1e93ea4219e491118fc2692ca7c8a22a8be843932aca0c2302ba4ed8f2d8cf3d59833e03c98bfc53d33e5470d224ca2ab80926880578633de59c40ab076070cbb47c1be290331ce9343ed60965d3082a6c170b6bd12346b4c76cf5b983272b0d2052f74305d242b91ab37fb2b0a26552d85bf0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f1196c2394727cfb13def892b56ab692a40ed6d30faac776fa58aa87c9792c8d897917097fa626dce2c9b14363b2c96222a1264296a1b35bd3a0971eb288258db9ac9f9690ab676630b1b06823b63f2b711158e064c94c5191c624c1a133e16d18b876162d4d7481245b820cbeda5665bf47284b18ce51e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1194f58dc5031c470f5ea2a05bcb3d125c57bfb1fc0bd0de830a8b6dd4ef8177c0e60ceb061a55f4e4c2abf4dc8e250b2bc84fec77c473ebfd3a98f8966b538346728556ad4214f4c7684c64de314ecc870f9666e4e88566e4529fe6eef7a247cb636573a8bde5c508bf8cfaca4025672915b0ff796908bbe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f42b6dae4284fd8db3d047ab440ea68e0d9e957b54bde72da6637eb0620c9bbc57608a97ca0243dd4850688e6b4d1883654b9cadd6b50904830584127372585a9d05c43716f758d0e7c257c18ee92d40bddd178be6e147898c1ab8c3ed69844a6c0ef37d0c1528613e2683f2eca4862abd056e50f2edf2ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7052ba561a54ba7af7ecf46ee4deb6a1ce851281683d6d6c67290b020da576880375501003314dab3000b83774ec2d5b2a7bf53f95b98a2a2a4e518f1558c97aecafa81038abf2374b6aff259682caaee4ec8ef537cb23792e0f8410d28b5fd2cfa4d4d48900674170b7aa11456e19db7b70496b35a386db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1145133ca394b4380e6bece4b29e8944312000a3b75dd9977c7be248bee79f3a3ad5cb9b4ee7bcd28817d49f2b8b8d832205e7a8211680dbcf6874306fa61593d34502a48aea725b423f923e4ba670611c886d7c1943566b5ceafcf9f2def811031cf36bf9c0b818e4792d9a73963b7441c362e902596e772;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ab645e8155bcbb375495e0a360120651ae0e0cfc4bf118ece97f6673c1916e743921b51bc0ab2d06b1c23972647d1c41ba18442b67cdef39855db87296f462f4e145dbf66372a1484ddb67c47291b5df9f3c88353f926d92fd2e596ebf6c0e480ecfb8c7fd79a1dcacb884e92b985a80902f85fbb9162ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf08345d4175a0913f6ae15bbe1a1fa0965864e25dc5107c267745690e53a4126c6b7f57c29233d949f9889f487d4c7e8af6d30ead356974b57d0adce76c458a8c660c84ae17c83692523213a9d98cc340b7d12a899d1cd040a82e27a0ed879f21e96f3ad925711730919f7b06751d9775f417c6e3af6a563;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h641aede767b2d98510dc24d83adea33a581b4fdd62cc426964ddd9d27c771ce30f3f2e10cd6eddb58ecc4cc5d34f3c4d3428375230e189fa5fcc475f1f2321e4914f5df908ff6d3ef02ee862efcf60c313f4264bac77e12b1412c947eb698a7c561b85db84adf649441c459956eabab2a3fbb816c060d8fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h868dcb0f1e8bb2df684d5eba3919b9ff18798cb5bedc77b9f313f18f00a7d559a68be040180ccc305b3da575c629301c3d1384e427da665a2d711aad788cc1e299b7aa4abc0918ea3dfa906534ae17ec8c7c0170bf864a4a5919d0aeee6ba2a25f6ffbfd324d20e58853b19aceb13562de09ca4962985dfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h352d0909a36f728d2c826ae09e2ec360be8cd91b550ea35f80c57884ef68a1480f313c49d6c0387ff002c582e90d3318af749915c4bbd13766243bff0ce88b743f4fc755a8237adf2975cb1bac59935e24dc9837e7aa37532f2475d6a2ea3f00e89b527a3e7f8f62c73f4e7f59094eaff80c24c4901105c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h159e20eff3d18dd11495b7b4915103c6dd2c53104ef9c379d22f676faa9f44c7eeb0e43e74417af06cc4dbf11cca5ae022bcc1b68ce74f4b93a915552ae70b1c0efdf55fa66603115d67beed3ae6e5b75e8c3d9b11469064ede8ead6ac06aa73de429013d00f5339e0c590d13ba1e0c5eeb16a1c55bc66783;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d410a0735605e5b7d6a60f1c7e81a16037d8febc7e587952592ded1a31f6b275f98afed79ad68cd56cf10036d8cc06917804607e45a3e3d4669456275f9785841fa5b9cf11d10ead8e4560c5b286338e6c0272165dab6c9fc639e869b47176403e429238e6490667643d87569cc6b5edc969dcf630af0dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152437433299779f5c75fd9ffe6f073352def43ac72d2fffe076f6274e0c10b0f00f0b45e24878ae59fceeca5b3666f9df191e2fb86638bfd55ccbb682cdbda50a484db9f45c76a2d6b4a506f68bbfd7f092b461232f97276d2c6a3ef56b94e120a279181f2e725960a0041cdff817cdf66e1befbee47dfb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e84f8a56d675c0cdc527c5dcc8de5e7cbc8e99223bc6b8f155455742af296ef3f488ef58faed1d5e833e851f564f549467c6c431915bdc474fc77dc3a8f404f74a20c2c384722cb7eed436d5108fc68e22840291dea5120401dbc81baa810fee531b0b48f60b8f2b91a614b075dc737d9fb4d8915ae39b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a062531804ef448052051322de4f9c9a9d739e1a4b6ce4e85104a53f8a82a8bf419a1e5204c9c64c3fa3bf82a6d1426ed011c1dba856cd2662d3fbcd17971d79857ccc14ac3923b07e1113014698369468d34bc163845e2412d2b0cc8517879652c5c68f03715c57ef83efeab23d0747349c66a8e8c9fa0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6444bf046991aaec6c707145d8ab7c2e818bfe691a56106e34366b146a4d803e8df7c0245de142308e6758d7b629c4dcd8366b0c515497a2b77c450f7dc5427cc4d8a7174ee7f4d04ce1d33b9d3f0c4c5fdc635eea0a482d709b907d4ae6728916d25c0b2fcf80c35cff4fd87ea54f6a84ac71dc0448f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b174cd63a2cf17d6a69694ae1d6763d4dcf35dbb7152723a30f52366054e86d318516b7703a6358c66c2c6f7c4bc123d9c4be9816122ae79a074ce440ff1159978cbb6566afd9968aebfee3aab396499ab2d1ec0404fd5a75a3d97d5c317d396789439b67705ba307cfdba25702bab62eb0bd2c002f1a1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88cab4ccaea316f8ffbfeac3ef0ec4f84186e3f59b93b08b399dbf80424baad4545cfc6fa328918d44a210b2a7c2d508386354b3aeb7290c9d4fce8735aa763b9ef07bd81207aa48cbd03a73729c013f82d899375262043a97c96235fc6306e4f63ce7158355e9f29b83ef578951094197907b4feb651500;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa8ff605387188f7f98bdbae6909e6ebef4d50c95076c72215792e331150b56f1bfe560a351fd9f125b0843017191c9cde3520313663cd18ee866fd571763c12357e179012eef1adea56f1b181b573001dee3732afe7671c00dabb7dc8d496c8336b6787581b6dd9e6cbab8a6acd30a63e16cb6162d3ce22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad35b67dc783a1dce6eb4a4a95a10856f0a8a27ef19b381229d98977f2537a7aff159eba319a1dd338c2fb0ed670596d4c1616d5bbcdd923a95e19f56f07992100e32aa06dd33498b68f463b00dd5b97a3571c0a59088e1f8ba305f1c98498eaca22400987941a1193f073e481bbaf3020bf11d7a8765508;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169ffa0ed25a7bfae6fa838442cd32ac90db079858f19b71c83eebfb42ca5237dc1f0d44dbf4ad50eeff614cc0fa732dc4f75a0491b91e63ab9d79ec9702ec089e69d9376f215981f16745ccedf7d98e80981b1cb31990d622c35adc5c85b6787c520a7997423a9580f5700c05877af71e502c0234b00f622;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e026fb20706ae309d1cbe33d4fd617b79b92c9c3b33717ac1a612b595d72d3852097c041f5e050231d5495e936fbaa793193215997c7540050702532ed4583b26be11b9c36d790cba862b35d7a7dc23ac097bcc32bd972d3753bb3bda2db8a33dd34c69d7888d7965ab9586cefb58805376041c9b832ff9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23e4829134351ea9c7f99490d7798cd8a1e8f4a77e788289cdece42409faa2572315e49e43a801df4b636e07c607cc2b5f603924d619b060302260ccf5ec8100bbec3d408565a6d8df8bfb775f3403e77f3e1554b508acb0cdf8b3cda537b7af5d34d0431dd9f9fae373ff14ff11b7a97639b6147e39d486;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a97ada868a33ee31d2c9fe64e70021c9068c0aeba8ab72c1f5dd14fc95e17d0575bf2251a3fe15d780571d807f6c712a67bc2e3c3f6339e8274dbddad17e3ead6441cdfa6b8626e1e18278d468e0ecc0db5c035b12e045f586b575059c40b7a4b466e390939f1efe676992f093b3d679d416c3d81630885;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbf93b204ef8342b0d52abc937c916d13ed37dcc9626ef35eb4611add11d04309ff58ff0e79faae876a68053e63a79c2cb44ed1ad7da32875c12432244fd246193a547f1a3ff79e237c43f878a5759387f8fee5e7b51d45c4181c63b06e1abcbd819ecb2897eb16e311d9778a228b676a5eb6cf6c200dc30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64bf0d5f05aafc01ba95d8fa1b6af2ab9e15c384c591aab9917d9093a2135bd070c85103961574d413e3489e66c823a6e7c08503ed26632b3a9db293683300321fd0f6fff194ea41a5dd66b4fc3d66b3429cf9eeebf1df396d6b1307d0d546cef2d12f1bd46a839fb76302c2b5262b779d862e7854dffc45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133dbf782eff7d4e29bb2faf3732e76663f4db22143d4c42ca0a4e793f44bc9771d7287f95653a408b32ca61d3481358983d77bf6408f9eeea88faec7bea78dce6da1a86fcbe35990900bc0d8caa9612fd3971e9f9d5472b78344dbb221ff84621620d812d309869254060effbc0570768fb7a1e74b363ccd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173c9b77b127dc19aa86e02f58190ccdf368f0aebe74894dac5a00cf1ede4105b338800dd6d7943098d8accb35101e0c13580269d096847b1a4c1796a5247f509e9de0721c1711909d2b3a59cc87de96eb40e4273afc26b2121cbc948b57cd58260d8a5c802884b3e948b477c97acdc6dd0f09684431e2b94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he83f7bdadc774c4516e93ee176493c2d6fcf31a7e58352122fcf35ec453c091ad8d21c04c6dc0df3e238eb36c9a93ab45a645a2af7feca807e1d11259548e745e2f89b234faba9b591ea628a7bd29885e23f9b0a7f16c7bcaf289498067c3dea3c01538a2ae94a6cc1d589c7a867f0c426349d60bbb3d875;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4fdfb929c86dc9038ab54195fc754d1f9493c077c040bda5e2f8e4c49661d236b6d809d1a9b70df49754bb19e0d97ecce6a0e389d97cf2ef837ce27cbc32b318cb50bb9019c1b32c368702c090ebda8962488600e37ea3967b5282b55aad5d72aab1385e8135caa71c61e4a9eff91047c4ba77a66310f4b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35aca35305a6ffa10f336e64b9b0fe596b687714266e48082089792ab730bc1a8af2e912fc0f933601ce1f5b45bc14c1eb8d0db53aabf1a551c29c446b720aa8a1549b9327a56cbd8621e025d4a8ec42954bc33c671a1811b5cfed7e66cbffb88c8cb25170087638a43d7c19e81b45976fab1e4138805cf0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f2c9f4bb9659993359fc95e66533699ca4f2c805fcfcda245c1e7edc2e0b986ee0df5612d89fb46bd7d8acd26032d3351c8c32855a7fd713cede91ea1e04be498d52d5217dc00666d0ce0271bec0a7e581562987dcf91dcdf167e963d6bce4f96974be575292527a9ff21e2dcbbbb8f3a2f3ca39d17c94f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b63d19771d4e4d6b82b491d3565110854d74ff47d94832a954d1be93a591a58873347af717d26e4122db7a86d60367fd7fdc46c1fa32ffca1c0577e330ac134ae83fd0091ef6fb3d8f16353c72ef17fbfa41dddcd55c7f42cc8001f1c50cb3098004f0df1e43f403e1f3d37cffd4bd1991c183d50df2354;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d122b34c8c544e16a03312c230de13eab01573d060714303c9204ac43f51a62ef10a841c6a8eef6f8bb32d817d957425bb1df19bef983787c34a7eb60050942d935cdb204b6cbd232e9a93f25ceb1058df9949be915ba14d936ad246bca7eb04bbe3f758b343cbedcedcb8099b431d7e018234b559c8f6e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7e2065dc6eb75fd58ba79754bab24477337ca034e1079c23e85cda67e8f34adda5fca41829a97144171440c049cf84c466b921e73bae0d9528612cd45d445f6b7aede5aa1dc6078cd039dfd99b304804989541332cd5f7e10f56840af61d66fd9071ce069613235adc565dae7f41f2b6ec4758f460eba0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9690450e307acec1da68eb7d283d1926384eb7051bfbcc1d13aad33b10332e8c45b9a2880f6a5bfe8c2cdafcb1af0f7c13a0052b7a72c22ba6351720d7fb63a97528d9381bd8ee806ba29408a25eb9271af755fd4cdf60a42a2a02b24ca4d4b448bc638545a286eab9ae4e5a4678f202559a2d2c5d2567b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9920911dfff2cca71818b626bbc5e30d00e0ad5a8069e37fafdbc468fe9be7fc61698f7461329c34ae013182b83ac683dcee3890b61337908991648017b3691324473b90c118d3452bf30775af3fc8b5a7fbb7582682b8fc0dfed4c01dac73ef8665036f583a467119ac271f35ab1089a101a104faa450f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cf3a16873bb632daa89600d39b3e52c9ea3f45baba09a487dad85a10e7184b51e7ae2b810b9fce3a712e62ba1d3d0782348fc1b510903ddcd05c5af2bcfa3d214a9f6f7a66337da04b997febda46cc46bc6fac27a2664b48f27eca73a5798838e9893e1e1fa380695833a3beb59994d575c9d1c8c71bc5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d061de39e44efed8e9d362f4b971ee805b07602185524f4585cc5e53c7c901bae57d75a6f56b5de0052299f5d84ff3b426aa53fc5da6808aeb2f663f3c2260f35d01ae4aca136d40f5deb7104c4d99ea711951d94feae5206dd8ee664467264868ad54d97a651fc1809dabd39d9613e977600457cb702ff6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12dcd523819006d5f1cd67d5d1c31635c60f46af72ccfee8e231528dff3e5be3a9ed2e0260c66e6582bb7e86b962347b3ecf5943f69b7f18cf8c8dae67e461125803c30250249ef85dd46eb0d1e77974eae07a1ad534b49be7d956d024ac51072183975baa59bbf0b43a8392e9cd2c637d74e9df0c91e22b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135ce87feeba25c1c9e2352b7d05a2ffbf5cad6f13b3c4af5602c078ad69c1f0c194faf019a8ab585ff42252469d0096f6b89da6a805ce7390c1b20c1edfde1510f5f0db1c30e5c9f4fe482d90cda92597f975f2cac003b2be2f057b65161a81dab4ca7269b2fdf0fab008c05af4e469e3a0c816e8f1c6742;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190e53f244ed5b18a4523614ccf227d40cf0e41fb6cda7c5b6679cdd2ed6d8d18fe055824042b347c16cf3dde3236d703cf485aecd5bf39cbd9cf7e3839d30ffa6a7668969e0582a18193ba273b490c3a2bf43762bf99a06367bf131e0b45aa3429272e3988fd869e6037e82b34e3b7f30ff93134f58af293;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h700cf0618ea51f205248ea657910b5bb044c57b00084b76d3c7413ab88a1d52ca910f3d1119bfaa3947b4a2bca738a4345b199525915aae49911e8e090ac49f83f01f9e63e8290fe9afe08c325a15ce6eee1d6106173094e0134136ddd46e2acacb66996dac97ee7cad517c51ed2bf5e90eb86f625e74dc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf76253497651daebd4e9108b718323cdea42934cb4de2cda5027217468de884bcc63c67c565fd2e176d12a9a6c5df4e8a51f34da4a9ae9f5124cc02fb832ecbac6d8679194b9229ead64c22a473317adcec8a37a82cf3e0ea166c9f9f322641896ac3df7b1d81f5032156ac42ea8c5eed787129413a6e5d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178c351a2a4df6fd142556ff6367d7ef0735472aba7b5b745a0d16b4a26d4363b67d42b393794e427ed5f91bee912b71fd33368f39fc93e2938deae7c008a2afcf5ec41ad58ca386a48ec9a590edbb957436a89ec85672ec8453489b1e7e785d7ca6b3db9e5520b3b9393c5e04c11cecbe58b32d75acf1123;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcea88b725caf49e4e756bd77df229b27d7af390e27dbea6803bbac6bd00e3932dd88acc6ebf4de2cc1af126bf0d7b6d4b1bb2d3c53990c407b7ae5706cd39b284cd233bffd32105fbc4340778596daf98575c92129ee90491ec843734cdcb13dc7370fbc3fe8489d779ab6750dcbd37f6a0fd94b646e9606;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41d45c75c88fadf3da1dbb9cb953880a3f20641e004eb779ef30699847ad3cf3d85b5b11b827d7ed3258f169e9682d82a1122389fcb544cd1ed3709e119963d4fb47ea39612b8293814a43be41a72c2680d5c08b75f52a063327cf7043013bef8fdaedc7f696ba17cfb9235940c75cefd5870adb40fa292f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ca05bc95ae3ac4dec81f4f3309e5d9ebd9a6906bfd1c55a6335999a96a68ed25064d097d0f2b05148d07978798c530e9f71abb203efeb6a5b4b6fb86b1e0cfb8821eed4c00d10da3b2d2186c1dd895effa2e9f933e88cef14c95dbbc7b5274d271b2a7bd9ae1d5ba06363f5e48966ea0b281fc06d8ce452;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8279483009d01700b81a5667a996df25996769ad0b74cde9c8890eb5381921b2fbc87aa4997310ce6ccfc283122d2271dc8d7b87ca6a1738435277f237c73ebea772995d5fde0d425329305e92f0aa866d37ee9b7733c32a61cb58e1b2eef672be20135e37037455568398a960913acdf2426edcf23dd2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ae2753fffaee489608b821c7335728674a5e00fe90aaaa054bdf524b643979f2b85fcd938ce593010798e19f85fa2fc814c06db1992f306c4c1e0f139d195a1bebb1796aa7dc11611b240347888f273692b0f6d495ae73e4bf8d4642ab097e71b66d77bf391d83fe12c7fb37c1d533a6aaa675d73af1017;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9bac1fc50090e751a86efbe621a661474b8e32f1272da0249719c582ee2d4257673e8111112592c01457e05add2b9f1c96221a589dca28dc62a0430306a2f9492099a7b4d1df8a6878c79a54f3e6358dd2d087972afbb23a80f3fa8236ca67da5bd5eefba3ca797061f6e7273ef08b4ff59084195bcf1cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dab934292c5a7b5a3de4372885fae3c3157f313917ea30a2b4928b9dbbf1c76500133f34f8e7f7ea9a3baed418fcd3b9bcb9d200a82a03fd5e34c0b98fc1a768bfa808d27f4c0af2d393f30717ac6f9d85e1ce0a8ca6fe1bacfeb8f33c5adc412fa09e0bfa7b9b4638fa81e370446cad4942ce179b4c03f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h251055c6282bfa57228028384cd3af8904fb28e1fa31bdd53c7e13140fbed8e7f3b66788ac60f442ac902b69393fca90789fc5e2afc135831f07b4de8124e8e86cd82534cc7d7969c1e30fd5bfe4a3bb927621fd406d8e71107347f9be73f7f049f4f67d5d139e37fe046f9c6c4a488ece93bb3b8f28b8d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e5e2c6dbcbb5742d4bb97dd79446f0957f0a44a935fb2c2990a1f848a84e74b3e914da48d868f4521622117030440f7a544954f98d1ae27ad9cfebdb1e3d291ddf74de7d3f2db10e2e7d02f30a6841dfd3f22d8ba757927219b1a545f94d8dc73e8280b25baa94780f9b456aafb611b9c7968473a70eae9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a676508dd2c193295e8e4ea88d468dc421e4d622a459f00a34d174f62f7690037d544b5406c50839274999b26b1dfce3d517c1a91c9fb044819fcd77310778b8d283e2218b726d9ce9095e1e425a88472de176817ff5ee428c47f72a4d6978f7eb8e990db629794902ce7ea0f3560fb0edd6c4b364c00b2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f200a6cebe9759a5819e76fe8ae4fd0ed2f4914944d64a6a7c82012cf222774ec52d19d0785f28a2a54bd816237cb3f4546dfb35da35a6ffcbb809213b4719f1ebdb815a7e89321332b55f7d3a312adaa3d6dd175f4f0f886d97d3b0b95ba525c43906d09814afd75ad3a521a512fcb6d18f95c096c0b09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc90b033a9383527085e138aa5907e820d3c2f7ccc6f2fd1284569979b377002d44099dfb44d37c64aee05f9b4767358f77b4b14984f1a3888718d1383e204c5ac37204d0a93c3b872fd716a84ad598ce0ea420bb8f048a740c39c4294927623d3d7b32c97eb3008ceda7c66bc632312b1784b3aa6d3dea09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c33b867fd6180ec98e9235d96a532661a64c1449c8cbebff90fc470396ea378008e90a66dec48e5b932f185efe15c9a4de2202580fda0b3c9d604a8965aea5da2851788930dcefd09a811ecf853f016c8d36370faa64d75487dfa0dd231d25598f38b6af11492fe3af740fe47534f68ace7f767289c2da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5de74b7b906b50f28c5e02574fda29abee697842bfad566a723d001011d962d072d91c9bf6e43c0e872f9729b845b54a858735b3dfbb388d98a69efb285bba8b578dc1aede708e9afd707006202764334a95cc624260cebdbcb6e6921c31b01cb8829d4a80d86665b84673c79809e486e83ed42ecd4e74a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b516bc0206c8f7b7cfbeb1c3d179c3f3377085eb06ffa86ae644ebb8b36b85c5e65ee75ca323d4e812dedd69ded0a996e2e4a0e37f74832af3b28042584739f9ead31c29d672fefde6ae46766d3b390b58f7202e6dcd3f62664cf9ac8a52233fbd179dfbae9ab06fd16ed025890f2758c94698078933d61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb3b510b7f907bd9bfec5523ab7c94413357fbee0751400cffe28e06444f23e4f0575ea4dc683c8e14d4e3d7d322bb211006c936a80488016df72a8f4fb7443b4aa7404c5a15cbfddf2a66fc103a58d47e6272c625f49ac89fe9928a6fa86f18adbd1832f812bf06b139c07afc45d40d40a92c05495845bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he36065b818ab3f6c5bea1451bc7783375230529cf116f37e69e806fe0d439955d15fde991e5ed4c051ec88e740dd933f2185c4fe973cdccc29a5a0901594816846e43cc0b597ba8fc707094e2cd77949e5b1f4b12123e5aeab45d090ab63cfbcc361115d0c8b5b524c1acc70df65a42217870f111ad831a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0c5d0654968270197e2dba841fdd6310593d0b9741c177cafa3ed04bd22efcd58c38d80c6e795f9b152044f54881a7e49b017f1693170305c1a7f8c6c19740eec6005efc98a74733b8f7bcbeb6bb54289975b64f09951762c484f65989b7151592fe1a06f3d0e20d715d7a6d9f0916619f6dc9f2efe028d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184aa65a167320623bc9ad3d3f35a85aca6c75fb2fd735f49ccd78930883f20159c3add4eec9466a20c9870fb82c148bb6a2cdabacc87650521a4a6dbbb40b499f6ee0e0e5553a366930125dfd86cada9cc6baa8a27e4233810b956124930a81881c1118a91f4c6a2af94188934a4ba4e0718d7f8f41a5f8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fc6c9a57e9b6d048d4fed5006648254c8dd1b739fbb33df5421a09c99d284e87495539397580e05bf350c51c2aa79ff55a8a32e2b380ca107d23e261feb6aac557cfa9320d7ea34f1cc105b5a74f7cd1447f9b984b76a64ffa17163b3e2f91f51d3103691b8971158b35ead8bd046d12b9fe28ef89f4e5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb81ccdb1fc4ca191a616db13988b21b6342f99e969309a8cbd6dafc1768b0efb8c29f2b01ba78fba94f1009d55ca30663c865274381b1df9fad09d62c6536a17b537d94b181d13449947bcaf69ed29413dc3e4bf7aeb3481899d8e2099b1177097d7f3caa30e51a2ea5442e819db4f49502d97d3bf3e66d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41d04932357c5dc2b1b67191301f005a51f763d76ad36f52e1bdacf39aa249a7d85a1b8090b06e3d27515360d0eecaf67c03d9a50da162ec985dbdbb5cc571cc6b7ae36e90e0d4bbcb588a9bb7aa59762db556e4dad4f92282247e79c54687298197f11f791b2096a4c9aff820ddc654e25a35f362f03451;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148ee4f3de815d4c7781c6b689faa672725571d5366e8a70fbab5b8ec610f8079f56cc6a0d5eb03cf6501a284144f6df6e8a89e36a84434ea54ae6249271a9895f7a059f91aa03cb073ec6f96cc1187b2a3025697d1a5b2ecc8559e1267b3a84e06366e4de29a5b2ced83d0987d8471c39ad4bd5fe89ed790;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b7f5b9241d1da51f4bed54dcfee47eceb4f6358cffa2219690c45df014fe25f6889820d4de3dae10bc2bd92088d8f4cb5c2f3825cd8036d7374c9f181f7b2f24f3ef82eee11a7aefe91b0023fae64524fe23c5f63455e2ff5787e43df7e4deda9ed6b55fe41cf9fe8ee4236fd2daaa2b328047bdbcff83d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3495188ffba7c8d4d53ec0cab664462c255ca3b29a518052736e714e8082f05378c3249a0571b0777ad3d157a3bc5dcf4ad4116f01188c70f4900a9da44fad58b75d292de9c250491971ee13a913db2954c56fbb3bb3ec2e523d2fb337934c3341d8d21287f40a89d58c916d57924fb73bdef4426d133b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5ddd5c2eaa0e1d66830415146f541cca55964bc99918c90d127a4071dcc595291c4e6f400b0ab01bf6866dec555faa76c40ea1c5a25d8211f78d97a656c5a20eba16d436c1d9a5789cbb1de40837f223d9c3bc72244b5aa514cf52882753dd7b5abd60d870e30f6df2e73a875222d680aff849a4bba5115;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4ad4300c6229ccfdd76e05040d6644d13da07da19371dc51d622260c1902bfbab3e0848a6ecd72f8558b0bf892d1aeee27777b1c0915229dbfd887f47766c439d123d5dd4ba5891610d564d69ab85114d1289451baca470f39c61cf141ebd8a9e3d84934a7857d27a000fa4d4fafb9dde37f7444ce1e396;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dad8f8af7d5972227dd722c423ae018d93acbc75838d5952c13508cb0debfc4966628fc996a16096a02e11878787c8be1ab96765e1c9636b62c438d07aad4531ec37fe9d317050b2a1c4ea29d7a0e738928f14441e88ba3cb1098f6b4ae8c730b175e1e8bc256538db8dc90efc676ffedc608283a5eb1f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0b068e319a853f142c48a1348872a60917d718fa869e70a8b00e716f3b98be8698393e8697e9cb9e1be7e48fc20ac093fe73d8078fa58a819d572c6424bb280a19e1994c936a56c731f61a3bf95d03e30b4f86ce8760176bb47d89e9417115b48fcdfea1ccae2231245085ff1bfb5e3f8c67eee119961e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43cca7c8466a5ee6fcb087b3cff1eed0b7648c9f76e614f73698c9beb4d77ef4339448bba6932d7faa53ddb39a13c35d4fc63d159933807666e68ba36e5bf4d151a43cdf485367f5bb96d4208b15d2ddc8ee948483275dd7661ddfadf3d498bd64c1bfd1e65ad2b0b949da6a00e1f34b48ea01a733f291c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32e1732e01bc82e0b2aff9beff1f8fd1503d13b897305ba3ca522066b7766bf42cdd624afaa910433226631b46b6e501d765a982831828afef7801fbfb6bd9082632625a9ac980b0594ab3a84cc90073614e9885fe43f41bb9b891e7f991dbe595af33b1b46bdaf0e19930027edcd420bc6846cca2b3ae05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f22d89fdfcad40db0c6a382f48b07fd81490b4bb895f67216d0732a864c52a648866dad1f1883c271e6b4dac5a61e412ac09516e9cf832da3386cb56fa586e3a6fd9f655b14473cf69ee1fb87e24d4249ac9b903285e4f6b8b1c8945c0adf93c37463d4ce924d96539f832644cece5d325c00480a5d161c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbfc35247b6ef91a36498199108b4fb6d2c361f6e3e7082600a22be7448bd013cb0a3125efe10bb3b09ea5001f27721129782ac31d82b96aa963a16e6352c4e622e3715a0efc7333e092709956c9516f6b1e1dd8bed8e8d66077c2bcb3b31bcf9891d868a83b3964e1b1ae528a650430998c95b1944953fc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7472510e0ca6ac2c575d164b976a3bde087c661a5a761ce495491cd4a912932fbc5d6aa120dcae2d51be196e1c1bac2138fa864e19ea545721e705202504e884a96fe8551387b422c46099ff660c6711ab63ff834c1944dfef707ecce9c7f4508b247787e2cae38f43ac196b8699648a8cb5a302b93eb4b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef24ca636d70237615d00d5450673251ebe9781dd18cd0968f6115bf8a13fb2aff0268d017222ee12cbf907b30e7ad24a1ffd2925e01f2160a26fd4ecc71afe67298d937106ec9128a691db890f460a526318e415d22cfa0bdb50bee4171d6c7b8b497905fa2abc08a5cc54ffe8d4596fabd13ed867e4e86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181f9d46af42ae0d32a4a83ca9732b9b0365f7b7b7aa3c9ab1d433da6e116866f4fedc7ced95002592e18d54208c9ed0c56daeb2ba1f328b4f412a6270f156b082ed3c3477fd29f7bd24ae010184adebe0340047dc4091a4528304be27dbe68a530a6bfc32b122f8c3615cee451efeb04190d190474ef218;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h436fef65ffdb5ee2756d3747b71b7f15d40e7905741c8a8396dbb62c6b6e1225d22f40507a8e0e3c716544479f30061dd1de23eea86592c7ee46f671167f982f6059e7bf65167b82d2583f6cfe4825d9a239809e38e3dfcf5911b2570c101b354ac801334546ef2cedc7da29b04dc07550984a106ee3648f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab7c161de0a34d5f234fa71954799684156ad6740be6a9acfa356db129ae553160f481b30b33bd6f634c40838022602417e47250f5dcc23752ba9aea7e651ada53e20f2ceea8ca49786e1d1fe100bccce04e7bfc7e8d4dc8d678a6887c5a3fdfb57eb622b13bd18ccbefce9435153d32504baf75debd8b52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147e160b6fe54b33c93e41a497d8e27ea16aaad97569a27b1f667dbe49c400557d6f6e1213e290c48bc0b8eddbe1a822424ea70d4b534ff5c8f6cf971a878a64e8df89f450f49d0d72cfb2d84eb2290d20fe469d14d50c250f78cbfab004da7bcee08f37c8ce76700af906dcfb8822262d381da13f6a81004;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f54cf2f54386fd3643ff38634cac9994ed87a5d73313161dc28498d1cfc2dcb44cdd9788d556b4b82bb130f93296e7ad7e77364c74725e0b30e098f4b8d20aefbb9eaa30a376692650db7b6cd3790b40f382702e5800ac5b679dc5b1c67cdccfc9a2fa966c0e1fe1bb8d404f2d69223a0c28207494e16b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ea127eb8a4a36c040b372ad3af0d369fa17436082eebc719ec3aff0fcfe0d3151ba61158f266eb26e3186fa2c968dfeb1dfff228eb84a0715d35657239568ec52e48b23132b01a3aca1b030032767dc85762c6d4251f1177b2e46228da787a8202f550c7af85f16f64462b9fbb7d26ecbfdd7c02f1eae5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187f954671f661ecfe69db24cc0a504aae4c6f126cb0faaf8835f5e37bcfb0f9949d6071b7f4e7c84735cb90fefb7f42ce92914873be047bcbc025c9ed14cf435be84e3ae72c4ac16c238184907ad778d2a9f927376e68451f5b5f63f135b83b99d202e76ff1e4bb95f70863a03518ee47a87a4e7f965d47d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1050447769bcfbee12c608bcbca382d8383945edc1ced3b34d23194deb3e31d45f807809923e85848a9b46b9940f5470d77fb5fe91c135f98e727fe9ea65bb5bb95229fc54372ba2b6bd27d089db3a3043b82b390489d89a38f7dd12da4ae79961bb462b8da6ad7cf4cfd661aaa36c8f211f457321594ff70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf191dc2aa66064386e125e315bb14026b9c143c407af58bb8fa3bf2299fd579fc2db9f74404f9cbfd5e92df8446e2d4b344b03b0edebc7f5a12312812b589fff5ab77800f5ec507e9f4d65fd7df71cad70a6523b21082a5536de65e78b86a6b9b98b8d13700d63043ab8afc022c95b5490b0f779bb05722;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h983673fac3b63918258a37dacd8c14d147fac9777e67ee77953657885e83d6fafe61b60938b702162b551ab616c2cc3c5813eedd62a7f0b034ae7b87af93a1a1cf2a0f36612f4cfd8e7df12efeb18434e0e9eaa23df2b5903ee7fa718e4f10dabc85894a2bc5fb546417111d4e5c44e74969bc530a2b74de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he808ff0a6900bca3d002a1d1fd380e709e972b58a6d427e350f1fb3ecff1ae255ac888e385d161936b12df1c79b649849458643272a8b5bea90c63e1549d262110851fdc91945874efd5974b0c1a9106a8346a532d58d5031fbdabdd2726db1122f36cf687c49a8bfc8bd4a1b962fa2019d194272b0209f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2c004970fbd439713a293070362d66edb60bd3ca2011259786ba1cac0a6468eff02e78184cd3fc92af2a3981014b38bfa3d1c23975eacf6f40a6772490c626191eec943d27ab5d7728d69e69241a3df6f680814a45c6f5d9a6dfc04b27509ff7d161a47d21e21dfab8cce06e6f80fc69ba526cab55ea60e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32272fd0ce394d64ee4cfb207fc3bf285e1d4b8bf23534c1fc90f456353da8f6967d3a74ddacb24d68696f79df53f4a00afa951142c18d4e43cf273cef613a739a0d49fc3ac68d7cc7140912ca62d91eddf4cdc6dd0dc0e8d6e479fdec3ba0205786c35c09a154ba3886af1d4d9e28d705557eb0aad2db37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfdaa0ad091d29b583c49e519aef34c3f81336d3efd5f3a1000e9df61fa41ae5d596c95dff47b7c62b2c8fb1a27d221ddec151a2d91531d6526e2a63d0d2144c619e2f0ad7ca86fff0e83a5681880e7298c6cf1c27a2c9f67e4ea5016a059a1940307a47edee7765cf147b143bc050ababc2a6743a5b6a3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea440307fad43c8b21f3ad403ae1139ae8f9ba70170c2a690b0e0bc067ddcefe779f2b159c46d6b3db3926992c4cb507b02f7fd13872cdb28bffe9f0a8e3697ecc57b52642b86042fc2a4ecdb1a87c4c11774267ba059294494635543cf4b3be785cc7be9dfffaf66c43b0cafd7a46b2593ccc8b6cf3d4b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c1837d87847f9795516e5f0bcedb971e02171812394001fc44444fe89b7c59f00ff0599192869c35b8d5e5fd063e1fba6bc81d480e59aa370897e8ce19f19d8062de67ae5c384acc91c85b30c5a1f41b32d921ab8624b6535ef8a3b8494da5796ad1661b5ad427f3882223fa53937c36133bf3259247815;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8231a893e6d06eea27b987e5735a1a87053c299d50013fb97097f597b621a81364e58ba1e020da32ae17cb9e1db064f1cf20ad09df5271becea9e1452fb90328a3258d782e7250890cfd8e4e33de539a383d6494cfb90f051a69ca1f7251003dfaa55980e66ec31d2ea55eead4276febebb4dca0556f2ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1c2f618b5e2a0ff70433e1c3b69f679654c41093a7fd45d7047bedbcff29044c2383bb2eb62b2563809451971aa2a2763c22b0c47bff0e08308b0439934e5babf7f3bd91d2bfd487c3dce19efadc8070c34bc7a277117770f029d9f315299070dc970fe1eae2034f704f1d27759b5998916a4ea8839925e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee23d034b8b137f2777b11427669dea05ead2984f147e765a40e1ab794aa1e948d1917fb3ab0a477d26054fb9143a76c814fa8de808029f7e4461be1edaa398a8e6db17e3b3087667b973ea3aca18a7b07f7a04c166ff4e147a96aeaa73b3aaf44aa2844bca62b4264d84930b45113e062af8b2205129988;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2240236ca23d2104a50073976fbd57efc068a92817187b085097268cf7c983bbb7c228c1b86b5834003d32efba033a3ce755d0e31fd6931237132c7151d20bfe09f31e0bc5e82e9296cd0d687afb8b14d2faf52742f6f88021e291fc602fa4110da531b0274699415a649950d246ac0bd2e0baa8d914339;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a25f2b4edfa57ae4753f55ebfd654be18c311d093b5f67d86be93f4f451ac3d7219da16c94782a2d34b3223707f7c069ca4a19680af8201831f800b535e4da67d81dba1c57a07d392eaab9a7f8686677c7822fa780aaa838aa15822bf63c519ccb71cef9070828a8c5b6dd2df532cff09d4e108b1e9b2e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57779028439cf417b1cc1e8594c93eddcad33a3c713e65d7d5105a37168cb5cfe5a80ce95c17e340cca576a96d2b8db879c00779e543c80d0257675c34ac7a89a1ffd6e417e91414dbc7f4fcd3f0bc2e121bd79b24bbb500f2676267477cc161f361d6e3e415078e7f67d30a39c832cff53da80fc64e73a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46b324a5dfd89ebbf3b394600494b384c6956463f8f69e56b337c6d2eced84221744bc093f20b413d38926b26b8d0a5942fdeed0e7ab493e4f51bd81dd0badb2edbac01e56e6ef513689f0f552b431964bb200ae8cc838c99d872bdae1e9cda6f97ba8150a430277fdbabde3c4e68bc15d04e0a62b6a8c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c2f598fe9061ebae1794fcbc2b8547795511f57d8bcc80b2e42fbd3be880712ff31c064e025c34fa396d2082a144831c9d3918b93aa79941eeb10be0b926b0dbb06a644420cc3378df8a58c3e8f3dbbd6688489dd1d260f96874705888e5b64947cf639987e4481511e89bbe0fc79f8912585bfe2921aad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9890e0fcae19fa01e9f342dc683c6dd4de6f72884784401db65f2401af97522335b5ae9e4f796efdb1127ac8d45e9b41d11f5b70f9bfe776bab8bc0bc244df34bba7b921d76408730e093f12e228cc26616828f4eb9700294556979d330f19f6fc9e3d23d6d3abab85c5ea81b31b7dfd81507faf651fcc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d899459dc3994812ca24341dd226b910e07a69bb8d031636a92cf9010c9989884d2bb7528dad0106793f81a811b0761cd88b8b9a12abddf9ed29caa03eadda8be6b666051e0c1963b8910b0333073a918a16ed18585d98c8e674060789bcce9604fd2333291a324a7a4a340351f8749c7aa5d04ded2b1c69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192aff1deb880b4a45c78033045efa1dfb90d5705e39a61f5adfa85ecaad82f067ccc2ef8f90547b3f438f6facbe0405280b52a3f6360be838a047bb4db3701f396553a4f85183e4bcadfd8b95b34046be82031d3d34e74e93513a3323c05c4941afcdf41f27255ca90efd5f19b77311c99a8d54f3e1616b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e451b3738e73bc77d2c6711abdbe4c9a680c70740bcad9aef18c2d3b3604f7c364b8f1d70d089db5309008163ac76b9cd5050d023aefc193d79e718336d73ffcd41f96305861555f8fb17b0c933b4c50fab4506bfaec47d6e4fd308d2d760f4d7094e46da2b39413db7a543be8358293bd71c75238539d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c549b3ebce11c7e797c726944287ec4c28416d4b143bfbf98a873ec0e97ce11a4a63cdbd79a3e976d7d000856e8a2792c275be007a2662b53bbef19c647cfa229fadcb37741415134471c19e86cb2b72331809af27b09de5b1904c68ef501c1345ef15c846fef7b83de782779e4fc69bfc433ba9b578eb2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed42f5b51950faf3446158b9645a8617a1c35786b2f2a496e51a675cb3c8cfba280c9173284f62bc93543f79830d81e44f07487e32f83172f02e57981c55b9b33b094006f6f3cdc49e8c6fbda71036efa8b6efb709aa890b20efde92148c011bca74c26be9b3592f9201485f924204d07daba6cb4097ad3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bb6aec6c9f917c70ee95eeacb0f9f73acf262a4afc90d6097ee5b8ef93b87c9cb43ebe8bdb75bb0ea06bf9ad9cf0a6a71d7fde811426bc150a9c5e4068e5e64adde4dcf13d4c56129c04c307daea970265dec52063bbf02263812a3c1c238565879a4ee2a08ae18da3f2f8d398e97673ce2abd68bc6b89d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb550a7f51943e110218a82a7b08341ef8eababc95da7150050b4ea7fffe16a5f6b0cdf754bed7b1a26a31199de53abc4671ead0c3f9432662cde8a4fba853857a602db62fd6f0d90a746bf517942cade8bea644852f7240dc2b4fea5f3159993433fdcaa608ae63699c84cccf2460a5f43ebe7a17ac755c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha37491887d4aa8631903e83135c6e3f146f89d2d756e8ad48851dc1377dc69bab1e2bdeb130cf146ef1e96a901652d8627015c724cf6d4731e9f568cd56a3f1bd224ce9391bca676e2c3b3fb1a3d67439aaf00e046a3140e20e2835748d4c00dd8d8306632a9448ddc96cbe883a6429245843013ba55c87c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h290f0ae5cd26d4e17cb46a6e91f7a92373f68bfc183bdc26d8d4897a500bb9d982589dcd549ec6599aedeae368b8030867304d5008edaac828ea6d06f646cb98512e7fa1a5a606f8ac682421289929945749ab307ef7ec6b4cccf6e0e10db689ffe5e215f1b5959f24e3f36e69b7461ac836a81a2bde34cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181fa085705b4f45f26480f67841b52f3ca5d91cc3766f46ffb46ea57b8d4e9e3ec56b7cbd582b865c5b2844c91828ce5241818fc7cc712d53782e127d5a5334482c9328ad29a717a9c715a6f7b90ce22704f817b7d64e0fda14cecdb6cc1c5d4cd1d558ee14495e838553975376aba361f96b5f2ee83aa1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44c18a9f736ec617f6fd419e23e1f8048145a0a9d9c0ac14e7c277a35b827583ed2ef496f6174a92cdf4d9083e587504f6fc0dfbb22e596681cc43c3ff4913cc96c515f97fb93e795d008ca6445390b7206789125d56f2312f60e62e7e6a53c2b79b88a71fa390020f1b0b4c9d990d31921e8523a4b8f73e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h767686e8831e8d554aec7038642115265cbb85975f771ade1a00bd89c29a9d4bd2f46e9820b70f670d305724c4b6d57aec568c2ae469b5ba7ff39ca887abf1fb79fcfed4e298e7c71b6271959f28c090f0bff2eaccf074e38230f61444e6a6e3ae42463ff09ee53eebd5427de3cd76a4d04717d8be5b5ac2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf82fc9e030429fc6a83c1e514aec16a579b414a8e5ff6ecbaa393fb7a1ab28f546d3957bfae7c4a4511e46b0b7c09a732129ea0fead5a85e638ca4260ab578360186ae6d6c961ea169867c03fd5d7079e60bfd29d0d7139dfb8132d3f24a7ec525a473aaf99c54528f0121bc6574bf799eb7c1226cf3bf5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf392cceb28eb51e2c203b07dcdd002c3966933e86ad36915540ac0cd5edf8c0440e2f6dd4a6c8d248e988711a406157ff942a03dab3ac9945c62b176d0bed759f71ce9c2fd08096cf957c9f6d7d22f0270ba24beed4aa1587a8fe3d5be6b75f6c33c31976b6e804e375efec809eef615dc79129185d87421;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf33daf50821e12020e30cd11dfd3dd2a072c1a275f441bad9f3df1111772bf21134e1a699ff5850abe753815f9f7fbc70edab4be99ccc53800e487b5de67cce6d21b3f512f5e0b22759d1636db10c11950659b5497cb03fb253d7daba596f57d07d73192a73bd5b683014a4ad1cb893d9a65efa1dfa7a8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1370a3f5c2130b98dbc9a2532b42677eec048a3e3a20cef78bd9b4fbcca00840df4824bf335544964349e7bfcf9a7f3c9d1a57aed4012d109063b196af01c05e514dee74e99b73d8e058c508b806d906d2f3408a60726db238c8fddb963bc0c492219acd1035dd98ea6d3cb211ebd59f11113f58cd7a12de4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cbd32f2e295ff53501cddcf680d63328d585b5206979144cf64993fc7b7b976ec3d8b2eae7b7d2c82387dfb12b3543849e9513810271ed36d88ae76a704df66e4f32d4f00439d390a0bd95a8a9fded3c4a7c60a3fdedae913f97888fa4ce266fbcf859a9f3e72ce1fe359d948ef789ed3a6357c212a2fd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a8cec2dfbfee9ce57b23e854443f8e9f3d8b53d139c1c8a5181279d6bb51c4cad68ea2437177089fd37b5157149bb2e0533c4e85f91cf457178763c82563eb01994522a856a13ce6d2f86a692cf44212745982597ba5661ffa7b894659b43726bcc311f26eaab73d03fb219121f2a895db2f078763e8eda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c59a41ce4d37bf5183f33b668c0de271c59dae87b19a3c55e98d7c48d614f3baebb36855b6f510af4bc6b1d44e1f3f4cebec9ac45ce2d7d25b6018168d68b5795cdfa0eb0c066afcfaf903f27790b1b429f1f4368917281abb5775425b5588c249a84bd1d36ee9df98913932cfbc6f98e65f0951725d7fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8782c41433ecea9bb59d53bea59c1344e46f769b7dd9d9b0066cd7dd99ffcfb06c0cdab1884f48622d0cc091025971ab7d04ba9feac96361f4f31faa5da87027767cd71a88dc4ed1dfa54a4abe0cc4ef1efb5195b9dde8d0fbf37c85b9c2d4c67638db6b19c9456b840a8278a5aaeeb56cf574569c3ee755;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184c5b93a5a0dba6bf82a297a129fd8ddc8161b29869330e45caa085b1809061874d60a6d1a772682bb09ba57041c89c1f412d2fd99b9a7f6fc7e517d08e5634b259d0a1eec24f1e9a02bd764394af7f9646f823e99ea1e2419aafeab3cfd8e17c0d122c217f852e318495766269d0b249d59691726d832cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f26a4a13cdfd2d65ed7b944e20f0a00f15eb2b0ced497d1ef3a3d99398a30ea089804660646a9bccc7f3c3803256e0f0f01c679b75b86d351232889003eed10bca576397b39a024a75e6b54359ae665e88756fa16f46912d74c467004b80d76b33245fbb44423885b08b6e57bf0de2059c0debb29e15a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3408f01d3e8d6a4906855aeca5111d484b4754476e6791136748597a0069cf18e47cd28b57dc33d82d75c2abf09d2a329ee073194354d4754665155a1988eb0266e9e5929fcf79105591ff433c3ce629b2e72ec78d3088ea410d08744988a5cf13eb03df90a93f5eedc4d1619bba686efb7d8eabb743a04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6647d62d4aa1208d6cf06105666e623474c45012495e94e0a13a9912da2219021152c5a63a4b3979df48a41155f1e5f11837cc4757933d1e8df97b706dc6a1dff39990434f09646be27f75fa18aea995ab1c1a1d6ddc26b04da692f638bddc14b397368da365e470328e0239702f0de965126600433502b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc40bc480be2b955424c561ead9c9b7ccf40be2d688a1f157d0df72a8d4a398fcebb7d3cfdbc38cf995003f2d90fb2a7ae736beabfb1fbc21fdcf55f5470d4de8c28e62fcf70186c697aea279f521f374d7775af20e18b2de84dc8f5d40d772a39905aa9c1fad4e2551788df3fb09f47b785618ac4091a848;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128f867868f215233c15dc7283edb2fc1a07e169cf1be83abbcb62ef0fd333674f5a014572ced8f2ff6f85a3ac9e89957a8413ad1b4d572de47ac62a75b32d0e7cddf1015228034f56c551e691e58a8e437b474018f21f130103d1c89c59a0b321eed17836e445f3c1f9d86ed6c861930ca31a01b39fc26bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a539a5536362fd27a1e7b506eca4116472eb8edc3b2e0ff3232f1f23e2aa5a346c0089d12e18c2662e16dd80f84718e1146b5a84ba6216e9efb7dd67e1a3eeefa861452631e1daafbfc613e61615b86b88d0c4a02c76816c491156ede80fa722a2786e948bf64628ed6760e8f0be4711926f2f1a78930313;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70ae94b69602b2f4d6f21b260f028c9f336a6960b528e371bcdd2af1f991ab47f50819b000e9060b2dd0e8a11ddefb8f214bd1d5498820b742542bcbbb9624349864777959786f764be665144aea9d532b9289db60a707edea2911cc3cf7d4859241cc217af08c5f7af14175ef24dc4e1b5a9926db6af8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135e802d84cd4dea1db1303085f0e1a988050a84b9b8382ca40f28557c2970cc4aa25011430a05269a9b205f6841fceb7b3038ca8482196b5f167d6c60ce76b77a4799f3a9feb00de2a986276ad229eec529babc3c6badd32b950ac18ab6683157136d2f1f6becd15e4722030fc62b7572cd07b4ec92f905b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8a940936be9282f12b66e452187f4aecd4d5ec9a2fd164e7aee4b6a3e43dd220ed864560c9ae0539c9df0ea1190a3a4a23e9f3d441b4289ae7851def87d1835fdecf003cc09fdc634437e96916a52da95f02c44c2bae4a92543ecc62caf3adf8288431b7012140d9b8b7085ac939b21994dec47f6c54a8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5829f221ffeff572466801f0e8255c32adbc57a2e8891fc205726f3c15c80fad0f3eaf46bd13b680d14707a021f19b885656d55d385c6f6fc71615f24dd7b55f470f37d3a2ae61a4ff4f614b66dff6b322af4b97d808b7aa707b60aeed39b96bf4ba0dfc97e98355cc533ef52b096131e4a70f70b053b91d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1724f475bd9aa930acc9969edb7d9def82e15e26f6695a192ef0b997aa092153696ea896e441a564f13eee0d0a64c2f442889f93ef00320f0a7d4cdf4f5d18e5dec64f06e872070badd6ac07d1c7fbf2fd95a59df1e080a817d11c03812231c8956a5832caaecbe2d3b973d6fd4e0c2813fbce553fc2b59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cbcea19a7e60ff433ce08aa6fb9bc791e417c5dcc5669d22df1116d95a466c2238681fd283aef2c24c3fd1c484b01e54f93923f646e501452b2067485434376abdba90498471d122d7c877a9fcf3df25405a81489fd47f6c4920de8c0d072b92d386e6e29176342aa08ab2dd6188a35d47325f2473fe2ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1719a0a6884de03703f261b0251e17bb77b2c1ae9671f69f2cf239c2d6044e3cc15b7ba82820eb1cae7a0b09c6e8899d884508739e2a02aa54a3c7a44212bdfad725f23aa94178d6c951207923eeb86b72cfca1b98fe8a78f55d4080748d0c5aace2da59126b051a8ceafc2d780f7b7aee49de857d8d907d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbecf1c6177fe310f826327ea034963ca3a845ed21a56bacde1210e4aa1693c70121a3ea841b22a03fded736706b37575502e3a53865ba6d4fb9874f81347a8a488e86872c4491529009a45d99b0518ead225b60dc60bdd84d9af5e694cacbadc28f7c177c062afd5f0263c16c615933205fb4cab5a03436;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f96a8435d564ee4b9a830f2ae9359653b1d0613ed90a0e857fe4cdcdf9eb48998c22a6ecc42c6f1b75fe063c2279c59380c38c8ff8e5d6a82c67cdd7f0cc4b25961b5962af984bee1ea348e7c13885e7bf4f6203f3e169a87a1e47e2fea65ca45ebdaac45545bf1f62528554265d36b6199cbc82abeeb131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had73728b109e085187d78ecc44980d873232038117c41e88561784341d1a6e874b2477737b5049bcf31d76e7da323ba3c07c924fad6075adb96f6011d9a755999642af06e8e9c07fe2702847db5a683529c526293193ff1dca895d9d801432caad8e7d20f96c3e3ed7fb5cf8cd4a2aa5599515eee112e7e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c4294413af59a001a9bbdc2ca172a53d8fcaff59bde5c9a40dd484a450b9751abcbe298d264f799874df9720f20679828d151f7db20fab6cb38492a9bfb900b4b0b06144aa49cdc9579dff910b32529ab4d82fae4631e22b3f1b02d226411ffd47b75bcef80930e3683cd43c422d8e2ee708c30ca1a8ac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7c1e61d39812c4c665c10784f877033ef61b46834b0d1b279bad7e9d882d880aa12536bdd3ea593629f068017c82a4b95fd1c8bf076fd7fbb3e88fd387f47eea33f386d21933dd1fe975faa87ae3bfd5579f3bac24194ae5fe4bd509a4fb82ae54a0e9f2aa88bc992e9f9073ad3923941f1f346a661f174;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf54b580beb3bbf33b284586808eb845a79fa665fac5fd661be89a01afcc5444e92c8af5a293573ac04caf20952693e4055de8fc5620bc6fff9a9eac95114724b47d5b329dcca360b4e4a41262f0ef1a9b58c7e8d4703358bac0d03312a44e212a2f71817faabd1ad3c2c37a537ee351c1803d5d9e1de8b4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36f017fdb2ce615d289a4c06d9efa5d5b5df6dbeeb60c3b62610bad64c0f5c2d6d510da3d0ebb8f67e046fd6623c34dfd6c1037559457c6c929a3f12a32de7d31dd88370a558bc8d956cc05570401e98dbaffc8f46df45050fa18bb6b6c819b3fb75361d804bf37a64b639267fc23e7e60d7490265c3cdbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186a7436276dc1eed6d98e98cedb9bd40e7a48f83b3a770757cef0cf2f2ce8b2de516a164bd7cc7e59f4a2a2f6ec44912e4dc7c9257373717ce6cb221c85f2ec23ccbc9e7645d6d86c3a67f008a44bada6ccfe82e9393ba28aeada3ad0e4df9ef481ef7e7d6f26d8e290578646b111fc804c2d46d750031aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e906b26d6edbd8a9ed2d3e1c090fbf20d79cfac0348c9015cbda184504d412df0cc8624fdfabb9d1ba1a586c0c3b4f15a903ed33e57e1a9fed24248c92ba1fd63703a8743ce6287e01a0c49f5693e22e261cb836f2cec57256b554533adebcc422c2d636bf3407f083f1eb015a2e8fe2cf0e388f8e697b40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h445314752a2903ed99bcace49c1b6969e550486268814953104c662367d46a038e6f2ee3c71d1159fdb44c41588d17fea224c03c2216430eb8d9cef2bc98623a6368859a94be98a71326b0039cfa6d895c356c30f2b320ccc355eab2b5b6813cd0af0db9e413020c046ac97fc3ec5e8a13a1df53a57062f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ab4f7da6a60fdf3a3c9915be4bfe776dd3cfcc0e48c2d5f2fcce574807ea84c438dc3637b2e97f2ff8f6c07f413004cd21aa5bc8e5d3e0a83b0f3809bf9af5db51c929a517c7ad4a968ad2afdbca97c73188cc260f8f4897230f3a6c8db0c94072393e68b6deed8f3f8add49a2def627fc29c7f9f478c31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45666ffcc05335f4513fb148dabe5fc543124816080072cdb0a8d7e563201079779f63a1245cf36ed947d73fe24f644fdad3575807044da6fad973fea91452d13f22ebd5e4100c1c997f532ba3da821594d0fdb65110855fc4e7ce60630491e8ec97215e267f8278a3685dd2621a5c2bc0e8af896c1af2f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133b9b9ed2854045a8427083d4702e8a9b1fbeb678f081df417f3318f1bafc0157a42bc3041e22b5442785aa23c50be0516a83aad56dd449eaa6c01e98110831bc5254f2f98b3e6127c55e01f1b2cda629dfb24a2a7a7058849d1b209ba628b394df0dd2200a5ad121f76902b8cc17913ccdb283c3b0822f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42592664cfe6ff292cbf9421ae2d23bef2492e2f20a3e7f4c8c7987c78e603d396f87ff420ed0870ae1873a9c0ebe54e47668612920812033f9a310e92065518ebc74b21c7866db37b7683d11b97e7e41d4b6642d8c9e128cba408dcea9b21b69bfa9c491bcb26fe7226b4fa4b07722a72434950a1479f53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10460131c23fea085731bde1dc7a7ff52fbd3f5b25085dd24a25a4817a016fd69aac667ba3732914c6b04e96c65e161d6e4dd731e8a16ba35b7a7b5dedfbe73e41de415eed16e278605e26b251219716164c19f42fbbbc89ae5c0516704ae5c9d1a6d638499334c48a9fe37558304943075093a6917b9796b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8c0642cd469fa9a4cb767e5f7449cb2c9a7464b8e7530bc0bb0d5adef2f5d26599fb2f10b7aeac4f4a7d38d35d47e8dab587213029ad09fa39431215db8fedb64f9530ab67cbdceca09235e9bf057d21dd9b1e624f952d811e85d7e67308bba05b3207e63ef4a0fc43ba58b54afdd1e1f6a59061823fa93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h621d6e0af2c24335fc4e69c5e057345d97c43df9853b3c1b5ce77f1d16eeeb402ca35b4aaab826200401002782755b00a94a60e573b611531d4c6e3724d729d7dcc69162729377c7775480b89600c7df121190aba8683f7c3707b15f220d5e9264edbbd01b111544a980afd00020e6623ecfa8823b95b1c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc290ae71f0545135305b0693a98432b207c787e7d0431eee70b03c34f0e7a123b27bab9103329942f4a13ade76c79efa35ed0a5e3e0efec92faec302009d1fd6c894f3d77c8b075f004167360e857cb6c256d3536f88eaf60b31c20a80ff2ce8ef9c14c43eae6905ec62f73cdd1f71bdb586341e2a97a9a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf62ac16b468a394b7ca989819d1315877e652d2632d86923fa997307326a4613c8738394f00cd977b95a8ddb4af5ea6ca058c84569d82e39dc56a357b56ce08ec339bd932cb8007668156478bedb87328ff1903f34dadf0d82ea7d556d5cf53f0a9804313814cb404ec37f95eb4ba2407f45a39eef4de1fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16df8c135f12fb698d3016949fa0345bd3f1ac3021e8e7bc8c6e7bf36186a68c2d548b3d2dee1d1faf2106325d08911f2dbb10663f51bb4b09321b1a60f16dab4eeb5049d7d85b00951ecc8d1c66864e23b0ba693b4222d1d13daf4ceb006eb809862aa261d70113b62c4f1d976b465f3b3fd3820043d5bfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197958ffe6acd3ef2b5866ba2914bb6841609e9c01a8e442052e9f4d6c69d281b543a97dff99e928aea7147b4c063c08a79db23541125313c496e8968fda64e8000b26748b54cf26fb05e543003dcc7db3215465d9aa5a8e7afaeb95f18cfa6e324ae6b70ecc2c48a9f858da0cd00252753771c102060bbc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd995b3f0d8256d5b1b7fdf5146aa4de27ab4b7d3fd5efa81d45684a9bea47201434e09d4c6f5cd3e507dbd8e2945a9490783e121790fde494aef415f1f003cd587e330122c80ee323ad0948c824c78e8d25a671e6965ada9e38a94c78dd41138b86d27a5549e384fbd51cad24d0b1ffe5d26367739a9a32c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha03c2b07a64f96a5899eb0b3fc2e4bd7eea13ef2427185b2ff478ec9fff6ac68e1b072d870403d7775b52ac7ee83785c4fa8e43cb505bb211b1c223807823391fa638f0225ae95a3e254a75155367e00bd0aab99e9c2b0a09ddce9ebaeec1ecb9d70f4d4b8933800cb5200f78ae689460e3e2d7d1370b985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166ab4cf3fd607d5b8ff9ff0cd04acfce3a403f95f6236ee349f90597459c1009d8900bff4f43e9de986bfdd7b554def994f25b5bada423a3e4a4271a0c64d40401b30e7349f0fb5344f718cacd8fed3e85607063d154b1db1e748b2fe6402155aeaa989398bb85d17dcdee4d4ceabf1351001b2d37e41b5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hddcae98b950a0f8e6d29326a07e453a40cb1db562be102ac68b8af29c6eb07253dd482ff770cca555eb2e4a8bce2b48c241e68ae57ce186442e2e3e3991fb247f83511ae4d8ebeb3fbb1eb125e84ef82eb9fb791b34cca91d19bbde33b278756fc001473f5d160f673b0eeb41f69a5323aea3f087793cdbc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf303800924ceca96e13b6c501637f0e19df1bd179844ebf787e754b4ce6282c78640e2b089ff2f4e2b94507f23ad343e3eeb223444f265b43f80c0262d7f0f86e415f9d3931a5cc030f8a903dc38ca251a8286ee1933e5bf369748ee552dcf4710073e8ab1e399dca1e34fc9bf7d4cc47167d64fc51dba0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b7dd5d6fae011ab2c32c49acb0a9d7f0e14b7f5490048f0d7cfd96acb5393370423c64a9e0f54ede1f0712091828054c4bbafab8f2ade52b5560f6849b44b9a74d493fb260d2adf2c22956a8941599fe72fdb805cc14348fa01dc9a4583f23eebcd90daae4f9aa7de2061425013645f406547eae49f34bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89217555e7b227111fea9b78d45ee020851e054296b5df789566a60098b42df3cb35f27c38543fb9e73d588f84cfac0c85891ffea4d709bdae70aafa01650798e2913a8cea3250b856e66ada876f63a23aadf24b91a1d497e78fff8c7b52fa3112aa65a0204916244a20311c3a20c2f156e4525e117ed10e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9aaab54ae975c6195dd97b0d1207270f61e18c0dcf669de64d629437200e98d02fff47b9ca1d002b63c94bf9f6d3ec848da7e4b7ff3ebcc8eb1ba0b6dd2b86f411dd2aa9c654ad847befcb23e0847a9fe56c7d6b1cf76c04bcfe7087e2315664899da977224a6a4ee70cee84d5cb9eced34a049693d2ef3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c73b10328e8de776595f23d689498313ffe856924d46fd993966edd659a864845a092b482d7c1d1d5638512ccfb7f69951fda7dd6acbf370e76f9d3626b849e20b092b0937c31a73b5671baba00de5b13016b204cb6b0d3a7c1e9cac11a780ac4a8495e2e5030e2a1ccdb7a9354f3834a975a9a19c50d81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e26db2b6666548d046eb384de0612d4ed400f2b26a8ea568dfb9cb47ea02c03c86ff1e1984368354d0d228510f7f23d2c5188fe3155311c4fa9e69a4eb0765eb78d7f81562ad9d168142c04f2d00a143d1182dc1deabf8b50fbab7004ad34e617f301b2f4c4afa7d88282ad00486361c4fef43d566557cb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116a1d464bbcc32d81f76cdfa284b3778745665f6991e822b3ba880e9109fd7cef3c29844b6d44197ae21d856d39350f95e36c9f65c82e9784b02c40ef4257e06e38fad60ed91ce1d3fc7d615542337b47088b7eeb87c582c8102b398d0c6f5dcab879b0067f2a32ebe1fabe9091794ab8373ac8865eef5aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160d302e77c12284112a613070b7b77eb132b29de109504f9457ddebe2fc84914eca192f76030483df51b4a0fd46e76218bcc9289733ccbdb58019968cfbf0418a36bbcf6e4664f1a3078b4ef7528f8c682d097eb99e583d8fe9b90e00910309ce52c97f45c8d59b3a2081901a12264797249bc3f698f6540;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12536c6b33d20788b386b6e6d6f6a932af76196f0eaf641f1c2e6f8b07ca1ddbd33329dbbe9d36d99c21ebf816c9b5d6149deb3ee7b24ec3f495b9437b21ac3f4929cc567b05a84d39d648b2d8327402aaea023c31c547a5c3b8dfd85a750b02766b0708f4ec7d5b8b592eef9c89c5f44c944ccb5411e1236;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44e3b254e1269cd8be415e8b92e78e1ffc6d1ec5aa1bc5f48a4d0f2de238af4831618bf514d59e67813fc702400c6be597e3ecc4ffc58fdac30ea5b06fa33a7cc20081da98b619b7d989005e847f27946b4ac29a236e56ac7a1e93224836004c29ca30892e4f59bb092e5f7e3e002f5a3ebdddfe5ea1e393;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h960228df5126cde3dc24b19bc608be935ad3c734248de7e92c3a5e9cf2916135986862d1ed67546c640b92bf1ea2e5754b58f39b3d12c8cb5e1c2eebedb7c1a7c1f79d6ad0675107ac805c4eb557da7a226229a1b80d708913785cac09998968eccc123a3d65fb393a564ba860d990231fd142d6294200f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b2526c2e9c63f88cbef1d74b7e1d7622c9117e1ea2896ac5e832a82f34581ee023b1502d3b7e67ade106d08de36f5ff069d7f49723c4a0269693c516040b3497f0843c9e1394101eba6dc2fc78404089dff33f6b8def2f900768cc926e0db90d3541c4696ae9211d950c6a7267a14cf4969cc37ea2f79e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e7245a5020b466c47b29a4cd647995a193897d3f507825acc4bf4d86296f376a87ac003b206fa3e64084a3317cac817b56c4f39ca428f4187d4ca0d4814bcf4c2c8e640992e2852a0d390942c9b80da4ae79a9df3b625376ca7e8b306519f6c79d7c2c26a2bfe85d43692c421fc18899c79ae9e9ac93d72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11585b10319c38e9c138082ff54e1dc2b53071e51c46a70c50056752df631fe9313286beeb31d0c7f1c5b7e1c360ef1c14db8a43d12be8ff069a841a41f61fb0ddd7aae43ea9328ae02aa3c4f2758f229395708d7bc2893f77eee32a9e1a4867a7acbdb554d091a0132a4d02d689ed6fc7695deda5e98a94a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h858de82cc4c0d018c048c26a3022bbd808dd7efae1b286672897d60161d77baf477e39d0bfd7a2113965259a4c65290aa9f602b32f35ae807fcce2910372cae6c05caa36e55fe177f59ea7d4b574420b9abe6ae53f545443d59a09985050f18088f69705a50d26128459fcdc233632573a1f570174bae780;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf0a47a0cf2d09209873e0fb47d72ac76aad066480e01abda1b284057c099a8bab97369824b14844b94b6c9c11b225791d625eef75aa78e6c04a921b60a3ada03a21449f37cdceb69e0510c6cb7841d33c7206fe35c3d0ccf439a073d5fdf04c571d4e99df110c5c14f67c42d0a9b84698045bde2a10a051;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab3417cd57b15c2c49fbaf5bf0744b17471999567c3b027cc53fd4a9ed5d34b1578f6fa4eebea6044316760978e8ce601a70e48c61ebce27b1e66a6bcff6a980eef88b97463412a6da840ce872939b9c087886f3db9eac74f01397bbfa970385ec46ebb22ff5cd694020857d04f67f9aa8c4c78b40cd2211;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e53888b5b185e267a6f9a6c60803967455b8552db50739609556a3170e8b0640d7a12857be398bcb0e5d8f904764c7cde8b23f4d6b7cb6c54826a649db5fc0696faa1e5b3f38cf1181c8a4a23439fc3ddd51546455a237df87bdbfee827c2805bfdf74f6149a487b7a79004b7314d06c9d86b5929c9ddba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15055e80cd2e8086ac11678acb199369b3449e8833df291205cdf5c0710cdc2be83e2021f9e61d93a141d67c703e11193c3a0ca2da8d3d9ffb50583b8b83f61662f5b1093d323203d67720f83d2839d642ea17eae463be1da5a9ba0e62f2282b1ae6b4d386c186dfb3369c771fcc29973ef5bc773b8c74aba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h705b1be28849ca1fc96acd53425fdfeaf327ee641fe58fb8eae86c5068dcb42ac4efb8a63aba139e12cd6b77753b3f0ede92f6d1c563b5063a9e2849f2e4d3e425c0b9fdc11b7f2c9877bd3249cbe0e09732d858671029f768eee394e12fda22d3db41b5e09bb7d2d564e7ed8436ccff0d1341edf9767279;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a2941dca2ab1d9f421c8ce73525f502c23499b54ed0d6169cf40e3d4a95462118e17802ddd519d3abe25ec0ad7252ff87e0aac43afb3fb399e38d964a344207fe68fc2339e10cfb4b2338c0b7d6c50c8c5a27a993e144108e03c3d344eef56ab17b16fa2074804f24191fae5f0cf17cf73ff69d9c362b63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8dccdb37b78a2ae89863b894eaabc73328c013621786e0053afc666fded89bfd6af3eb48e36e293f20f20009eab6bb4344f20079c3e9c6b6df221b1fafcc008ca04dd74a43f12f7bb6ebfe3b19fa7795d25b56c04baf2c9c340f340fd021eac915839d36c7458316a2e47d80e444b2926f3e5de3d7a448ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha14412954a0691897bc57fe2114b23d9c87c45f7f8fc7ab918eddfa363e4ab96e9151a8277f4154f779ad01dbba742bdb2493e1703b21e02a552d5924cfa4eb1f69fcf2cd96d7868bd97fbbb3ecf119e04ad5f0de1da620bc4fff767f8e3a0d1f3d9a6b1e5b30e66cd710f8bf0cd259c12a3c262b71d7850;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2e2991aceffdb90115b1e39e9955a9e1fdc0603ea99973fe449844b6ac8d873108b377e3c3c739459db13fe85355e867b89f7901cefaa2a2b55e28391e568f0fb0ac53123ac8aa2254ebc7967acca0d8918a01dbe7215c2f3a811024d3f8087d03debfa1ccefa5197d045c2c76a2f6aa77645713c02aea2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162a1860343b1d409c990d07527ab8562013b716cc179d758814a51fccaf834694e7d85bb3fd7a08346794449b35293bdcf8e3f3f5f52ec062c7dd664ca8a052d6090ef098c1a251d73855f0c0c61699b60a39582e685ba1a92532abab14379343ab35b04fdb6449d1d8e4e1e0acf837fe6365dc4ce0326d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98b9f1af940db13c2dadfd9a0b217847af84dfb3fcc33a04a8b27fd271a213ee5b05a4dfc8688510167d548ec714a0fb8caedb0c1451636ef207829ebe539d66989e1168cf23bb0f44f44b1713fc665871735a289831e54766236105cd7a294720abb93a04a001244dc58b1c8fa2d929e101b859870a71c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1230fc08896ac5a6e952b7c88ee2b59b160d62bc9d6b86e108c6d85a4ab5522760aa5aae5f122557ed3abe02ab9fb70cb8a34057eac7f1c550916f2e9c27441c0fd7c309fab4e149bd6ef716b1598bcb723d24f7d498c29f24d1ae7a4d892e384a2ceece7952cf15a6310a9f73bc7487094978366d39dcade;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b6f656c493d9e535b0d03367a735e484118c7bab3fefd93889503f206d898aa30087138075cbfbbfbf5beb54062b8a5c22453e610a7ea948c0c05580fe31996519ca72c036f970b97357fc74d4c0b92dd96194c79474e84d059087b811a14ec0db55c9231685f8eaae95c9d68f9d9f5b4863106741fc852;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc89b8f9ac28def470ccbb2d901ba18effdbce61e86229a415744951a69307d727f230eff306f798040d1c34b7aa42c4fb54f44ff81523fd6432b5e9eecd5af9cdbeb6bccda493d60f0bf462e5182b3486cc7b6e2124ff73892550f8c2d135f0046dab44e90e35ba89e1d4f3de114f201804b87fb357737c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a9ddacecee5b42373e482f500de2ab3972191e397f873362dd8f718200e0866a56a3379a56c0d25680d01696f1c624677287efc80324354761fa8cb696c08602ef83ba0493531363910768ed3c7c199895fe46f05cf346d0fff2e2cf529e350ad9c43c1f73affd8950d9b714f2078fed9a0d823f3f9bcc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120f4a60d0a68048c5f3cc0ed48b938d778a6c338f2b19f286ac21808739a5229a6e8d52cba0d79b1c3b96f149c81968969d98d9ac88f4a35263243a378fb33361999ee8c4483ea8b19e01fbe258bc3e037a7540a7bcd0a291218ef6c686dd75cddadbfb563008f3425356bf5d0a9a9705ab11cef2054caf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b1e59d3090caa704b3be0ce0e3e260427aa312742986405f3fb47987df872ce1fc2921e5e8d285e88b17c65190a9a906049072a5abff787822abcd2d489f8421a974b3f0662cd2ed31a5aa9cefb3badd6ed26095a59947e22874fd196a4e885b409764f2107aa8c045db7dff3f2e6e27f00061d1a766466;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1854ada2109ef9d444b0ebf1383516c7b77bc72e8a0455e00a2b22744ea7ab0435c8f123e9f6006c4263c8f7220e3b83695890dd4752fdf90f92b6691befdd8f0d6ab76a0dc9ae1d79f0214a3acbdfa11d8482dfcf06b672aeab41e3de6440951c9213993c9f49d007cce9c631e75d386d7a9a87768753c98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7fc9587904fa922170981228920b64bce43be87d3790572252c4406aca9b5d5267e130cf1882ee7ed7e99c884a814b4890a0166d95b24994a1cd4e7785b93a223401ee95e497e5226757b553c0af34e4c8b067362780bcd6f79ef2671829b412ecf365232f8cc2cff3f04f215bf0f48791e22e8883be02f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170df6b6332f4bd7f3245599f43fdacdb60b8adcd8245c37f97d92c18e022303282e9b071a9b4e53c7db5ceee4db39faebe4339ad3e6c075b2e3a676c3b31e787a7821042f058b25abba7479f2b3d1753306d934a2cb63a463e7f2a5bfd320f7f6ea5c8a0650b9e9905d47ef5309026c176eff9bc8689763c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bd40590384b1f2edf890534f7640acd7dee4360e963471502240fdd38f49b261297ddcc988a408096269c6cb12d9c598b9bc2e4b825d08e22547a5282807efb78102bdcc6720a69d869d09131139f71f229ec0a5209d13ce81ee9c622e5fbc7dcdacc4605b7593a1886a15141ebf648312548abc4ecb292;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e5f50091893bc58ab6c44b45eb5dbcccf5b10a3e282b244e433eb392749f702aef429d1722d167167c563398503d2cff9b7116d8c91c8954edb82ca0742feff3c5b7f1a1b7792f3bf756d1dcadfac0e31d60c5b9f2a78d9974ba5f47fc9f8eb1b046c663dc15c966883bc1b196def38340fff2901944820;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc51e87c3871f79102b3d53c1e8e32272696dac3bd1cb9c9772ac3c34bff882750af0708616b01f1b775eaa60b53ddcf7eb379623f8b60733fe76410614fe44d69bb3e92a8f11c844de84ad49e87009cc88d32e785f40d7bff1ee35666ce102f53e47494e04518a800f149f8f6794f868111168988d1b431;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h532cdaa38e82fbf0981fa2dbb38cf562f4c3e40e5630e6d77a353ab9e42be1a441f05da965601ee931152e39090c5d8687bfc7427dfefa28624dbe7c56250b47664eab5a5db2c9709fcb540dcb4a0463a9d0c4d806fbff3b1baad77a08afd7208bb393bd069b0386225d853727612cf75b81a5647b47165d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7b91412d0c37fa17f1e664802c36b5a1fa8950271b14648b44aea92aa27127297c16d871501e7eee3c54edc9a11e9e3b180810d40dd21fcfd72d6a8f230dcafdeab273b18ea6bde1e2e12c104ec6b1516d1e19b5faaef520b066f33597c57c2ad120b9bcb24af72eb01c29b0a4c9d2222cb79e8ce13c8dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he625495a963d6c5670d564a9f635977673cf30097b2a1ae0a8d70bd0eee017e676d8c92db7052c1ca7d0faa783e51c2fbb5b7b5eb61892be7f41580357df073820b326d6d4f7705b3b3ee709e253ac29e2095bc100a99b7d1e2609916b71846838b65277cde699e20181b84e53296ef32f34d8996b85c5f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194ea98085126d6d8d3a7bf0af694cbd927f77da0ac48c078a330bf17075adcbf3eebe094e3fe6d6e7581ff6551cea7e3f7fa7b48a8cf1a88e5f7c710a21f0ac3f9b2c6c6bb597ec09b0988d4f9e1f35bc6f06ac1a2e1206007ba9d770e177787bd805a32ad3830ae3c12e046ac91febcf9ff32e14a6f2858;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h843115bdc615edd3b84ec8b5b8004a426965736538d0e3b1d706552517b9922472f611773fa776b88a1091f3d9271e3fa089b679c8a1dbfc40243ccf95077fb46a59ca2c37176151f022bf28a3fa0c935b7a407ecc5c46669b82fa5c3949fd54373fbf5e6b3e5be46f075ae3acd35578a1b46174d408a051;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f35da1c7c4d9b020160e7ee2f52edba72e2ad8a67ee2118cb89b49dd6514ba05ad1965b099d82fdf04170c5e1a2708ba7eb351afe9fd09e526a9685d007451e4438871cf77331aefc50c7c02d049f9aaf226ca42e9d3ce0c18ba9f07730cd4d8a1dc3bc95b534cee40d135bb3f5b756dce08bbcce7f0949a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fa13043479b0156fabea032b4183d7782c30f75ef2863c06e8756643b050ed0fff3574f0d7393c39f1e1324b96b699334f584e028c93ecfecf0d14da71cbafcdeacde702acd1d8f212b3f1fcdde0164866dfdf840d0d13ca6939e1ee7bd82ecddff2a3ca948c0de15af284dacb3dd468c63d40ef7f330d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h731ec1f7b5f0db85365860185c4c676727b5adce342de9149004b4a476204fc7f5154aaeb0ce50dc74d4b6cf5d5eedc1db3d1d907748c93b7c9eeb53e93ffc0838784c1e09f5cda1b7fed34bdb27061ab5f0a9bc7984d8a8e8ba9c2b6e2c20c9efc84eea66f9bbbc8d7bdc8175f33d85d1a2dba21185995d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e63747298537d017f8ceca7088537ff7af6c64d85056a5d5a66037b034a8525f950d12542993f22b7159a9b8d268645c851d190be05958dd359f312fd50df102f5cd9e7dc4ed23e1a2b055820420c9c1522d9fd42816e033c4d8061ac770e7d55488cb21f9c7047202417249f062856b0e65e74ffa2ebd15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13112fdb5347b52547274413053305856a87a89c128fcd1cf12bd29e994ce55b6f416119ac583f2c6104c69fb4bdbcc1a6f4580acbef483c01036a56dc2fcc839182054b63b59879fdbd4cae7a6c3a01e6acf884e53e6276bbfb85d696f9a664af2b16727bfd3a83b903e847f9246f4ffcb4f0b5eee686607;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3bf1d42b4dc24d3fc7e3e494542b96929ac6b8acaf06a429b041c6ad0b183000d429adcb7c7b629ab9776060ba56a3df250ea75b2554d2dd56c1fd737fe1b5637da755a89660f1b058986bfa122a1b9452666b4ee8fd06baa518067377c6acfa0f3ec97affc0d6cb1096a5eeee63cb3d39df2394dd8c4c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h500b46cf89fe5bc30bc0a1b56747c69b3b0b09e28727c1a041eda5021f6d329b850423d159c410298eacb43934aa94a912c56d24cbd1104d3280f00e5c4a4df700d7e95a4a4736bc1fc3e99975ac80d1dbce32d2795c2179de2e77597aa12ab76e7ca2f22fb0d9761a6db44699e6cb6b3ae4a511e3937dff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114576bd192fa42b3d61553653846cf8ac7303e3f9d033977b17688dbb69a6f5b49d2f8eb86192b546fb6cc29fc643b2fa59ddb645cbf6882f520ba7752113d344b78dd18ced89b04e80fc86bb71952c5a94e182bbbda2b4fafcb766e7fecf12aa870cc0c55d90847fd942dd2764dc3938500428cd0804944;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd17c175cc39c067ff42237fa2dacebc24d96097d24b6f0e4d91c4b6da3c35b81b57b5fe1fa8c4b99d27f4835b0520cca0a697d892770957ea14fb67e63c3ecbb7d6627810f899a6659f397d434890756d7875ae052ac0e50ee486b554f58e1dbcb00debe3894c1c8d0cd8ac056bf1aedd2642d998e1c5cd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c30e25ff3f18654593c9f19b7bdce7e1c767b8648fcc743dfe71f2577567b38f0d4cf2969f07406c3242a30b64e9fa6e9ff3303bf524c34ac877e9fc907cd5fb736b5eafbd1b23224404e39d48e0ab56ed6128617e6b45a68577070b70f37591880954e588e6d6bbea88a1d0c8397ce5a884a270ad4c40a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51feebf74aa739ba131fad718f375f846138e2ba65b7dde34fca29cad172145f39dfb7f2b60c1cac55c49835969a0aab87a254b9a6f7bfa049f77f4ff18f190e56c700d73ba704a541a4b6e5b3a7bb829c42272e6bb50840f72df435a87cbf2600222f8ec20e9ee23b179c5933004f51793618fb9bbb7d44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7890f4ac9087fee836eacb1c31e9bcfc14ccbcd61dcc488a4fcbfe5f40c9489411d56259c248cb7186c0f378d2aee62a17a6f4f0ba4efd59034629bc6b5a56f67d2d64d937ac3465bcc7d7a016a625ce0ac7311019b878acd2ea62029c2c03ac3b81f3ad38864a6eabde068fa0bbac75e0bff8968031f6c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb4440e5cfa1108bd4ae89837f596d19164a60c394e9456bce44b8cf24a0bce784542fd3f079a3a047ae7704f91fe6e6bd06c1f7ed23185bc66233af21252e376dfc5a777386fbed61a5623aa9f5507e4fe8bd8ad8062e6285cb554dc896ae9813d2bc37e1243a4e2bb851923b3fec047869d4e09b9af1e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144bdebd1057bdffef0955bcf885e9ae57aa067f0ee6362fdabdc3c62efb0597e91960159cc881b7dc9ee83872e2099c9bd1eb77739567c845b0f912e9910663e49c59625b5a299b248de34e835165eb7c4e49ac1738b2f8ebe8bd233bc8db49e6ac9421f24de604d40d64312869de0107f4f5a485d3a8e0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f557e84e573f1d9bf3dfda8ed068ee7225b7c9b81c87e55e8d192914caa425e67d715cbcc35975fb45e35f6b9c8e8139927a175cbaa4c3062f9e8e95c434eaafee5cf30899900d0e626f3e4442dde7d4053a51641b54f00d320380139e2440580869d420389424c906d344a310e693c69a36c1c44f84efd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9acd6819002b25fc82aacea1504bc8fae87690fdf27b75e38e887911657c178ad99ee216b99d06a742bf51e1f7a2fbe58c1af544406c8cd2d7fd50cf8071ef3d57bbb3557bfa53ad574b684ebf4e2631ec8cbd0879c6165ab3a49b7eeca93b822a05099d59c5672badc51c2c99f95ff6035be41b63f216e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0f3dbe6ac3d51bf697962682605cd7b944ad6dc75021923d48b2507828b6d53d891d36d1b3afd0aceaa7df3a4bcf722c6e862a938d58553e13a3bbadfb3c412b4ba32cc4159d678f7703a55c06a0c6582d3139ba60398fac75bce3f5c71aeaf240f1bb4604a32eebfde6842144a735f3ebb0277487461b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc287ce2ac71a691a9c00ede73b6ddd686789aa8c167036ab4539ea2e5554124849777dec2bb6ebe82fe169b4926118faf618a5ccbfa086f1df85bd83fc01b3bad900341e4578548b308f274d54c45c5c837d7af463f3698aa02ecf3d8b3b6acb696f50ffb76a849c5e55adbab2a79a6c9895e12d44c99b0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16fbf4c25db902f36d44557fec1f169d251b155b349a0ed9fccbe2b5cfc40fdfa678f75fb337e138d0884f587308fa6fb6cde6688566c0d45bbdbf0e139e3426705e79ffec3d67123956559b9010960f831c14e9e052ebc3f959003d966fed5aee1f4ba2747d4328d21048d97efe1c01f7317c54f1d2ceb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181a3d8219795d4cc197cd711bd4734664248d3c866f5ec2689b544514b1a4dc6195b655a2ad0763653404c713f85b5ba13322215a6e88619668e5dc0ba60712cea70fcf3b299f8aa903af943c73815af30c0ccfad06061838d506e75c0d64c985d113cbec974543c96ce932bc72873f1e33fcd185b5e7709;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1387856fab2fe074811e1ccef46b85eec4265232866f1185c8ca0ff131a0d22f1031b919edcaa2f9f75208e104a3fd9f7d0a904ede57ce6c7b11ef0da38472b73c850f100f4b57ef39c0ee902a809295d60bab38dee5f913033cb729ddc58f81a233c0d35e9006c85a15bade746ed867ab23a649da9a6cffe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4cdfbc7faa675e8d23469a3e47388cedaaa20e65f78bc9ecb1ae4710d0c9b5a1ac47ba5d9c547ff3c3aa9b7cad4d3473e8617385a634eb12c0c4f636ed006169aa9d8a5d80ec4f9daa7069df63b5875db8a0c1abb55d7ee2c85e0979e8d54ca416e67f6e364a14e4ddac7ed131753b340a28c87bbd25e68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fee0480f9ccfdc73ccaec9afaf20e7d3cffb1a595de9295b38b72ca008abda8d2c7bb70480917c57c0e8520a9a6c14dde3f6e25d6eb438c4ef5e9c2a1d96951a16448aacfd73e8e4a8760e55f72113c2da08953b78b873fbdc076658efd30b4aa8cb086c01245ad68332b19cba34c1dd705fdbeaa37371a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf4cb45c3a04375147c8f204e4de2fb8d615ef7d4465f2fc4f7e34b099103af51c40457edd24b7a1e69a7ae82f54c21c5419dc20dbcba7be0fca3411759f4c2968405c8520f3ba20512bdca3fc10b267c25026a1059212902e79e55439375ca16db0ac4d094d2ba7d0f67b0801948c69baac0bc83331bbca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d26e6584c5c14a937172ba78abc564f21a58c8a1e2607a34c6bf49af6fbcc4cb38d5d87e38689d10340387b856eee76d88447bd01867eafe88baa7cd361815fd93e00e77adba0387d732a3d551a1b593f3d813e31a45803a80857a228ee0446c804b28010d72b6c4d72d9cb7bec86715e7911aa9967c4a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5326f2a513713a8e7490345510299f72808a53917cd7e3a70cfd0bfd2f1d1e99daa5af2585c44b4f2c244af45674a1033593765abe298109f321a14e664d1cb0e75d3f17d3a083bcaf9c2c989df6d52a5bafb516be74e50058eccb6438d01831a566f118056414ae219f5baf39bf8201a803b5fff6fb4cab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h464037614475f1c30d92411bb7f9ef15b82508ce72df0bd2476b397ca9c5085523d734de5eb779707bd89fdc7eec1f0046874414a139b63a6f0948f117d5eb44866d6ba0c9844fd3ac0d5baa9748fd849d9fac94b7c2238a0c877104f4cb8ef26a3aa2d132012ca342804de55b92f082b2b3e55d26616455;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14343582a14b8c4809edf01290d80e6371ba61efb56681379805e6a60df2096b8565e93383928ce6060599210f125860e5cf2a8c0189023b9b2f2a443ad429469da8b8f21bd2453128e4182cea606393357c0837e6c0480e171c122f3aa0772fa755627f2619ba11977030e7ed6e66cc5067120eb873c31f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b41def7026d09525a8934134ac4846bbfe2798e6b4f37ec5711a06eccc94b3bf58bd6ae7c520684d712fe87e8507bc58c11dc91e7bd3d1c4a96356febe62c4c2fb58b9fef7a148ac6e8b205619910fa95e76de2fa1cd878e0662bc09ccf549bd04b49a80a4bdf2656f387e30a25d9deb4adbef70670d2aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ba072a3653708447d52fc97932eae550c539c7ce364f8c05518c2361ba1cec77adcc5ff403eb190937d569e4b47d0c82dae3dc8e6802b2f1447b4f8b8441e40ceec8c895d295da1f01af413d7555756da8446153d8ff94d96423fbaa0f339144f2d3c6ee6121ff96b7603677e217283e2a006197645a2c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f9ff2fde97961079a08ab9ff7a8533601e8504764d2ee99b286d3013e80fbe58547c47ffa43059efd16c7eea0c13c4f4e6b973669630fa583680b1befdeded8fe04e9e4f0d9871d7761d451d454ffe9917202059b5b7eaf70af71c5f244e1b07c73c3209e4b540cf22704436d0e3d08f77f25a4ba75bc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h482f1862586b3548ab568317bb9a5eaa77145f11494ae5c33554199fdebf566f0444f323d9bc754948de8435db08102e4e0c842a260b5fd09d1f9371b95fef5e9f5cd24ae74801acd6f02482f2cbc70e4500a50eee34409e3cdc3cdcd2374dedfe25e7bab7397b7190493e264c6ba4935abaa2c3f8f6906c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c438c314bfca7b9313e61ccd394fd351b6eab135147c8e969beff233279938440784b71838775673b507582d28009439b2681f07d4249c5bbf10c0c4f7e0b328fa96a5339be5a993ea837ce086b978f5968eb90f354d2ccceddcf21ab3168f2160d178d84d97063a7df0b062c36e45cb25e4488fb85a1245;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had38b87a134957c12e7882b3b2dd1db1072a5ac4d50f1f83e7ef612e598e96a2ab873a5c9b6ad98850152fde92c5a9c6ffb5586e86440697d66824e1037b8789429a75efc76474408c1e01f58d06eb8c0365b7362bf245e398b5be2ebde23eae507e2f417c52e49189aa49e0f3ab29b2e9d9ea4e3a0f41a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0e793091229a40d98f59eb1cfb3c3be73a5d18b3eff49a3ef39ec3b5d0d1b34c20fb2277b72d07bd3cd005a8759c844ea3d265519d696d74e6812145ecfbb8de9212eca0c36e2a249785b40020723346f88fd210f612f690d32f0f9626a6df7e75fd2c4ec630c2d3ea8bcb6f32c8bd4723c6a462f1cc7d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adb31c35fdd348c7b76a0a0ceabbc99742b1e7d91ad9066c815b0a45279895d31eed24610e98d906a187f21a47d69b03a573ad198845bc13285c207188ee46b20748bb2c74a128368e924c80e68185deacdcc4cdbece646d91159c77e55853d202fb7c7f53f0de496ab921dc7c11344f0a4a2b0e34c669a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11738857d6196eb93bd35a3927a2ba415138f1626942a06ead18f4d9d82c7bf968afdd1b867bdd9c71a3f0e0d261575adca64b60d93949b2ac8ee247647cd443a2170691fc9dfd2624bf5f1cfb08933d37dae1ee15ea22fe3e45d1ebb0c348045911d17554bfdd6c485dcd91b39efcc9bdb75d8b82826e56a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0bb50ef16d3f886f8bcd7cc300a77fb991d22c3441054a4653043c89ad33d283c75cb4722a31ed768828955d6bf39757039a6f5d0b5119e929fd80aa1644d2b16987825b996a469b777b83e3118c409953f5b4e37d29601d6050c788dad64bd4677a62c38baff50f77751f2c1bcfa5d9a2568627a5cf38c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d3d10a0d972899e96798435382191b45f3de48392345c07eb67f01d13c0b3abf95dd7f51938f90a10c6a5ae7c5d22ee010e5defb032c786c0339e2807808f05878e8a23a173199d42929cdd6b7eaaadacf5c20260525e9304e4d00d1d423c3bc010318bafb5119acf155f0949b8a0e46260235f9eea2bfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f7e0f630d3386637f6dfdfe9a9677a81dc2d41cfb6000da0c55426af790ef2f39199193476d91f18edb7769ed752bb9fb232cccc7a0f3b2c8beadc62b17fff80c062bc1b9ddb3f382c4d329c9674b05529226f9b78a1790373f2b05c9baf1d32314c343447bb64285bd040cef959681f6f2609c3fb6a9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5c92ea11bd71e44b9b52fa27a53388ee6804189ce705248b9de2d42aded1745bffc47bb9cbb0827ec33e328af4a4c8c553a690b48f62432a55557bb9242c5e7d3d91e04bb7b64bec47818e52b6ea924eef6b2f9881f1fab2b044592277769870716c486ecd817ed807b19720f2c20f82679aa5fb80b1912;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0ade1a9e054daaf2c245a651eca0c2f373821e7f2e5664e98127187d32b60721b2380bdd5a9756e710023e2cf4ce1890a45dc95038babc0ee4013d419e5f146241eb7995609bf479f51f4919c1878f236b9fb82a8171231117140a93eab1b157b735725cbdc07eaa3b62fc446b189d1f7d9010e9faa3d8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f002264dd0144176352d82ee3ee655a49f846ba05c23b38571fb4f3f878c7b569491ad4ff9a83399c1090eabaaa50e04e9d97b4b7d78679939672b90b1d9f3b35ff1cb3c6327c15f50539ee76607e9a1ee671f861cd7d3c768cd23888b708649520929b28dedf6340f24672ee1feece198f383decdf6868;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128da7859eb020f5712e59e9047ffd77833aa88bac7136097fe2484ccb258f684590aeabb7c64626beb9a2afc5435e057ffeb2691cf38bc947adab8710964ee637e1cfc81456d5630bd191305185496de9fe1eb91918af98d3359fdbe0cb3799731ede9ab1ca2bc9dad708d96bf486819e410c1a71e8a4785;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c49e5edcec4a0a0f0b35661c3f2dad3a811987e9ff4fe7edf12c5090ceefb4dbfc19c6d86e048a7bb0ad5ad401002c82f5c27b43ba909261cb0e144bd303660c31ac907ac0e180641601574871243622ea23a66a36f2450c7c61d96adf91f249bb5f40026363e9f941470837e82034d1af968a3e5a19d4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc94933fc910f7117ddd367faadd6267be8a931c72d9103c1e1b4599b97b13b5ce6c2976be7ee03a5b36343afc9b8f7dfa7ea49bbecefabf32093e3f10022af1c81e4899f05b6c6fe3842851f60df8863334d0010d147cec468bb38a527775c825c1b0bf826ac5b2fb1d19caa49be72894f1579a0d9f80c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h859593a14f9a4e1a79931bcadc9fb956064e8839f71798e7b92436a4dd5cb07a2619f779ff70e8c16f32c2e0c0afe69f55056f523dee50207963e661b555ec9c37bc3ad5faca356ffa5f31fe055ab1a2a09058a1af22db8365dad612922a58a1f465d934759523f20695ce9eb1784df756968f0c35efadc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7690c84fb8f70686d48b0a244dbecc19e8da813f4715ac68d0978164def139942e666577d5a2b26145aee01e6bafd5a444ece5e804b2548daedcdcabc3def24118e8ef959e30b95397518a29fd9ef8aafc35a2fa3560f4c0de5b2ddba0b4ad08a61e04bd8f0dc3bef2ef630aa7d549a0c89619d4363f3a94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e5a2ff3f8ef170a187cf24839be9ec43c7877daa4588323a020269fc5945dedc68d9db208725affbc62162e4793d9e7bae51eebfbdd2167da44db08fef1dbf49e628436913a678ae47177f700709b24c5d50e15e9cbb7e61818b4fdeea439bddbad8bac2666350bc577d74fb0f88b7f07fb606d772d797c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1374096386bedd81b04183eff129c372676d27612acb8cfc5537bd42023ff337972b0a0a3fe4c80055e325dce5674b668cc1ef118c6273112e44a600f75cf6bd90f7015913aa87aa1ad2246375e23e45ce1223b13bc60542a7b1ad93e0b6bee64fc80dfe0b129c41d0450d216c7fce9e924aa07889c1a76c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50d02df8d9d1c4544b5ec5bdf7fb6c5bd66f8c4db6b2005debc5a81239885e59dd6e1d13340c82eeedee7e81b5fc7ffdb02fc6db3e4b0f016fb5e56932a9cd7c68c0931edd4be298780e38d9fd325e18f98b1f3043e5303ac76d953b7b5be00eecedceeab251ce658c1d12b9a81742b797eaa23dba47ca3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc010adacc906aaa80ac47361d75f0631db483d47b717543107b185be3ef7d58bdc1667e378af3517525dbd33b04afe26d2168494a5442d526a7b46cfd0a2728c962ce209f40a56436210626ea5d2fad93611d69818d01bdbee7856dadd2fb3e9b86dd3bd3600cd689c3b0eda76ae32beab59a7a85889e83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bfac6278db4299dab4e5abd8357691d0bbf2c12e0ee33c3707ff79be61a31e438cc7bebc24bd0c7e19f266561605197af4261852e17088aa30a7c313ff148867da290e33543cbf1d2d7ef49a81a1824b44002f4236c5d5038d3a72c8d8bd5b940d32bdd567409f84bc1644212779c9f2e0bf7fb009274a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff5b6a174c33179922a2ee041bfcf2d0507b2e4d1f58f60c552ca9df42b2918786260ecb66b8e003d3e28142dd5e0e6fa87a488f4d3d794b2fc74127060ba9722f3e014ec0bede8aab2b18335403a5f0ea7251d41560ca8d8d86f1986e3c6d1162e533f2e08290e8c82d0d01e3ea5d537bc9980a41fc36c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h292dac132829159abef45e84c81c2d1fb1f8794b958a180a3af35fc7d1dea7a4ff37c079284821e164b7e09e53be1de4f2c8e25abbe8ef01837fe20418af4940a72cd0b07a40ebf9d4b8e740ae81d1664a4d0f443559d5da7f075f080cf314fc8c318916d300412518a5547af469e0d38cde8b6a1bfc7e01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102f28307789eccdbeca03ba56a0b1b4418f87dced1173819e2ceea59633e96c0310f3e4903c959ca1220c3f6c1ac85ab5ddf63d2c63af90b6a27752fcf09faddbb7beac835f398ebfb9a3cecab654c2c22c83de622f5ad039d4fd7be16e54f61f5fa6caf0cc63762263643fc26e26970a6e0c41302435b0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1319908fcd6098956a2b49043e3442ec21ce39fc2a76b9263a5d07f3ea19ff0f5496168286257c842a4277078ddde9e2713a628f8c80be1c99d8d7a4d0a56c550df78a46d724ab752b8a074802e54a6b41cdb0c0bcaf25ab78a40b43c05e87468a6b66cbfa877a0b243a2d9716ef161af895e171e37ae2bcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108005ea6275fa60aabb20dd1423cc67cd67e9a4f2c85d393965d31c6dab728be5498eac5604322b5f096fee01eceb4e196cec1c460cd9e5539fd2ad77529dad14c67411db8ade54e0d5758caaf96d7801551715acb3fa2df0eedf5370213210db3bbb3046072abd311a5b3ba57b03ec8efeeedfa576e1dfa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6be53c451a7de47f52f9afa80ce0acb6a4c78ffd0c075b2c61adaf7ea4dedef0e2e94a3412a3ffd37026221d2309e15b62be861be484c117d6ed48a444a0747a5a19e33f1b07b820e3442f9bcf542fdfecef438411613a88c6ceacd3b7644dd12c54b8db21dd921712a6059ae4fb7271019068fe05bdb9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11843b3b2c5babe190213c05d86134060c9fdc26d11947d675726da5d99cf154ebe077605b6229bb9fda05c7a4d797ebbc022ce0929a83ab0d28354aadde15a25c6253388c662dc13ab12f3f8ff455127e9a28033294e64274ecb8ca75d060168639005ce2018158c34e05b07a385f37005d3d7b7216419c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20137af575c7dfaf3c890d28d0b9d99693e80e4b9adcb3aee383e938b4d232547f7c8f07f161dfb4a9021741c389ed1af5122d4b3871e06498522e3b3dc82c7ffe0cb8938cd3375ff6a6ae04ac613ac41b15e6f2625b1ae2f55de61d29b835cd6d74a4cb0a660814e9746108254bee4e06bbcb4485403491;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d2adc6476c345692164eec6293ed752e325a93fb79a00ac4d8728ab7353ee7a0419d469d4ab1647afd41323ad2fa009c3b466739c1c3009538bd5523e93eead11f461c4bb86e91422172b0693452b4580a4ccc1b81f35087a653880a41d5550c8deefca6198053da5e8c59b443ba8b198345fe0eb03dd08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf922a5ed516ac560e9ab393434db5ab2e24a3b0c84d5be7974e70ad6cdf27ccf213683da9d9e44f5fb5208e67e667c72c54461f1710a07c41c3a258108c5bbbb1232de5a595d950f8cbfcb887a5882428f1eb5cf80a8c6e65144b9b6e0832c05958b4d73ae188ba3232c1f67701f4fc64b5da0ff86ca3838;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144a10505e13696ae176f0424d747c7311bc4e457b6b77a1ac4d0f962df185ae80ee834c8a67f660efe03aeca2838d43cbcece5d80f06cd036b74fe46a3d2b10464a99c31fdb2c097e8b63faf535683ffb0aef7a634cd11a8a964c078cf63a018a2bc50b87e946db8d262678b12897dfab94c85e88cad577c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e9d757186fd80e74dfa0f1c4cf0860e206cfd282086b9445ddc70b84afe30892587ca50da7fc7025d0f963f55c052a6e5ce0a41d61ada6c7b2f0a064e579c24af7641b970e89e823314f4850d1763b818cb996026fc8c312169e34971d8d6e3b4c9e30bbf0520af0599b2b0c0c26d50bfebad3600e791b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4572c38e779623236a59694478feb1083dd1001ca20c222382df69381538e5c59a4460724d5cfb84cf16f2911f2b5e9e633f4166e42761e3de93cd5223c480050d533517456bc8676072c963cd8f26051491ae2aadfbcc223d76e30b3d56e2814a5ac380c250591f73bc700913790403c95002ddcbc02522;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192438283d1d6f8ed1564c03aeea1f8db2e37025d2b8f793026b6252d999484c0281a4dc04ab49f04989b23ba5fe32c130ff8fa9202e57c9394defa3ed0bd59c3f1e31c7acf725148ec0c5ae1dc3060e08578a5dc2a504f55a47fba3246bede9e7d8f21aa9d235b7259032e48659c1a5191c56d57a7789fc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7e76fe0dc1c5d477031b85425b080a986c1a116ee8ee59676fb06e264f0acd82dbe024cf7a7e0e159f28eb7f543880575bf4b89e90bb676cc4e3a91365eabd5a581c1689316008873e764d6992f46840cc37e80a3f47a3265746f6d6af1e55b6be7c780ca079d62b88b1eefaa041fbba3e11d7aa733176b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13145fa9460f6a94ab1c2df9b8620700ad2aa8bae39de73bed2fccac94132e2d6b5000d60419d3f618f53b37cb2321356fea173b6eaed8d6510b456e6cc51d47542f1e4187bac2d459dd869b2db907d29e2cb5967c1dda9281499776906750585dfe0f75d0b0183d9beb35eb60c780173e3c57a43ea2996b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b25011f5948b81093b3f1727f48c6c31f917a7448273abfc28b6b33c03cf633769fb4f443f42a0830b520d926bdacc0281cef24f306d9bebe77c67f7fc572b24277376931bc42329d77a5de1cf2ee03b480f5bf0c2e8b4f28a25c5cb6ea11d03e1d79b543f487be56f2a3a695758cb7e0b9d270217a74476;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1352e7e9f642572c7d7cea98d7290ff15f6b1326a9067279a54579c75879451178b746c4f5081603b1bccd425db4dcd4531ad7778984124596ca8fc3a8737bcc6e272f7f919e09a63dd6a28f16eb239d92a3449c9f884852e5317f37978bfe9fe1e3575dbee31feb23f370b1c74531a649c381b395bf369c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1073fa3106c34db7e947681132b6da56a2c197fc621a6b435d4a036adb77191dc661297cd381fe1fd59ee410cd791ced1e92c19e2ab4ce87f730bb7c69a688f681894e9f05182edc40fb6c8464fb47069cedc50633f7e9227382e91cda363ac9142ab576807a3ae44b6dd19017591113fd2ba8efe465fd1f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86f97d37ca7238feaca734beb4fef20960a4d950b4b861c4e81726bba6a4d02e1614c43bf0435963d25b91d2df4f8e041f65572c1126925a089119cc22d32ad8bc5d0a9e33ec2176bd007899a1274974f75f95e97a8f4f22d298cb26a5f5ffa129ae4982b6e2dc1fd66b82bbaa65cd4375d68027fbdd01a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h472dad5cf1bc97b22c6c9cdab7f2066a752763f89ae1e567b3e06793cb9aa2686a40487444c2277e3ff41bbe384b8de44bc39d2f81b52cd40e3f8933a020db4ca9318490071003c05ea8f684e51a094ddd78611464bfd6451acf2b0fa543d16055fdd707cdd0c9ed3752042c8972bd2a9a60cd79544c331c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10eaa1afded89e0467954cb727d73624c5c9e81ac322bc23c2d356008d8e4bbfba190d4f7991d8da4c31246d1cd65966f38532670d4394f3ff3ae0ad9558a0b992d69f3ab828f46dace292ef7a656a07551e9d483e90adec3aef8d8ff4118699aa738db420cd070c4a08f70529e0a1250c93eb0d54e24fe9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b322b17d47418eaa906599168349e5006004d81c46a36d1841207f9d0c703868f8ea49ed78367dd983a22f7f6a8a97dde981ccaa63bdc44decbe3c08f7b8ba98fa79a40bb6b66af22b7827a148b6dd7f4d728159e665da05c58ff6b6cefe185ee32f22daf7a836714d67a9d64f57e69d389cddd1e0f07bd0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17eb4e3e1a9b2b97646856fceb19a1f8464ad41b53d836ead6e7f844936f8680395202c3514ec73650c573457de7008fb719292a2882d233df7936406ced89f8eeee9760090dac8cb47b6ce6672b31fa9777868bd6d7d34f1b6ccad274f0c3b026716e119b96b5475668a80be6c4371f75efd01c43706cdb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d256826b8c5c6ff21bb36cd251cbb6ede1c72db1e7874b4b1b9f85db60bc22f34435a39aedfff5255854c8bf9348715b9ca04281f17d64ce50bd108c427723f3eae9c36c195234173c22607c491d1d000b19a86088a86117b2dcc009cbb2fa9ada121a0c78946a9bcf482207e36158f9251327f7546aaa48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f93b5525608b6d3c33e2cf00dd7686c5f3641c079bac2dce89416ceada4a372badfe0cb76c5e942d6852304cf12b01b7e97c79a9aff2df5252ef0f6ae5eeb3549a0e15a2c8bc51cd14ec8526bb32996ed44c306778bd226f1fc842a9b7dda803417be65bc53369c960dba7150f3a1be82eaafe2ae0b0f4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1996a8abfccc666a05d38b3fc0b7ba1e140e87ec5a6752aa175cf025faee5cf5d051bbb45b3e015824732a35cb7c65ffb055c8dd0f5210a4068c813d7c9e1451f33436e8ec75dbda2d6d995b8e119a8d849629d1da450935ec4e4ec4ac826158b13c18b4cb8daccf50c27689d222258098b8675e91fd816;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc308e478a7dedd0c02721f893a3d47c90a791f47bafcd83bb4fae129f024862ce0b58cf41402adc74bd6662da2460f664bcc622255b53e720272fdb15dc91bbb49ff91ceedd8dfa457d7b22f94c981ce68c1ef4b17b9a459ac678912d1ca9f1bc03e35a3a0215e92157caeac3c28e6ebe2766c413ab2a884;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90561b8dc379f82d682e57b22f696a043bd66ab57ee7ca5fff5a7bc39d44b774b8ca11254fcaa80bd0b30ff79ce5c04bf85c83c13e4283363e257e9a2b7401b01a70d95ebc0aab8e59f4e9e8b256a0b6cb2a6725f9590f71521b8ace9ec160ec19aa9b98e5596b75d1d007dbb6cc0ef09e916caaf809d6b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haac7109888011df2243eefe21914808b09582c2c64db4669373994080ebf3fde2a35f483cd8993ff6531208cc5e6b18bbcacbf002e0afa2a9f933f6f32e7208eb619a9a46b465d9ac4550b8ac84f58bd08af3342c0969d8c9e278caadde07e0abbf2c337b350d2a1a80d059ed0a132fa59d67f80a94b36ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd168dce062388279a5d781e2726ccd4e3ed73494b0c85745dd682b804d5ca6584396ab97b3439672ab53ef03edb77b0e927811370962d6c7e64780eb83b31af03622fe1a505d3872339efaf05e4bfc23ad2e9787cf99105f264cef3a0bf78eba4eb9c39751e2f2f11e483d620239fa26fc2d95545d586680;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d722b6a4eccfb9dc9de5efd81aadfd2a7e321a46b2591eebdd0fb43ed9a544c9cde8f53506d833999a9c62f6d8991d1bd409ebe4dd230d9205afbe2006857c81be9655e204e43e916680e32d6119ca08469793787f89282d2bef6ccaaf89c39d304062afdfdd5c8eaae2fbfbc4bb13d1757dd0c1e8ce7e25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172389c7c2b85e34edcb69c90be5120ffc3d1fb4b5e354843042c15487f930b8feb3387d44297e92dd439ed30ce28bf3eb4f56657f8d460d74ab898aa0471c1515cfddc7b781d36af75b41f8fa269f67a2e8adb00ef2ed4dc3f324c42a6f4584b4f8fc66173091fc079bbdfe4f094129162aacb5a1d838320;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4ded545a9b0ab40e1c67b7829001c39488f6afb0cbe48b3a0eac43ff9a6f3ddfeb8f47be51be80df7f504d994fde68a7712e06aa51aea2ddce52b871ab6f1ae6cd6aae645b8d0d2fcf23abda21165dffc6f489afc981f0c111ce455fb9669974337ae64cb36f21e357e9604e554c84495b33aaea2df121a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b706a988079d5464a75f5140027ef22a307c6dbb02b308be01ebaf1033ff4a84a8d2ddcb930f5d875df8d33d71c0029825bfee71778247f61d03312c20eee35f86ed22da2d6b96325e0e4fc24cd3c4032edea43688118fcaec390d2eebd40771c0446c187e1379e36f4bde4471ea93b205f021f989a6c96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a2378302a007c0e4b22506881a082aefc336a85e99e1a487c6a79dd56d82cdf4828135e31df8ef52c1754a53be2eaaa7fce46f56dc615c328222f0de92001df81daeca8534a4a053cfb2b5e73ec98962437330ddd979333875accaf15a2d0ed13e7aaff62a41f0d50c253bd6c591a63bb9f2b4e33453d12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h442c61ee3d6b6f1175d5679d5f2b06e72c767094839c4a86cb947a05cf1405678108b394d9942e9016c88b7292517c8695cb09d0612a9f3209f4a26e1f19739dc8753caf68537b22021cf9c210c091b8a0adb7a1446dbea0b53f58df89fbe20fdcf1a3369e553a24644f9c7d0228ee05767229060aa07b49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b198e6061fc98f1527f7c1c3dd4eff5b2ca80d2e48d75f931f401a40123d5813d57d8d04a0f9ef3e7dbd831b2c7f2dae2fa50be0f2a5dfda5cdb5b647b4142b62dff4ef90cfaef74e5c926c336b7318ccd4633e3c0833419b9f53567954091341120979d8fa22472bf8fb7c37bcab24bbf320f28539807;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a1783bc994f977d879f7f7206a21aa00711978935dda333acb7f1512858ef3d37265d44c47d9302ac2196de0f1cfd7811ad6e08076a23a6c6faf1ca68ec2222406a53a189d51fba6462eccd87fa3d8bdf6d8f2d5004e25321f38dac6306b157151854bf326951799e64bcc3cec3638a0bc0af594dc63bdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1488ce8f28f4762ae6786872658559b56f2d4fcbf094de57ccf2e7ffd28926a0f3f2af2e1918d6e825b708abe4fca3ddf2b653f0f3a1f83be6144ad48040fd107999916a8e04c472b4bd7a890c9670a250d8a071afa331fcf630b143d835ee79552f9e2b7f68215e9a810bee5da79238bdc0fd7b7205d6444;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h145f29c802d372532ebc968207df14d34627114f67999f6a1c11ceb601ae3f0fb98618128fda59607e0ed4961a74755bce70d87701ee5bfd54659ab948e64e253de770eb7036f483ea77c1770f771a0e88d3cb3a3b82440f15dfc707e33a338f44547446dfca216def0b844c6ef21f8161415c5102b9f489;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc884fbb01d9a640ada2afe2ff06b33f928ff925013ce5f000d53ec054660365dbddf0eca95be7172f66457323dc5b357eb8ae26fb12bec3d6bbe310661e95c955327ba344c4eb38fc9c94307078625eb927018b148eec48655501200c0a96bce1afd9961fce9f5c9e8ec15bb86ad55ad0b242cdd45398f66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h849d97795a7590afeb14d1740bc6606069c2c8d527af962a975089dee4b872c0bfdcfec8b847eb585315d20522dbb8beec1ae69f0713722437c547ac69b7de9c58b180f4756b9dd7d77fc72060b2e171fffb98ba274e0112227a6ded2d9d32616dca6d71e2fb001e5c4c90da545cbc612660dee92ceef9e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33918ca8ca0aaa7ac553dcb08775095976006c52cfd0f23d20a199210f18510d465c696c6b16b31baa90a410e912e9069874ab55aed6d15a84b9609e3ec5847d9ff82b92f0e4b6a9b659059e747e4ef6c23a90b0c78d61c334d2e12e487c2fc1abaa0698e6d51650f09a1498084be7a6e0ba36373535ef66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c99dc799492f88a958a295ec606671dc87571c86a5f88feeeeb89d99959f8990aea1ece371923e5f8b739328cb45a85f349848a932612ce7a64b8b276d8d131b0bdecb0e8ddf980d1ece488063ba03f755042848d4a65689cb098a0616b4e11d299f85d615346443f96711bddcc1f3807e1fd52977be15e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179036d2a7b7a44526e932aa35140905a102cffebe1aea930c78646f803ca47aff2ed7da4bf86bbbf377154086551b71e5112fc754b20ad685f985b4e5699727fbd83d3df325aeda98b46320b377a20b61ecf673e53df177b4712d6599206e55de60af78732429259a781e270afd52983f453c047333aac31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5209ce3d50f2bd68492d186adca9320b2d5d467cec9eac6fc43a1d13319de8ddb4f1bcbcfe0c279a5366dbd454ecd4de93f61a3d0745352921712e28286e605c642e82cf82511dbc595679b805e7ad59097cf52bc739d8590a55afc6630ec59fe9ea256c26eca58f8a0fa193e9c1b2f2cc9a3add9b2a387b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4f9a15e0c43e3ed23257efe18c747ddb3987e9636e29bcd2a5358a588257809be462d47e4d5a446457fe40d0bfd85e7778a6b08dc7f9a8b08988f295b629d27d2c156a61618582b02a1a3450bb6e88024d0abd3c456dfc4ca9bd465a4f4c9f555016866a37929be3dac1bafa1b1a19a24cb8120e5460388;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d97feb35491b06bc9b43ba26803a6a179baabe189eeba8c46bb47e809f93f9c67053e4f9485a434c7ff5f81f58eae6dafb1adb1fb84edbdd83a7cdfdc82cb28e15a636f85531cd1a13fc84aa0e61ef97be67249bc6d1a18ade5aa3321cd873373acb7bfe08c41838404b6c09e4cdc413d74e13a6c03ac4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f808f8c8c37f561ef696773f3078cb47fe8ba58e9a4092a437e1a91d2f35cbe511bb4ad2fe5f937ba9df995c0901dfa5d722347bb5e592ccdfbd7499103e33d844a08880c50f5e695a38d8068fa1847695dac334c1b41c64cc1c52cbc0e80b1612225e099f1aad80d993b54ec49aa5cfe555880dbfed285;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a935a07912c9ab523e8d786e2833ad81764843fb464d02eaabb81f1663dec4761dd5c2e621ef8d9e5944d21129882d93963831a4594c3c5d7e4257b6c9d82b1e7c65789006ebddcb7bda5de8dafeacdf33343ee54a0a2f8cee283ebc498212236effa81dbf10ac69a839397b756b7072bdb673c1628d97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f67297fda17a4ee7e7c8eced65df08343052fbf4c9c33a1b4b7aefd5d0160da1ea2b2ddd1296e05f26530e06972f8555e17d5dcb7218495f2adf1f2faba8b4af54ffe05757160db366e6c62fb98c09de0307a4b7a563fc8a79dde9219ad35062304179c66edd181c6fcee992a54a12af540d536c6dfcf83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1258f4cc69b68060b9859c1721b95d2686856bd1ba8bea5128f8cf5f2edf4dce93c24f6290c261bf37d539fbae38ae4bce2e622b3531a0ecb2c30d72d66e0e7c337e91485bd222fe8b0d38e19b8cb2487abc23db7935ef66a3ef4a8d6cbf655ef09637c75c12c593e55e0037d2b7ad94679f45d9f621150b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60bd53c045062ae7d0b1aa0361de9930cf22e24f80deb910ead831579513046457196848c73b64ab13623a783d310762ad547977ba61b128ca9fdfe1a8712597d7de73244796585a16fff92b0ca9edd21d3512b402d4a0934debaf7d17075bf76967f98bb6d868549df426eeaf2b70c17c1ca94a9bf154e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b5ed35c9dde0e00f1ba33cc011d6225916c1ab2ad7051a250bae51cfab8fe649395b5ad9281039795b8242e64555f341004889ddc55854d2b34292694a4721e59eded82dcdc93cb1ea63398f922c70ab1cf53ce571cae4c93ac33c7bca816bae5ff4358b1ee768f5431f20bf267b211ca9a68ba71486a17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138ea3165cc1cea25f503b3edd01003e4e3ba7a09ad7978ef1b6437aec1c7e59392c713d5b5e4e209be4aaa369cdb872927eba6bb8a0074a453a5c441cb7780b9915a1e44c591f4706c7c4677a54455c53c26b7f1fc1671449b4df22cab222352265847fa65549cbc6c45c88940a045d2964e90c930b31aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0e7a99f28359c43f28affc7846a20643f813bc0da0768606d712b2c3489f46d51dce9115f674c089a0fba0e61f273e8dd387d472054455b61405ebb9e9492fbeb8c8ec73df89fdf615c4cf599e8170e57abea09bdc5f2611923bd6b137b5e5176064934e1c8ceee201728b6ba2d25a5340c33b11c240aa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17187b4e0457e35a4138ad156914cbfc97e877fa0b312f6894e2e33547e308f4f403f9431718a31240879812800e38caeaa72425e935bd51087a65109d8c88947b8d185f0741a1ddf45999f0105f96c4f0ae1be7f8c6eb0495b82c504667368689906f97b4b6512506579086d7b7ece792b97a17ca98f18a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c5ac57c9e9b1f88be78f8ab6397d1f307fb24dec828740a4e71acded50eda5c0e751099b0978979730fc9bf8f2b21f5cb67d44d507b976ed048b2be7eedc58db28afc95d688578992958eb0ed90ccd79b476480cfbe7c7e4c4dc1ce45e121e5607f821b7bbe093399185d941c1709d92205e0f17f3f1896;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89867e86e7561b4628bf43309a8948fa9546c85d76ed908767e29ce26713521540b4d62d6d650425098388012c83b3ed24252abb4dc187985883bc1992c6cb72114c3832bf6813128c7ac4e0e1eaae44d631c691978bc1c3bef503137541c25474fa16f249990958c57dba930a7a209f8e1ae9255d3783ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9267fe5ac15bc3cd7badd60ab0d86f9e9a50f2a886169d5ef96db74b38d5bd2cd8aa4713ce6824c2ffd12f33df648dec8c2e7401310759f31cd324ad404dde954b43462bab492081dd9870b3096faec665fdcb1d212cb558afd063108cae3bbec92e03d52efeadb5a75654fc1524e77921975dc1f2a189c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h491b8d92e0ee48a8d5082ef05bd8e11b7c516ac7eff0a9acf864fabe1dd03d6a3b7a527bbf9a3db51654c6d8e2f101cdd34f24bd3dcfc169df04bcf61469f78d37d40626e5e7fd46976ae129cc217bc99326b46ab4e05f2e46a59cebe6520ededaf6dde3ac750489f5b0f379cab4776ac54aa03c900f6302;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2eb80bd3a2167007b2a3481741966b28d9d9b964c17e727a3ed0d46b731dc8e66efe12273aa5d0e362ad6014de0fd99e0b650b562397931dfc0d7568fd8a43adbe87000eafcddac2832230135afcbd4eb5278dfcccdc419d498b0703978650b1b0617cafaec901cf93d6f1e82ec45c568d7587a072a354;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90ac60308510c31836dada081ef0ba3434b73cd5c4825f052fa7011aa6a0c0948cee9ec177f840f3d3a61d3c546d70494f4587821afaed0cc35f1f806081c73f210bcdc6bb7d82706b1fe6424fda2f073088280b36044dcefe78d524bd95a6a73a4d2c51a884c27be4d9e7f00a13ca6b749f8e546ea92ddf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fcfecbdbf12469868750cad9f5f55876971b665d881c5b67413755d6fb9101f95a088a162154b98f253a165fdd174bb3d7ceadb9c07321e73ca47001090e443e011d00e9762c4dfe1cf42d5cafadff418ca76a8e4cf81b72a9bda153f7dfef91ffad6f7fa20761ba3f09ce6dfc9fea23d92285e9f2d06f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1740c9df524c42141392b3b4040e70c92107200262cc3f36b7fbb0302a818a292df6e2694445d944e6a1b6ba6962a00cba689f77f45a627787f50b8ef26a45a3e4dbfc47db88ce42ee8b813e71c3d2e4d117aab0db7832e540710ab5f3c8e2d3b59d50f6f73afc5cef41eb9c4c6a868dd37810b80a032d84b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183f4f67e6b6ca34f731ea4b947ef96ae6ea33caf8f668bf28ef87ba511d9c00c179c97b338be04c653b4119a63ef95f07466eac7b2714c0bbf2bd1b3bcd89cd840ae1a4c832b0a9861039de08449bb5503da82f998420f08ac9a1c415b42e7d5f430e334776905efc2650b8f3765c141ae94cf398129ba16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7850da17645516a073431ff48a6332f7b41c08ef772451ffb9bfdfeb7be9c4850ede5cd91efaa7f9c534feb0335f17ca91b69e7629d483d7381a297c4789a9cd60478f33a91356a51c1fb0674f27e99beb2364a8be38bcd3e88f921d5492cacb19551023e8bcce7676d1ced81101aec2690771acd0212f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94dba837302713126b408f772c523af25504665fb24db84e17abf62521383853d0ca3411f8d7a1363eabfa82c905f5a547b529a5a1ad8a7c525b5ff790a73ecd80038be541f5ae9d54485b06244a261fb43f45fe48bab5c20f2d75f5f4cc94a0822d257ed60a0261ab65485d57926a49d25ab2b83edf43f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5248f5165a34b77145507c165a8d3731cf74a22aed1d0980dd238d56d503f41d516a8b913eb9c00e30c04e2fe99d2a1e5ea07f34e78caa07ea5131cb7961f0a7e9c06bd20c81dd19c860a3a46867953b23500472d4dd4cc4943a77d701c11447a559d74f9d5e7605df1bb77b7c43e9be887345354def5b88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1348034df744e92c3b30c51a4bb53f35482255c23b1af98256e550c41b747c727b9d41f3f0dc107a16bf4c2da315ea7b63dfa5ab0a812070f31de4c5a0f3756602457431361249c6bf5c4e664dc00953c2a58d317216a35d69d808cabdb62cb839b52c54a891900352db7fccc84c45f85c119631bd23505bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62b30ae7f63f50b8720f4277077dc1d613fa1c62465109a64c25c46ddaa4ce4c3563755a60da3610b12a1068c9614e2e82f67213d6ed4e7b78a03b49123c2ddc6ac30bb1121960386ffe84a6a8eb54ea57831ca8c1820aa099a7a5ceccbbe40a8aaa59a76753d3d85ad697ccbddc7ca7fa2ab47dc1ded994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd299b45268710cab67ef7ae1fcd7194fac05f8361371bc1c1d1067668fa06ab6c93e85b0e39d4df84b2ac82486732a86591fefeea3849caed6b95a7bf1f0e7e3383d951199f8e1be897acd0126feb3f65c4328efc81e7262a7973dfd94e043d02fc0029ca658d851a0c369c4634b47e5a72161dc9d9058aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9222494b1ce142480bee9a06117f95122975a04a308e7b563b6100a8c488caec98f354e42407474e0e531c1a8de9aba1e52e4fa4e5c9fb416f2c602d7501bae37deb91ec413c67603324dd66943ad32a5c2a44fe8a605671b025d00f71fec8b5f229aef7ac96b9ac7fad3b3cdfd34ad89aee5e1ec2769ef7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35be63a2d449b9f99b24da9bd7b7c5624cd978ef0bd40b725b3d94b45f3439dd89568a4c16fea9ecd78a8ca1aa51d46464b59291b7e6ec51659eae193597508f0877dc1616d81bc577b61e3cd83eb00337775b542d27a3863411bf203c371f39aa3cbe54b6f9352f053ec4aa5befa3c5ea265485adf0d45d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e5b5abd01cc00b8f2551c9ffbfdc991314b065758a93351d7bbf57970eabe21c22a36393e5e38da2a32891b9cca6091909cb6d68a3d061240ae792fcb6626591d041570cbdaf2dd5cb4e5486811be2507a59ef04df5189ae41e05d2eb874fb1819b359a08f4c74c7e5cc6f83b15aa85ee142cf173ab038e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a9d0850659f9ebaf7ffeab59b5b9465cfa7a2902af6159a8496aac8dee8cd8d8da33fb15255115b5f0483c4f4b5c66558a3de7f5a573b5abc570b764740f805980f7c3e8557da6b648fc978944062a653835ee1d9eb8383b1da6cf7da7141a13c54b68b9f773c1b318a5f85697222e24b4ca40aea77fa57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15791cf861606a5b3a26f71869da15d3087fc1314097050e2d9089f42060a204fcb36245a09dc2f0f22610677a8e88c70a277e22d3e5cb7e6e39c994e06bc58306f5e3d7ecd176c050295bd8805f11851d577ebafe8ff13ed522605dc833c8220475c5d1cc617ca6536ff07f20f5c4f0e065d6829d30bd733;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d218adef730b3354c0062e78e6c090494dad92ea377e1894759c88fed4407c8c10b47291a4cf77bce183eb82199a4223ab73db16b2cff002b30614319a843dcf30672e71ec549eef8dadd764bf0fed662259ed498b5f33af335c090e9be0e61414ff754eedaafe8727e9aab292e4f0a6f4424cfebea7e7cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a152f064788e9cdc0901839b59e27ff700885f5b89225773b8798a1db23d8068c6aa7dc08271fffd504b6319d71f95b120f10e6af52a7485b4438bf2d9c20ceb131762af39d9c639817db1ec32334532c676b0248ee091051193cce8a7ba75aa29e1f41653c46c2fb62edb78b6d0fec36f31a63c10da8cd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a4813f1eeb37e9674c7a7b0d901fa92864a0b8e7fe61665b7f19933a2e28d6d877e788ea8a166443e72592849b582b1db2210211f13939a34bd97f1413a1b89e85500b986437ca3456aa55ddd4bd7b75d8b209e57a37520cfa5166267242885345f2f4f6360a8d5b3d59dcb8d3cc354987c7b86f49b7e72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e9f2e915c0350687692d4746566d81f4cf8ef5313026974aa9d1fad123fecd7fe715b8a5d89ee39bb9790c789b1b40403dfe7ee77babc73600f68ba98f5562bae8b9b206376f3895081e32b04e4a2a24190420b26941b40f2613150248386f3166f7a59d014e5e77f8684d8c65ec82db7f1409da721953b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf13fb42411ead6ea334d36be68d8386d82fd05fd4ab194ae0234618467522cb47188e5dd1c1b9ec45a82853a93393ce05076f2528d10472ba7051321cdf02b1280ccdf6572d2e42bf2dbe7d73eba17a79f11a236b1a576ab80712ad8b226c5570f62a374ae2448dbea65cd5a6ed9510e93dfd1aa644667b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50d2915534566559373c078019703f8b633d0acb9f99f66e90a59a7231a61f68deb426815e47fc12f7c5193dbbacbf290a8e4334597e9b347612f424bf31b92b248581e5bb63163543bd01ef8f23d9058abbad9473ab443f3351b5845c0b707977fcc63f385a5049174d422899297a5122f4c1c4c2aeb2a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc25485f61ea1280c373418353a4b9cf07e1d7c7a1fa8b672b125480c19e658f778a7d12e34c2360de109381c06d380248de654d8ea12753aaca3718e7a37ff4a6c6afffc993272e7afff31826b04767bd98c5550b012450429421f78bd9f67f45d0e55e8ea760e12bde1806f399efff0df3b4363813e52f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198a29d59b7e5b6f2fb6b2420d3de01e4d4710d48791993edba066bf0b46de1a38f126f020058c9fbeb2dfcf7044cf19d35c5ba12add59fe23591d86e529426f4e07b0d5c7ae49275a826d37690b79f4e9bd3d1dc82fa368d97f578398060bf2e75f80181406d2953e52b7327ac1cb2300a1c62797ee02f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119585e7dc6dd9fcd137a7a08cfd50ff2ad20364be24769a021278db0d33cd132eb0df4629ac3b8cf74575280f8d71a08699f56deebd777c35c256bbb192941fa5db8617d26e638928132117aa062301a13ed456641afdaf1c656df6c3604289219d8883207d8a72d76f70506843099bb00071d5492a3d1b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c3b37124854e262d1b9c6e3de29731eae9647971fd1de76e5de42d4ad4fadb5b44a44ffb8950503867b69833e50fdb067e681030183e7451aa86d756a664d622d0002e0e16ae101d112aec8b26c5bd85b3c1e07f60e477567b75c1c1d70d11f80e1e2423a5ebe57b9a249cba3a333c292f3a34bd69ce7f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5587d6d3dd25a181a3375f2132b8abd58070d010e49ecde9f8a89b84269da86d674b90cd02e44a0ac0bfd0079dc6fe3b7fc8491b80fa8cdfb8856a0420f93daf59da2eff374cbfaf1257dc4ff2fe5de78e5e9066c06a8c573d7f1494d4f783303e00b03a5e3376a90805810581e0374501858f554fe92bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10cb1e2856bdcb1124d9f759bf64e048896cb436fa15852b14b9e191624af3d538a7aa242cb72ab62f1b35c1dff3d355a31ce8d2c9bd53bacb044f39e76014573a26c7d9798d0d6b753deec81d9a934c0ae38b964616a0ccbd40778abc51a2bd06555a6a7e052731fa3c64197231eb52251cb6a047a408d0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d12557cb5234da5d0dd4342db10de20ee2ec4e8e69bf7ba66c47f299b679b598f20b2fcc33b892495eff590f194d8df2a43532c6b9dcb2d47674a580acde572195eb14914dfa1f591d9beed27fd8a3616381354075dac0fbaddc166341ed8793c985d7bcdb8babe2b21885c47d41def1366c23c2ce334404;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9762a74ec7853256d197e1e134ac0a94366901fa08e987c5e93eb3fa62162d94e3ab7e31cd23dcddca2cc4196a7628f1273d358fac756d0f7acf6cf2af29622ebf0263d75f8f3700d7839bcf4e8bb3c43e2b4a75903c3322fed9197f50db057f3d9c72fef140ada53678aba44c82da93d0eb2b3dc7e546dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cd5b9e14fa32b232a88ef8f70a83cf6a61e35bc9b218f8ed2f4fae26e9db0c036bf07b4c54dbfb62c5624b887da073ad81cabec2cd001581ba50a0c01987d76db1f3a8bdf943712795cf5ea64217bbf85b31d888091b8db8b9aec2af16a24cead9b4e68bd89c6514fc05f05f484ea88499d4634e45347ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h206b2ff8d330c152984099cc04acf218eeb3978fb5aab2aa4876bf10ee826a275b48434184460e6ff3050bca2f87b47ea09bafb635c07c25de35f7a9d439071ff209e12084f41c02607206480d1ebd94aa30ec6c20b606b67b602d1535506bbd0c7d83762b77c1f99f4521a7f034f1abc93055e3f34599d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a2c325ebe998ed8c3344c1d1b7b9459a4f99063fd478f49596bee7b7a7ab0161f89d5cc9fd24769505f6ceab79a6fa04f53f4c48a6a68e087720ea8cd8d50f16e18e7d628e95c051850d0266359c8861cd18ef7b67e6e79764d77451f0f797f62c9082f80d82bc8dd06995a86305c6b9a0fc3ca1f01bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b91ab3466fd89e63244867c5df4df10d1f9edcfdef1b747e38be1a81f54a32b6fbbbb3246a9b1a09fcecfbbf2d74e0e51d476e608d1965393c8b385fe0d1ef1e7a3c88e167b5141135b51f0314f1c1e4a407c1e6ff20eb12ba487129bbe39fe2c72f5fb7739242eea2a251944c286fe3f405422a54f3548a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3d2d153f8c34940615b17ffd657bf638b33def8eeb0ed5d7ad8074ccbbe6caf3b62bdc269a6272f5e9bd7174d96ad6d5f266a75cc0cefaa9093c14fd2f412459b93be0455fdb4e3fbf854c4114f2e5593f162280eb1105f1ebae4e602e5450e830b7b5e0db008d990810b2a29970ae26956a17c575f56c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0236189de4de64db63c6ec719d7e99c55befaf51f320f845b00ecd44c68ccafc48c9029c0f0f1babb0c033880cabc706b4f338f3b5fa2be27def9cb05239f7758be1cd87368e1bb6c29bd6841f8de4308c657b28550ee121c0d8b9d56daf29eee100b5a6ef4092fb704014e738d5cf0787aa68112aeb148;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb424bc76bcce9ea4efc368127bae724ad4cd604e1637a163f1034bc657264923bf4940509048cfdf374d01e2b7a372adb6c383641f709a89b6ed27f596e343f86d46e731c917f0c8633c11da28ff859acdff9a6dd3f83be8cb8faf1dee61ff55cf28d0a57190fb3505d0e39c6d264c725afb96a52b4094fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30059105167e440894011f9192ad6e54e5e71e3f86489bad6c1b980cd2a19698aaa3f8f27f10f2a6858c523c34aae74b7a75f6d658d0779397326b8a802850ae4c94c1b69e70c6f21cdcdbcd2afacc5f31530d329f3d2767c1713afc366f2aecad167cacb4fcae7930250855e43a0a65426949f4a6cde765;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10266b669713540e344c033b273c58e72d843659584c17b1084e0af39ffd1d60275718e67244b6308a1f85b43afe1e6a7e173fd301ab051d8f134957c454911cf337275f58b14c41bdc00c98a819b17cdf86b15bccd56f28afd1065e7c3e187bfc1e938c33e752306e45b7795ed9450823f9b45e4e647e729;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd111ce6fa53af859773576b4d1896f39e65d8390e3160acbfe8a3db7e0e4731d2cc0b4fb8568c81361e54257b761ac886f774570c0344d0912505c72ee05455dace02fedbd635f9131d6b9be83f087e1390bfaad979b831b2751e17e63cf6b1a6307c4268b6a2c4e8bdb1e950c87b28b3cfa20e3cd0b077;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf20ebf993938e1cc371798c3063ad15ce2013dc25fc0b6a01dd7a06e7294a4ed9c54fbf9e848cec534083a92a030a3a8f855cb771b7af3f6b34639d3fdc42b745a36e4957af6d2285f035934ed01b39e4453cd234198e5827000006455600fedd91f562666301c9dd3dccd00d8b492f49e4300b218dbb19a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7b3b45e87dddb33a5b043662b1caf98449559a8cbafd6466d22653a329321a4878e01f976715d6ced75cdf9e1525f2928ea50b1b87a6771218afbba81088281066314beb547cc720aed5a82d8d61499bbf563f4b51c55be9a1df65e47619c180449bbc9f4306bbe9ff456138d3d1803337d8773d6bb0eb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5ab48b3b27dcfe490908dbef557f862a7a23ec8c485646f6243e2bc5d4a57f3f59cfa7635b697cf5cd51e5a7c5fb65c75d825639994e0656d5693b1df50dc643d3a4c682bab4c6d8ac19cd4fd378ed869afdf6a7baa0d50bb9b13636ad7bf52e8c36daa908582520678761015ed7774ffe02c371e762eb12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147e42d3dd2891b30245f7836ad0d9ab492b09a53a1f0c8db2b59be3b23b734f4d449138399a9edb528a75f2f84234a3bf104ea790cb527ca3610845ac646d9ac240f17659cf081990c1d84d59c4969020d4f461781c10e075764be3d819e9458d9b7b25e70f0dc26d11c3c50cf1932d270923c6e0c8603ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8b700072fdd2ab557eccd3c7731f818da3045ec6fcdbe77975abbd50ed3654565c775c747e9ced9541b4ed9fd483f620a16617ef95dc459d143b2d7d066024d021b65b3e6bac03f9670d454f49e7ba23e4074cc5bd9527af3ae148ef4581e68d1d4033e7c14b3450a6ca0a1a2794ecbd7a72320d6e588cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5739f1ddff843449ae3f809cd088ee4130982b9682993235ba01c31efe78c3051c03444f613dab47ffaa2137c28a80f6491f5615a6e7e9252931b4b97aa01d11f1cc572635d55d025de78e199502eaf3f184f3a16de7c4b1733c48e7df5ee92c6a40f344d2ecac28b6e75354507802bcc02ba8b180b0ea99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58215e55b48089f50186f641e17f94facbd89a4b7c764568600cdaeedf52dc1c35a531ea62cc74834a742f3dc8fec156dbafa31adb76319236ecfef778ef22e93ec1137da067ee36582f1baf341138659180d4060c7f31b2c7fc919b02a0d027a43f706bc3ca21191540dd2c3c182288c9948526482f6ace;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10221d4724a80203609f68775568361baeee7833923a37dbe209f7eb650c55aa1c979f65e6227653f6eba1123df2d77b4e13d2fafa3847aa7417c2b21b5c6c6f6712ae0ebedc861fa392d991c44c04c8e87aa04e7894beb13ba374eebdac5bf75b66eae98738c2f11cf9a15e4764922cc661b7906e5ee2bcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8ec182c8c31940931de31545e497f988b705adbd2ddfde1ecc946a54d1d8ab9aeb4c8890fb72cedf6f3feb79252a8b283c0b3eb3e326e72ed5f8d98b4bc8d06000cba9272c8148ca88d67878d1af2de7303728b297819c526d8d36455fb6e7706bac881eb6c08035a0ec0bbe45a57816157f306daf3ce0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170ffe3c7ea3501e7bca4a5e596cf18e278d1d799673c7ccfed809674bf0bc6583cd36f7534ff4d8cc71f8f8cebac5834eb21067bb62beb8c5d0356d91b1fadf98f9ab4a539c36ec697bd31d0112bae41d2beb7f3fea649ada56c3dd5724ecfff1d75040bccb99ef8e3d77b48d017c90796e059bac927be56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5f15e8d31f27858408464c240428542afc5e8fc9968cfb29f64d4d674a337e6215336a5e6c8698f20355704a20058b1defb85a512deeb024bc792a4d4d711c0d984d8f5d58762b36bc211fb30fab96a4e35d1e72cb9ca06ca7e8b5b7a971fdd2d04f3a6a8ef25ca0bd22e475f7c00d44271004bf135cda5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d38f3ba80df30ca982c53a277fa0b01d7de9fd7b7a41084e34808976a70bf360161e2ebde7918486fc9acf897e9ec2377f346f14ea9452c1dad1003452252cac2b604c256e6caddc01930df106fbd498977774699da12136ae370d93bcb3629cac0f0ab3ee990e2ada9881e7e8efb6695e93963795eec94b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0350b6e6bfd6b21c34bc4fbf8dd8022412a92e674ba8e7d382825276fd19ca2f8c74ae150106fb583a33bedf3410c08d78b8b940e63434e008364bff44df819d2548a44dc3d28e59158dea1801720fafe487f2e7bc51bc406018d7c939053c11e95cb139bc27a83bf589fd09f0eb770a5fac0d4ab7e4f4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e6d9b5418c7e5fc6be5184046cd39cb4d9c403efee9f6f04a48d546dd739fe66439f0fb16c48481068b2dd534b526cfcb5ded9112124c91d2c202a8e34f4ba02ffec9c6ae0077d9b479c745231d0e714b2afced9aeb994dc4a85518681731ece362dc0e817a7bc05d9c0a5d5ffe4a837daf0de160d383ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe6c4583a973ab8893b7178d48298da91ee09b013b6c899ece7c0fd495dd4fa8e9806e0e62fe580a112442c1741d1f4307a3c84fe5f65dddf1af846c60ee5cc6866f24a12077987bccd3ebc4f80c4068ee4f525a58990059b4a97c2130db642e2d356f1354f137220f258e622fef6d60493787035990d0a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6bd90ecef7fa097debc521b5ff67663580b585452c70fcaeba4228cefb14d1483a26e95bc07e8e16262c3a26dc6817d5daf991840978ee4a563a50475eb0d39a7c25357d0a612d75be369efb78517b147a8a14310d89ee4bcc525514243e67aaab699a0db66eb51d852de4337ffe4174508165f68fbbdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a91b9737a5d909a9aa703a0ee95385bbe6eb7014e6182ef2346bccfb11a51134857b6a8122efe20d5b4f7633fdd5f02bc92e348a183dc770aebfad11d65c5317a895668448118cb5f876126b445674eccb1342045978032c0ee6c1d07a8855664e768706939a5e9a0a5ba5685b1dbe2704e07e510ddacc09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d46dee24f5d8785bd1d37df84599bcd71a2da5edd06a257e3b6f4090c7adf5e9476c073c1faea2bf3b828ccdca304ee38cca91391992500bdfffe7a1825ec2cfb1f475d475429c285eaa361c5a445576ac371734f5872a989570caa7d25d587903536d2701c3f50b9f7a862c9d08a9b699fe66fb769f64ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1587bf3ce090522b66925a73fa92bc2dbe3e03b9a38ff3d880c66d754a4fd1964d8967775b26bc19ef200b28cecb8bd96ea0d7204a112780c05c1f83f9c6ef157e8942505a032633e754c910811cf5aece24881d4addc31a9ae734a85243742c3d8cfeb186c99c9af7d468f0aababca8a0ba77acd6af02003;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8dfd4d67b67fb7ce89419166da8328a1514566224ef71ab15f7b072d76acb6cbbd8bea14b96b2c290682504714560c0f460daa21e34d42091ccc3697d557e21a8cad01a1d3c8c5d7bda4b652a5dbe877e2a6d8bbf393341de764f50b75284c10d63c194ef8c11d669847dc891912f4c9569674ecc5cfbf8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf16d32ee66ae82e204ae3e521960e590c0714a13290f77e64f413ba9bc69ce5ffd84646f75b25c9f47d40286d3e1db46752ed748e5329f60faebd746d2ddac47fce8c2a47ea5c389cc4b8db37cb1a1d65e6f1985f1d40ff44e25bdd2c277756ddf8d99e79eba01387de97df202213e99d3d9e6153d98bc74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a64d0b1bb6cc2cf4529de5ae5243a658953187d30aaedc1dc434706b8202220f0ec455da97216084418f8c9140f17d8f7e916ca7b131b7fef1550c1772d74411ffdd89fe1dfb186f171f74e4618615eb17ba2ce036d4eda9633756c3b59ee26d672cd86b44ca4c29ed730176195e0e1906ac8cfe094ad24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14191e0ad2eb995dac23c84ffa3d2f9ab4c31b8c696070372a46b1fe92e0f3f98bc92abd34128aaa1f38355935cdae1810752b2981be9ee35618c4a914b4766bd44541e050f322f99dcdfbfac58b2c8bbf05be5e8b9bfe93a823c787198d1a7f5c71e18601214a88ae6307fa8a2fecc9210559872a0467206;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c031469f5df5374f7eddfd9cf7576c572f34d984f9844caa61f15fb6dee0b70a88db8cca744f99ef2fb96466c54fde686b0c17efce7740e99c811deb6e396b570e57bb0e66b0e6c4069ceeaf124aad974e482c39dcaae6cdf51d7c5a2e30eb623c113865770532641edf8d72b8d0ae5108170600a767511e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14097b0c38b1cda46db493f15c4c295c86c451f3c3f9e752694e5573c1839492a426f2b97efd43218d7a8802caa24a061e8158939a10788c280b01ec4cd337ea620fbc0cd18c52a709ca97c6c6be1a1c142eee15de805af7001636e66665e8891a4fc26879c94cf977f92ad77fa5153a4d4def76dc51d62d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b248bd8654156a6b89fe0998f95462fc9cd498f275cd576bc3479d27e207a61d15ef4acf78b858e850d0a0b34c6ca6f0c18c69f7049392abda06f3c5e9b5fe112a5aaf4d47a01f2cc45da2d88dd6d9782d478e673fa9bac6db33a5dc7bc3d108c6180148396daf09d55cf279bf1649de008fb07ed93b630f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7715fac6325583dfe8201413492c2766d84f37fc8c4849a89cf0363dbe3d353731fd36a78a2c6350acaa3c1be540d14b56f599cc632438e5cd7c1cd9bc322a0f46041c6768077d4a8121ba9abf136502a5722ad7d462474331bd8439575abc41f752728c9b78967f993606ec7ce5bb50be4697bab61395fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h371065666a048f83e306616abf05d299b59d5f173d80230e7bee5eeb41aa7e5ea5d87abe58093bec76ff28bcba2d263defe7b3395af44929041981377437f8cf50d42966676b39d0b33b3dd2f1ac324136c87c2c3c8432065e0dcc5712500c111ec33a765a8992194452e409e0847f8e961061cebd99d20c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0f5d62a825b224d043e36c8cdedd154b016f06cdf73bdcc0a89cdfb7c228e5669f246cdf074fee169792c06b3989171fa6fe0c04b96e777dd6ef116f3ab7c4ad75e2a3ee3d4e799d0b921c83bfb765d14f4a291746681b37af8b8f153b4dabfe6c41249306adf11bb01804e68d0ab8996bab090bd6e5ce8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56334d8e8528bac3745e2dc10cd8dfc7aa93e85091c69d906410864541d6f60daaa0ffae6274c0f9431520ec8710ce1f96df9b12dd88b1519ff774920e24fdc04b4c6845a65914b0f1f61e9484e4e52f90d3217a69e3bde5d8d0bda56d15e0e82ec2491af04de101ab619afe201aa4e5d248641e49e65a96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb191380d1527eea4830231075c6c9b2f8b306c788a083da8305caabae5edec8b9d9af4d8e7b3a67cb74d234aad64d980375fd33bd39976b6ac47b715fe40a66fc7030f89a67ce4cc9a52146459f48777c1f2fca148fe8bc1e57c8333c55f75f024bfd6bff901f4f707fbf663eefd160cc15cb185ac5c244;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80fcee5438cb2f86a8c9a0315e3dfd4332f53c0a40adb10e7a412a1d00a16e1cf7ed81fa4a12b64e78fa0b20615695776741df87d5bcce87107177e56a47538fe736a2cd2e2f887ba50dda50e37e857cd1bcca029ec58ff1b3a0d5a47153ef773e3ba80f296504d9b1488919fd53a1cb5cddba8c672885de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34c68528de2231efc6c1713a0c4faa2620b655d378f31b0001da8f1d4f492580eb9cdceeab0f96dd125f8e95c292ac3e48fd242898e65668e297790eea8fc064eb93a97fc04eb48dfa02e254605fe6c40aa8eb513c5086bb0fb2e4c824ba9c87e47b3f3c5383ace4b5c60c09d95c0d209fa76938b5676083;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82406543a89dcb866984fc02c475d5ea839812c281a1be078cc56745ad84e90e84eb4ba39e54ebdf35605345b9a482bfa74245661d2adbaddd3792ec4677ad2d324cdba3419a8b355200310ed1755a059813fdef5b312b442e08ed803d55bb99fddc9638143f496309a684c20bc5ba37127d2eee51d07fec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f6c49ad14876e72a1a01912c151e0b1e0ecf8a7bab34f1611127f8d52394eca4bf48456c84c44324384393ae6dd77229a015e2ee124bf70bc1fc4d2a656f0d7a6151e1f3729475d27e8fc0a34ebdd2d48fa87fa385e8bc908e5382b3ac0c4f1a0f633d15fcc3b3346eb2320c424bfc073ae17efef045f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b1e2a500556f9eef1ed1f920339b630d7af91178d03e2211135ca93f42302d6abefd36a723269be8bf2657ec136cae1b52c1ae93197f121c63e7576b8663905785db7f2aa0a5aa14177c0acb4d784c0a4599cf29141d29af5aaff587bc0f3d23f5b629aaeb20f4de81e52e913e53711623b6dfd991207a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab2260be6fb186c9722322acf894b19db8611aeba977f0ecb89d347ec9c2bdf0efa2ea5f7c0cf429ff0bbc5bcaadf97190bb835528b67ca216c176eb3b38997a139e5b43eab3ea9d504132a57351db12c839389bc50c96147a6a0dbab20ca773cd59223269796f5a483a3d2a98b9e534821564ebcc23b029;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190f08bf951ac24c53d6dfd074e9178dbdebd24d0e593b072ff20470602dd892ff0bad1b06673deea399eef6d41b4b4a4857db35aef143ad5e43763f0de0f7b565e3ad49d02f393eb91b76849927eab74271f982ee1801bed9a829506c2e2bffc95ce8e3715b231198e4979879bceed6fd33f690235409122;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77d5fb4f53468bb151b34ebb448f6633a5ff10b62d8901879d383f23030b63c2c65ebaf667c6cf27c0df5cb0dde741a4b3f3f02533c9428eaba98fe70d1fc06478c8f21ef99c7077bf5b968e46a1b737c93c9189652632fcb20930cbd8168c5aeec681ffeb0a095bca02ca7baec86838189ddfe20f0ef1d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f2c52329ec05885563440a8f9dcf8c7e1ad0be32e1d6898a060603c22129d9ff6f9f7eb46d05f4c0b3d4ed6fbe9551abd5f00ea0dde6d1faebccc976c654084890d85508131dd716aaeb386e7413c219cb9a0778772d214db0c3117147e1fa434ea04023488b62a653c06c253689298ac371c0700a0ce7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c80535fb46d5fa0b217318568f1270b4184116f06b00f6677b6a2914d5059a409db9c0425ace7cfb36b17385352f932f32dc2a418f7d14699c905c1d94c6c2b1cd1f5f416bcd84288406220e82bb664ed6fd74fb9f50bc72d788db58dbe4143ef36789cd06bdf72e35a73629a3a32c0c2cb514013276c64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2db4aede646931a8c5def5e058ef9948d197e9de1d68201428808b15bf0ff55421f8964ae95d024a9fae7d32a969279ea03a2db1f83f91fa3b242115bfff82f967736aa28d45a691027f8f63bb14e796b18f559a3f2771738b754fc6f7ea216f3b76f38ff0a508c4dca1ee1638f9a63719720f82fed09df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d41adf969f8baf69b4698bf423c4844ef4a8d9e4af79a87a33f544ddff2e6f5b11a9b36dffa00c4d3922e6a210ef7cf8ef59e59cb57837075e0946c4f03edea03e61ca396a7e22479d3583a41e07d3bf1af940becdad576c2bb4b91db4ceda9601aad5be329ece8f02a69c8a4f97819ae374ca76ede2e02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109136a261f92294a737d3a76197ad0db242c8758b348e193662badc9e9025219cdff3858e62aa9acb688506e037d86f4a6dd1242859711dad49649df5370a92c39a4dc2fdf848a4118cd0656189451f8bfa5ef0f622d80f0b6ab4caa1ecdec6835af15c69a1b15398f7bee57572d5ef911629c9c9d91d5b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1301452d9ef9b4faeaf971548a25a9f92a0c7493c00876dd5a496288c95fabfe661364e61f6e15ba2cfc4070ff225d8d42e35cd9e2133a8af6d9b9a7fe1ab0e45d78bded9a67fa5feba401dd4d07a366276dba8ae245677cf557efecd80aa68814996a2cab0de669d0390ed74cae237cf0c667df00a7c09a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75d3c3450d7ae35c7dfa6a1717272a814f1e26c3fc5ed3ddfc70cb11deb67a0f4465dbaef09988c4ca0f0e2369660175ab8fdb22240aac1374cb06edbc7abef7f9616f05f13bba5d6eca934950db4bd586be5cbf22e314d4cebf7cf9cfe59150f08f4359f072290699baa8a8d230b3b0ebb8c63d2e849b2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3e93900d01568e0d07001c10ce0cecc84c91da7fdee8c3fdff4542d8a3a701aea2602e49cda0eb079a7d0a04a2d2c03740e0e58eaa63ae4b60ef547c9cbc2116e17137c559d3b4591a38f1074521c11b26d01ed16e1661574930c254d3f4252950ef002ca565a8b3b04e5f10156b4112c96bfc2f3ef4b3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18bf1efbbfc70ca58f2a4c1a126f25f4b02485cedbae60a434460ff0831111e6fc5b75947baa2e1d494480343c1f38facbfb5ea181a57d10f8bee900cd867fc77ba5fab98d2048ce46caa8ada399e263f80c77761046fdcc41f5405f12fa4a1306d43185e7f3b92b9905300c4813f9b577b5d8d8a0b895571;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146980e8492e69314ac180c0d72630517967f560f34a71e1d6a6019ffa87e23f27258bebf05447919ec71b4838a72912b0668199bebce348a94fc84812e4c0a6ac2794f6dc14e6067f10ab189ff5ea032d65c06aa6b217651fda03f0d447cbc6d24527a9cff7f0a3bc9768385f4383f1a3a34a7d6450486bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12474385cb978dc7205765b7d6e212eb3891b0b022cc913e84431471eaf09b263917af441b53dd666659e8e2f169b00843d6342413d602153c34913d2e35dd865c7110c7b68065b6fdc3d0e3ba2f9e11b2de1a4c8d15ba6c00353bd5aa0b2e8b1b32342c555d4489a9ee342715a68c0886d284dcff5be5025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121e9b0eac81fe5d942115a5ad7efd7f3c52ef1d86e2214998fde926a9d17bb07f145b3c6e3f4b5ff1676e1294f03fa72969df19324f98a072230c97bb3b67be2cbdab3823341a9333dfe5bc2aa891d22339e7b47dd88c0cc2950e579a9c273b8498ce902a6c540f67016f50e4aec948d8b0855101af3f458;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h314303b6e09a3c6fda08ce6093270fe401655dad65924f541c814bcadea858479e7358bbd40bfeed0657ae475345cdc463e8cfd2710b8e4609c5693333addce88e984af91c559fcd57312311aa9d285e9bb8d7a002be8d6fa565b4bb3d8e05fa8c33971a363e3c188b9573fb7bd2aec2d41ab3f0658858ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8dc437da80e2f74991ed696abd3bb439089d2730dee87cd7bc68f5f7bf9edc12a0333273e360fcef8a420e24254ea38b8e35916058334c7c762d0f94e47375fd7d761eeb53e53cac29004aee8cb05b9e351af1a2da2e6cacb7c571990e2ad862eed9f229cc4022b1aaeafa164d60e07503f192cf2a0aeb6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71cb7b159639120e7ed55cfe7cceb21eff8614e1d7585cadbf044b49bef20bc7df40ff7fd8a6606ff02c55f7fe4859240c46a1621869c39965352933de6ac09f1e17a85fcc1fcb8bef82996cfbdea0e4d87f96f12a6db4fccd51bf255028d747e45f2ab9e32086090835d142d5e71b732039f5bb451ea9bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116ed9c6b1ebdf5ab07ec57bbbf57a8641f59b5599b2bada6d8cf9d3a6d786c809edfabf16dcaa7e5067e3227847e0e4b41f748a8faf82f8ce89f19af17e2a8679058ac8b410ed68937a03b64e72d8666436130cc50a76ec084193d7f6326c64669c8518d23071e6706e5b23519f8cbfba453f840e3c0713b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10264eec5c2e686cb4f4079115c1f7c8a251ae269ffbc02a3e9dfd2f761aca68c9b411c77efbf60d6de142e08cd6a40aa8809188a7a42bec9f0a8397e7e22987b3c95934f0e5f9fbd74b77bb5527a54cfed4591a907ea61e5169cc0a005b17119803f42b0992483edb2412068d2868fd61b31cd7cc095f22d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f10a98300d02e73a1a91cf723039ac20fc9e9d432f42dbf062d01cf6c3393e46c4bbdf5fee663fe4999af9b132caaa34ff5bc72ca90c01f8a578a598e3e4b4a53f7d259f7ea3acbf31109109fefa5b4b949d598be5c9bc126ce22390d2c933ad5a7ac2e1d02cce9d933cdd2ace3d86db1df4e0b55b164e9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1818a1638c0c8b372b718e25b384cb2ae2487e7e4ddd568e968c63f4b614c147a08a89cef20a761ead1e556d8438fe20fbdeadcdffe1fca5757c8efb761b3641984d9b057441b0aa91dbd5bb813acecf5c00c00b7a1eca9cc207eda183c4a1b0b1fe89c6ddf433c7af27da1485f64cb084771cc5369586739;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173143b3a7f26fc1845db6069e7d6b7bf6a41972448275c7ee90fec0ada783cf09b8d028852670bd870c9c9be15cc7d5b22a48dcec31ad4c4ffb96653cb5b0a91aca507d4d5364bf6e747a6eaa2ed86fdf280685568beda5c87e039efe0219d7557196b3796b2a6b288b82d1f414e33f6bebe35e85fcf39a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c78c969293713067b0cac924def659b0ffec1d38871f6a2b29fcc1d5a522e51758eb8d34eca403ca732d07a276c3dc12af4501e7a4cd06bcd8798cf823cc224ec245dada4f387cd9c0589f36079455f205a538459569a3dfca6d4334a38150b237a9a65fdd0ffa8e2d0e09e83a25bf257d4cc95f8fe8493;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9acf415763f35240f8f304a0ac489b35f3e05ad233b5d6b77ce0a1eec536ee0c1e383ebf0db055516a2fe46d1cdaa853d135f1d5d01944089fa8254e7ced72dc9db0795d7476fccee838fe6ce0ef108dc7472f8f771b1f35abcfe480498929b99e4855f3d54893e4cff11dfbc5b46b2efa248445ab30085b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c733b848d7b318e3693166b0fd4ede8b9aa9fa2c1f4a6b91641be350586409935893ae4649169503f055c681f7426645a727594372c64d92994fcb847adafb10e2fa5ad8e71e1a9b142019e5a448c23f6a53c2d5dc3b8aba528103cf7f113b99cfb9997a19e299cc463528a96be949af3b36f1643c47024a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37a67709b8ded89fde1864c4c7ca3ff8feb25c2587a5eca44fe8fd64d23322de6f5069f859daa385c6fd97ced764c3d2067605270772d7bf378bfcdb9b024eef2dd53c8a64b2256ee4a7e78f58c852d3a83e4b280f989defbf7124737100b90700d778ec36cd12854293c5458b801140fcf5d7878e6fcc56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2a018115e7630340235fa9292779739a915cb37852056f379cc8e2d5d70ec0300872fc9972637458b9f5af663dbebc45f17ffe4858545dd8ed590bd427434bac7f90c4b597958907ee63407960ffeb716ec5d45004e817820eb33dc4a6d5167a51f6fab068d2df8b2ea5991a8c92355d2a099fb87ef9a72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9f8e789333d63133b07e733bd9f9b935f11331155b9ed40a4f014acf8b6ab22f052609528c8802c848a8a9c4ecfb7f63a7a6e99c929c6191f7d8d98bab6b0c7179c326f9e27c26f1ea0578d7037494d2f2012739506257fc453c6f43904b3d23ec22d14cfd10d071ae0715d1d348652ecdb855750928f96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7480b1d98b5dc378c7f0b20b152dafbe44a13aeb5d8f75d928007de0e958d24886d7ffff50f1b9c07d9de175c6573a342600a246dbcb9298af8b35e68a7ad8673ed3826140ef60df98370086e33bfde90cf50ae16105e467d8588790a1cb16161a21249d84b6c2a674a28163028cd6e837dced670026c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc61521cb945ecbd5cfc79dbcf0eed81232e739ba19142aefe0f3e900327530bf1b70a8dec0e0a9f22047e95df525c6d8817389e4ad39ac8c2a3a01597779638eb8ce73af4fe13ecec489f158904120366c2cb4ce68c62dadf60bb0719f1234c74cfcc6a330a257a9b9f8b399f277dc289e5c6bb2e21e094;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4044cadd7125e41f698d95bf2c2a0eb632e5cac8fbee2af56c2b107134fcba6190229dffe3829b9e603e3625766e0f713fcb03a98d310eead859473ba3c486e286081ca021fcee0a115b10ff88eb74e3a74bc14f673b67ee1f8069d6995bbfc5090cfee3e1a41f000ac71da2260a9facb682e4054f76d1ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a25d17ad1c89b589a81a526798c30a805a8eac1f53e6e22a5c5cab9387dd00a67798021ebabc793c31216173b63904e68040c5a878f655b8090dc21ebc5112c477b4c5d63fb779e641c04da67b782b9a7f334bad1fe3280e02fc1f8681e30fff9ba83064ae5ef45bf2953d2cfb7e2d0f6711ac2213fa45ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc3ee5bd11deec82943ee950e764b16004a938ed1143676d4831026c22c8fb72490d351d7251bf0e7d16d573ca43d9d394897de33179e9a5be963397c037cbb19b338882b6f4d5277871cb5b4991ce5de37efbba0abd17ddd4c7edd3e08ff329eb3568872dd609e1aae2faca96f9c50be3e057bdac552a22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11164a8986ce724d18159d70a09a77aab9fcb25fd570533f8efd4da13c13ac96b15e6057e7cdc3d9122d8dd3d7ec872791a8e3e177ae85d0367d2e0940c4c64a6a21ca2aef7fdc8765937053a0ab0026da11a8de78638e0513f4dae558c4c456c59c6d7ff22614f116dee286caca180c0324e64da5d501de7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a88bf5f2aeb777aaefbfa97395a2788763b4e64aa82cf3c0c865e843f93d68991471c849d771576d25abc9fbbb789887f5f72f64afc5415268be0c79fcc312b266adbafb5b587f19bea917d1486f0af67deb2336193bf040b08196ea8ff73f339c7a1688a7fe99a1e609212ba401bb65730c80a03e9c09b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28a258c63169bb6ac470bf718a078a17e56d9ba00fa421664e1cf8a74fce97a07331d5ad8863f5e5a6c1b5c728a50be55446ae2f7b52536aa9000d370cfd2075ec2d70ef4166abc912bfff34a6cc955112d5172d64c8cf06e78c6bb71bcc545eec1d87724b128d9f107eb4b1cd015d4dfac21bd9caf6313e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2cc6b699ee7b927d94399472ecdc4fb22a62a65cffacbd2b731ead355f29a16159e2c0906b37ea9051d60a50a6e93d393c9f3048cae4f89140e4f9b9e14ac111440da1be688e37e633732855c6213803c75dd4cd73022a658e7a90bd32ece0bd0184f282c515d6712b2590fcee505fe4bebf8482ab1b45a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd7423b53e06c835ba73e7c0b94eda741134dbf05a5b5b9e9cf62c110863b2e04481b74d0f71651d8a6ecf7dfa91ec490cf9f334583d3ad0acd8ccd8023aa5f3728a71b9811aa939467039c3766c527e5d1c88c4d7c6950738cccbe8f2a5025b2aa2b41dd77a4df43872f5c8f52826e6f73003d29213819c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h990c432456597032aa5d36be9c65f10476a51f3970ff939c02ef40fe9130a5766afb76768bddcfba00692e675005817ca46cdc3cc4f8c39138465e42765950dda09b1ed7ecc52fb5b21228622a4151e20be86cf54153d5083a10626373f0f2c8cb9014f5a1075c424d8a4ace133e25f3b507919aef7534a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecf3ea5bb6d78fbd6876f101a185563a120d47ef1b7870932f7693d7ad47d3dbd7294e37e9547718fdb9da9e7e487d663ee9b56f8377bb588ac4a7918ac5a747297ef0d72cbda9eea5c4f2e227d62478305c7b24b6f50b45442f0e6d25b8c5eafc9d6b744e37c8978a216691f984fd719cbf6d010cc6b6b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27758651a95efcb6c1a6caae0fd8c2da835e561b5fe2e47f94d4247081f76599fa30d2ced349ef81a887d214fd65d9ac9842206b62e75203b6c3594178e713ef14ab7fd96909a37e14c6b7b37e3a13f8824f0c9384b925c387cedc00088847ce4ac0ceeb46601e0327a1897792a88b6e5330482b16e4f2f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70d84fe7b7cb3b90d9f9c156897fe17c703ba898b58f88f79043bb949e1ac50513e1cdd28f9e36bc3012c5f5386238d832c1317e1e4f53de025d2583cd9fb10f1531a24f958c867045adf64638183300178dee49bd7245e051ef20f283ae197dd87f6e8f7a2d8e49d43336da5d8a180f082f4b0d483d55b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1231f316a6f9b4c6520756da8663eed5c9845dfb722b7bd1799ef84378ece9724bc6fa02a102fcf9b9c255e188e1c4883055b4f35a997c320ea15fcc5a5082045e07857e7e8413e913201c410bf3fb1cc96e2bac9fa69fabe16da6d4b95e81ce1ba1862bafa2171d9268a372261d34fcf2518ac5a927c1c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be33e48c2add4de3b73e2da3b4dae1146bc43d0632c4cc014e435cf179138054aa78340def8ecd17f6d0ce29f28ca3214fde2c5d1a8963cae6a1f23047be48c705294cf6d839d3318a8c800904a5a7ea901bdc7a7dc9334dd31169e39295f8da68528a9ab29b2b5629899156c09da033400409e9536aa583;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f1556e07eb6cb3b11c7ef99b34fe908ee3efd8287b897145db5c0195f19aae1602e44b7655a2f8b8d45a6232f509b61204193a31921c3d1f8125cb872a4b4ff248df9718f6069d3cc19491d3c118b74162a531c869506f92a7bd5098e161b938817f5471fd856045d47a1b8d5a7bdcc5dc57cca0e955a80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf5a9536c8ba74b034798a3086eddffdf4a7fcd5ca65c30d2b1bc2cc7152651a0024fed9c53412975b4599f99b4e4c4814660e312b1a738de3fb2ee29d3d39afe319a5fb00044855dcb6411986cad09b790cc7726051cb3fd968500034c80195354db5e3e006b46ada7cafcb4f4d3d0b9b8b34794f92c0e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h290c08153ce9884c10652b347b22937958b2ab5dc50cf49b401a3e4deeb1f821dc70b1195169a28663ca7e98b383bbed59b05f270ca803a75ee86bb56e8d7017c62a190629c377a888c2888b3fb1829f72c0c55846acb33fbd779e51d031c74cb63b65fb1fccb62ef8c2316d11259c3a909716dba78c9c4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5191f9054257093cd0fdde64f4b854dac09568ba73f19e75c5f3987521943b54f19a430cdb821651c974f62493c345f5766ea8498c3c42ab55ca27bd55634ca74ca8d97c6b164611b1d3e495800dc3c0575ed04d2fb5ee0b6b9fd03e10a8b7640f176fdab6001bff4cb1f790a586702de346c23f077605f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c03fffb4e5c8edbdbd9db5a12e23165645eeb7746d3306b0a0ee9d7cb67a0b7e8e7bc3b3351d031bee2a06f477cc88345578db8b14b72b85f3f96002bfe72325d79f0b82f16ff5535b5720d513f24292108ecfc9b5cfca11bd1e6f7c6ee07f03fe8aef7e7763016251d29313b7d3ff21813e44ed415563f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f1b2a5fcfa811eb2575408e9a43dbd0266ba03d26303b15d163c173d3fbd175f122f0fca368a23beb4c0cb5f3ed051e4e06be185293a6398af78f5d4f199b7d99e1e857945b9f4a2888ae7a241ec0d2f2597156c805c7490a243b87cc8e2229539eb79e3a63a73cbdabb30003c9a5fb78458462c03d154c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec6e98aa25cdcb1f78be3ca41a764879d6bd1778410c3ea6e7758ce0e589ded86a0b20c276ff95d929b382e7dfb7db6da38c2b913db50acc8f4d946b3ffcb254e3bd976c96fb98585dbb727a93ba8d38d523baac9907e19add021c6e26ab1bdf284ce10ae31c448138c38c2d6ab021f5ebdc2f8d180237a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14246951e44921a08857d23cb5e2854b2d9d87adc94c806ea72b4a8f8c775744bbcd581fb2db1731cc52590b3a5dc20ce7575d17e93b04852a7a16d492352a7ce0f024cc82decff86fec1c2afcdcdd543494deccd3c9726e25e5f574e902775790e787a884e8955429be233a2acd88dac1e2cac47ec1b80db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a89edf0c4035854cac3cc41d722636858313f5d5d79fc76127e3d8207433fb6631c4fe8d385814323eac7269f5aa2c53ef863c5e38ed9d70b855996e37a5057a328721e88dfcdbf6e03ef813457f92d918881f2858f2b2d2d4c8bea98fd06209c9432e9b898f717a48b5ca5dcb43d4935d2bb840dcf7cd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdac1f42e3afd9009996a58cd8657fb91635eeb2596e289fc049d95482cb5b4a011fb6932baab4983a6c971a0b7accd3bdbf5e2c6911d999e371da45d72cbc39f09cec9115fb76af5ff6b52b8cef92268c865b4bb2b03dddbc971d8c609fa549e307ebf26e6eb25eb90f9d8850f9b04e501ab3aa7513b8f7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1bea771a84602d494a4ccd1b583728538cbc4a82ed37c33be87b1d8fde4970acd090a3e90056d82500bc2860746218bfd81021f424322c78b1a555598ce68c5ae8cdb32d0765fff1f2d204fff31f22ac476eedb78e4e5ce063465ad76ee31dcbe5be0bb224d8b715ec53ba4dc8139bd2a84d9ed1ab3c6c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he27131440a125e75eda0c8b113853e0da4a2f5711fca5b0b7bc69b262ded4ec83bd75e2745399cab273d6bcc47cd6aca6495e451b48861e9a01b2d22df6857af48ef8a71030ec2b15309933e4a1f43692bd72fa107547ba20c910e240f99c82f631206e98701901af3e355d0599b3ba6031069ad11b9b44a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe66ac1c6c0708508e551404ba551b4495597d61e5d2001b5f9a3ec1e3a2807bd0d95ccfdce1725bcb5ff9cb6198cf5955933e35e35aa45cdc736314ec1261f4cdb7a9953fb160784fa05249a8c86ca09533a148e669f14f0ccaee483e4fe286d0c95f0e834de07bcc7fc3b951ff7f2e268947b9fa855b05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c143a750a463d9b802f1f2ce558c5ff51d6600cf7e1c90dc46230750940f9bb9a8ead0708e60548bbc7812871de2bfe935e848c348fe81560fc68e12e0fdbcd52b3a8d7eaa111f2f9c6204561d83c1c573b4719958dcd001a9345aa37482d7061bbfcf12e88a5d6e9a12f5589fcdedb0a0f4a7f2940b6336;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113c5f81ab91a1f6bc1dbb54e50e39dfee06a9077848170bd25d1d8cff5e5580402f4afa9db84193d4e592016c23e307725ca3975ca6c708527cd95b8472a1e746da3a318d0b08e7e09ed48fce5bc32901ae236bc5e1345ac177fb46cb2a275fed5ce932ab81076e3b0f6d40276ce475af4678625c19c8f24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64da02aa8118cecbb0aa7f573c8492f447fb02d156389fe2a798ca4395cef1e876fd53e15bd31f95f7c6fb65c4ac7872113280c9008a9a377173edaaf9511ccca168ac9af9d106036e4c47cb9a961410ac077cb63601323b94453ea7d31be096fc05c131bee6537ac7d86e303c1a7240f1c5488e9a5afbe3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h225808b15fa3447c9ba1d6c22edd20e3bb6430c5260a0b1b6a2b5dc101357e15ecf9acdf12421f3b7cc951a6c9db4d7f3876f5728b4c8d8e42f809b8550d2261747dccd2c0f5e59e00def9010050ecee5890e52d61eed5265158b24de67c2e0882cb73b2539f4bca6b6a17b189b3ef2187e31bb48e4be0a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hded952571d7bc920a02a094744cd9f3c890ddeebb352949caf569cecb0122d2a68fbe936370ee9f9f3edbe2178d89c262fa19d4426139df6f6a63edd13fde6dd4a2a965d770e52c72c02bccaecb556b9581a5a223126e6bba9f1864c275f5d7ccda8f98970fdba4e57f11f2fb6ad5d3980865063f09979a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2516a888427fa6d4a9a474d8894da18f71266c4e68c05b396fae8bf7ce1dc5e3c250d12a3fb3899df551c0e4bf3eac4fc389db0ff2ed4506dba0f4095803381a7bbfb80b3b879816058b3400c98dd00e85252b0e928d4417598a3ff4c5b6a00cabc0ff465633a28c001e2bc3ab9f00f1029802dd2d8094d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7312b22aac42d1c29103bd909280bb9bc87f7ed7b63a2926c7ef0c9e3a30c8f5bf9d048be4b3038351e96000e178ad57db814e8320af2c7aa1dc6c78cb66668ca6044c30f58e6d8edf800cf5489b15b47e569546ac12df8cff8371d98768fa05e4b7cc268813f4af1bc11c72efc462454e98a095b8a918e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf3cf9d8366604bcf250241807ffaccfb3b1107c04fdfbb4be7a119a253237df32da830f07cfc7d238e69c22f00f666b934c2783d2b7fbefc137ae144113d742fe4f755413abad0a4665ce0466e3a30d3e820873b8cc3a5fea8b208fa772924eda39fa25adf04ed65c2502111e41bf950d311bf5a72d2421;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1431ba1e7541aec50e4b70c4747987e991019e8d828160aa90ef6846fe37b7f8ee4c28719d870a8cf2f7a382bea46999f83d4c0eac7402fd1f2897bc1162c4f7783578ed318dd9b2f8f2dfe7b12c0755138b4e02e181c6b1e97ba20e2e8a0be0f0e04cce214f38fe24b8affe3d54282800f9819de43f0b3fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ecdd06a0f90fea5e2eadd26098ecf46fa74617c7fe6eebeb9f1f28f638ae504401d2a702706113ae94d0d120bf85cb890c1c936a44e6d34e6662b07fb04f380cd081c95ddd322040adbdc9516b13cd316b8918a3e525fa90f07a29e7408ced21b4fbed467e4bc3ebe78370c7ae50d5bf7fb6e14fc93d81a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108386d45266090e2e03933a5a516fd0f3ff70518b1aab3ecf2e6a7ccdc03cadfceed5befe6a2596da315f5f7cdf7502e47a2ea013c8c3771b11444a616f7983a5ebf8640622fdf7072f15a40ca333fa24276db1447486549c3ba62d90040c4d786f5bdffc4d6ef5e767cffe038eb975446cc161a5b9b236f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h750baca2c6337f60004b2c0802423cae152c26a27d0fccb268a861a505b8b785a99d241e3e7c5655cf7e98e717bd6e8ac294e53a7b28d950be777b0ea7c86bd38cfea954782e6d24871c1945bb2f193190c3ab94f203c9f1503457ae9ae9d9691070cc60e70c4dade4d3c5a8706727daa3d3120a4d5220ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35d9ebe3140400496d315b815c20258f4ec340e547f97587a36cfd8d4a6be855531b8f4c9663d2d7e6da9ffd74fa4b02317736dd5498f10a6e147647b02c651c662ead97d15ca6fad61a63e49f651d10b5d483aae2ec3ca3e257f88e133dc5418884df24433616882080b1bc88632122a9de3726652930f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd04f67cc705f072664a914bb5c6b784fac76a380ad7973281daacb82d7c9512a0a19360358fc5e1de7482617ac1f6db2c6d05ee7e340a986d9a565eac2761ec038a46e5ef82545923501b66c9b14c497baa47a58533ceb2eed39445593f3e691e3ae0e05510e1b68ace1a46564b564f6bf8e632e713e1360;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h434abe7f15d4b33f52740a548c558545dfbc188514226dfca3008926ce1a390c939002080f4232c1d42c4cb2db3112371146450c620512a7e54680c5821585baaa9ef2ad88ad6e9633f18ea67fa3fcfdd6dd583fd89abad095a130931dd346c817409d1427385d66beff61edc98933f3bfc38e15294110e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8213db3d1b04700b91459a182524050a4d49c8849156cfa643b53757415cc7d5fc305629d42716408a8d3ff2b7333bfc197803d3b6dc5ed6fde469d61af5362781b271637023a42ffcdd88544e6e5d3334499e0a2996167de3a513b8e2fa46003598dae33ac92447761faf81e3cb7dcc5168900463af90cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6bf4128076b70eefabfcc78ae94a9750045d509c92b58742a8ef85b1573963cf631e00691ee24d50ca7218ee05a552c49b1d7217b97889d0da83c087803544854e62aba3d78e976b164c3d87490a2ad9baa161f6fa88c5b4bba72a36453be2453039294c12c6154a71a3c84e4052392d97c60ef157b25c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1817103f1cef17550c58792e3e2021a85faabba0bcc76aacdcc139d9fbbfbf6375368a60d7a6addf3244105181670283ccf4b5317e42d88161bdc2e9ba6be6ac020554918d4992301f4859dd265dd4fd074b0b656d83794ad6b049043a52bb27aedb0aba225968c7671f613e2c7e9425d3ee33993a13126bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haecd160de7c1f864eb1f4c53a0d4ba8cb39baf99ebfe0bb7281f85670992bb53f2f076c49d3526e5a6ead1a8f8f1b6a9d5fd039f85fff9e53fdc5fcb02d93f0eba98fd968881460a525baeac9f663936c34acffed493a055f84cd20c986af65f26d987ed359d77587ece89327632162ca5404d2deee081f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195ee0de99fbd054372b3acf99cd62ceb02a27ef622182a98f255065052a694412782399f68ae599bd99bc2126e7fa7f57571c59318b65cc402587981cf4ef1b9bb3534815b8919183f3b3aa81b87546124d760ee765e90ce2362133c33cc3e98cdbcb9440605997c9a2f414c02b7fc7ddd7c207e20f522c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175f279705f6504da509130f65eb6cd3a5777c24942869de9e33165bc250f2e2b9deaccfb3bda6fe1aad20a7dc60cd4a85c3660aa8532c5627cfa5bc57984e892d900ffcd15db4c51fcb11a3ec1a1b48434a791d4613d8875cb8d4e237c5cf3fad396e30d4aeab29eb0caa86f1beb7b089d04ff126aa45f79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e656d301c8907db04bf2903629f8aed1f9852275dc06fc66301583649090ac36b6c9fcc67a69ebd5f19b3bc4996c81ba5ea8fdfc1c0cab2074629ef6fd61c3b88750d0c5a2a566c9cc974731e70606e2a6d6d40cbaf5ebd954945f4aca2d979ffd454dc385df98bda1146414c5abb117b18d2489b42f2de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d2eac635e55ccd2736bbc83450400dcf51ea1cf03b729fabcdea8022f339d91ed65ae2a0122bbcc08e320ba16a2316503a637a391e5a72750f3d55578d9e247085c2ff6b2467604c9eb0aa1acbeee76e7a7411d9c0578bb640003a013044748704434c6a7eeacbce93eb95ebb1f512d7f85f9307abeffe7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d912969a69ccd51bcc05144c365d3952f5af9f20c4c500647b6b51e68f4ce94fbd38ceb3c2f718a2fdc8ecff3bbe933f8f3aa516c6076e847cc305acbc223db758725505eeaa2d979d0f94292d6da9f66a5e84297b52b36787c8b39490b1d77dc302216dcbaf52f1fdab8b130bb3c1218ad80a9c2ea93ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fe3f8ff39861ce7c1914c62418fcb5e8b21437dbee41ed4cf1ed1cc1d18d3153675cdc70a82fe7d9d7be33b1174a397f75ffcfdc3a02c20d36bdecf4df40d4041ec6213bb58bea99ed334110fdf40bdfe90ee1b8b8d0e1dcbb0a9fd846ca19f4ce63cb0522505e8b4642be79bf6167f05636d4a53608103;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbcd253a87bf827cd7d5f9831a49547f4f7613d96b7201f01d2e97530c0f89d00d6fb38f708059b27c197c26eb01eec43eeaf716fc8a136b62c518defb7adbb835d7fb5d8e8c1111c21697eccce76a72eec5839f0f2f4d4501269b70e67fc5cef219dc47dc39627c8964b6480e20bda84f7b98471ed8e145;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h112fb2d2c004fef41c6e4bd09262d83aed16922106ad9b70d0f44d41aa2993de6144922f8b830c04c995a7ddf1eeac6340c900d7c13d4be216045db45b67a1bdba552096f880efdfaca4671a0afa7ed39166c16909412c4b37cf10aca3374ef834419ac62254f9cad5b4b82dca5b668726073e6df79319c6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e31afec000102be626abe589c383908beb9197b695f930ae1cbb699772f4c93566cb786e2804aeedd5b36d3fdfd3f57890ee13fe0e71b6a2a5a332d4a56dbf1a3990c67cabbd74e2377d61e35c4d505b61940d8d0d6c1ced522630de83640cea1b40e7d302e920adb746d6e646a185e2b5f2585e4f6c7bed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bee9e0cedf19f97b583a1b248ff02f07a6106725a90967d9938f70111aa657f00a5810ce6957c8a08b9f207ca640d40a9f6093fef96c38adc7d16c29505eee6de897a6f7394a289cebbc47f2507ef87b2dddcba48dde104171e71b98b036f454aa7f8bc239abf032b1d100729273ebbe444fb7b28845f84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10072baf3f0feb672dbfbe0b3bb4f230ff8502b7c94817bfca2049e08043ba77c18453fb6e4ce8ba9be8792fad2586d0c8dd9153f7d29f9912b93cf236061bb97d4d83f23f611f28259f1708c3f5204dcde75f2a3a3fd5fd5a35c2724de55baf3cbb294a75e9c4b750096fb37788a5c74123d17cc0beb675d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79d4bf44cac45c79ce967e1b41db3469adbc11dabfe73cc34037471395e118d63a00e4833d52ca6e3a2ede7b1d1435e1271694a6e127c9fea515003968322e56069b3a28b54616b35de25651269e6e9950ce024484e2906d00b40fe4ea486698f7f22c9cfe4c63dd1b934dd2828e8247e1f345ee39d5b580;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59d16683a3c9eab1829d6213686e66f8f60297fdbed4c5f661c8ebd8b580487e6659cd2284cfbaa9893fec261258f2a6dc6cb4721772bc240a7e9d7532cdae8db8b51081313a1da372f57528a86256754ce86cee4622084580e7530a86507185b40233dce02c366c54c13d7dee13155643f40c1572cd3e85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1509b44089c915bd4a310074890d664fa68ab6e3e812a083b205c59902010617bb49c4a4c7a518200c43112ecc7386c83300b1fef6b015b5e95cff196c4cc257bd9222be383ab94176f9310e7ea9816cbf176d2c5553e9f4d4b63ba131603a04c068394dd96b030dd681963f583844101cabac3f8f10040ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d59b0017bd6fe018f15717f2b1854ab342fe39c31c2339946d413adfd2976d84bc3a40a7e5d2d109eb387ce722790735c2b8b196d401e9c13ce2568bf74b1f67020046e73096642329fbefd036a6a8105b578ee1379bf7f207ed801581ef2eaee18bfa1bdcd1a8a669c98f3d7c2f6290456e4ddbd2e6dbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142d63171ea7426e4cddb1e8cbe053332b56a07f73e10b775a2bfa47a0ddbc25eaa4e4cc741d37799d27747310a034a4c1d26db4b9931fad28d79814966f48d1f8992bc5ae38e83b2eb66d056efeaaa5e8ec62802a36b210f3bc22a6df336d6b93111b1ffc119ee3fd754d22d93aca680faefcc3e87bc1003;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58f3170db244c419789e599a2ce5d0e83c92795f571883cf2eee0b1b4c9fe81c7d6ba005930b6f366c438ddbe0152eef918b37ffd219b0bf8d75e1ce30ae75d1a5436119836ddc6faf2da2dd364efb5d91962debf0c173e6af9f9e6c8c95740e7447f4bf60131f8e5e181e0822b90ab445b4b1c864008f9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b0b8e4de8ac4b40b25189de60a3c43011fbc3f35c299cbea264a4e9fb8198d83ac26c5cb375c3d652462d4d9f009dd1ad38ac5aba1c23c7cf37320e2bca25084d8fd1a23272f7af0f491343df42e4c5de55dcdef15b7c3981b0e957a8cbc0acb8e6b453a415fa49eccb2ad8e4c0f6645858247abdea65d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1007e3f5d01de2907ef62b3f6925b342647be337b3b08e6fbf20ebca34265aed5ef7a9afdb44e28df68ee547fd3ef2dc9698447a688d6eaae776f331f40d061e5ba89def0c6e36a95f7e55a25d8ee2068ec2bbd33b2a55fb4189ae46002a9ef7092e80967b2e26ed304b95d555c536a8e09cd09cca51a9479;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe48998800f48616510f8b5202be9b7f2f85ee7ab1f8c2a8e532bb44559badbcfb42d05c08c4f63c61d38faf717753e7cd368e042927ab7054a2009c501736a92406b959154ce5cdf0a49458fd5ea6db1838d3c228c1d91519b17c4b11282c09a45e4c60369df865f915da65be0a9e524b62b850aece2adf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2cdedd68ba9027b496001b730ca451c3f9cd83fd17e9b55f57b702bbfd71ce171994e3cb404e0a36fb19e73db9b74edf224e0ef9947987979cd5c80fd92ff7fea380a884a1a3b475faccd90c2eb8bd2382bf31ad7007af3ead923618d3520feb9bb5cfc83312346847e2c5bd219426f8c4d6d19f3e55e4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161971fb3ca3227c38bb4481dbe89ce2b9fa91b67c421e7ef489a62008293b5ac70f56a5bb9ac3cbc28a83a74aa6ce5b4059cfd0f5404aeba39a9727b844c6fd1bf8d2fa8aa2fe4c4b16ae2e6fc2df107d2c2d7713aa6ed74ce4b119d46e1352e86ac1818f742824b7e38ec85cc8b7a2db9e9b9ac3fa2d6dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e2b7b7f6c516a580813cf6bc372e91252fa4d75a7f99f75e1a7b43fdfdeb3ae086ac797cae81d1d3f9b7c6aa2d7b994a50ec2d307c0587cb1dc501cb5af9e8a6e9c95e3b79fcfde6ee898ea0ead6bcd1291b49c108ffd280487819688a50288587d54e8b644c2a93864f1eb38cc5e818afa3b09183dc771;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c45b3bdb67195a390f7adb63d2b92acca4ecfaa0885634db77936fedf9de7a821f1aded9386413086a0e78c17381adf3cbadfb16691548a3cecddc95fda8dcae4cd4aae8c4721b689f94fcf7841a9c0b80c3c39bd21d69729a05ac40448fac7d8e2eae82901e2bb8f56c37bcae76b046426fde2534fe7dfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea11a7c954d11d855c92dcf7aa7d2fce7a979f5c6d9d4c4b68222038a23580e258bab137123f53866779aca2bd3a2f7e1f5e48081c11d866dbb44237c97ec3ceac288da489f3450cee2db8a05963fe5b12c9bd2be4ba8fc0aa8248c594c6d7d41cf757c71bc798da6f8f6a113f872cc84644e6df079e978d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83ea5f49086363032275121550ca2f3f282929306fc6b99b6b40d0cc0d66bfbdf100a79521d36b35ea1449b9b9a96f4e24e1a2ba2fd65a1d5b872e9094536af677c7220613e0d2658d18883a2a309c9d37c49a15f3f413747f2cc54e610dee761fa18e720ee02a6ec751fe621ca9816420a0e229aa672b3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb53515ab87afd27730d75daa7439408206b09d62a69b73bd64a0a263fbd117678c045ea1edb7272da151e8be06f2f0dbc696fc43e50bcd4d1dd242c5f22dcd4ab54f80caf0e2bd501fb460297793eadd3e90cf93b89ce70a0d61964857f07f99fe51c518a108b25359b6a938c544e9f1c14b99976ebd2ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151ffde5b55c556e4352d58d65507649d2a7de7a9837aec19ccb6659374e9f1ef780dfbef75cdb99b823eaba2fffef634bd36ef87ac114a887b535a307b2aa5b03782b8f501f43588376a134fb33277b71584efc39ae86972355c2e1492c32b076e917fa0227a6d015deb7a1b9163df054649e578a046b942;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc29ff671574fc0da647fcc4389505a14a551546eff3b0302b14954bad4ebbf0434040d6754a938197e3185e50cac831aa23561889ae66aae37de67d7b67f28503dadecd5930c756feda9f3b86ca688f820e2eddbdf94d0cd0cc821e575ab7d0011432ae0f5a1149088673b60a71d78682794376a03b1a2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13446d74de76ed14cfdb68a4fa0533475987e3d32dbea1a98e600eeaa46a5bde31ef0d96ab11e064aebf58a1995a3f6e703f598d9e8c4c41cf5fd8ae970a3611c81cfe9c734deb32c580800e90e93259da91751fe60dc8b8eac63f202089cabb1926230579dcba1cbe2f3320ab6cdd7448d355be72bbe1701;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4933abc8357f01714224efb8ea061696ca4672eff657bbcaac80ccce8ea035bc0e240953209bc51b884695e23b1e50707079787004864f619057f46d93a58d21c7d31c619361934c3f2c5f752716a9eb702d70fee8c4a437d0cd77b065f967cfbcf09cc80a6c981f61780a382484e05c55c46033c44f54a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab557a649b973043fd7e54caa60b63f0bf84f88058ff47ceff9aef8cddad617e7a48ea939934cd8a9307fd8b60fc12bd877e06762e07b004ed2c9849bdea6c185f59e3f5d7458f0adcbf1f9efa38d580b31ee1bb91afe6d2b2b66f5e7ee1af1f3b3928a02e2c07c85da7865e15f39d27272750dafe99ae10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca731ddd544c1fc0edf12d8742c369445957112be0a089bf1f036b99e6b627b0a3860bcfbfa0dde2bbc82a7d8e3ac27126c49c8146387993115ae2cf8d08f81e6fa68cdb30c48a490fcf4061b84d99fe58c7692503617898141b7d3617e89c797e9eec56d6aca1c5ec8a62953629437899092f13deb8f3a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe057e531b606da84fea8f77365d2378968175fa3b5a18ee5177d51cc46cba7e28db61dfd6a0ede0f4007199ea1054cfef19341bd2377bfaff0b7c4fed8480b74c059c41ab035d03e9d355043da2f0c848f0f1af0ec783767255d32a3b01a48cd090353cc89b7d03b3120622cde3b2a2c9932187e9e1ccae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e02a7875f97541be5a40d7dfac90ec47efb3cef4152a3b8f3e7c10a090c25d466e542ae728ac64ed6e0d1bc289996fe9f48a342db6195fa97b02f3f2686700956da964c7ab4938e74e66a72a5363a46c0b656183721a75aa1ed4138c91636747c0afd7fafabea019bf8dd524ff75c240fd749b23364b653;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152e5fa491ce137ce989b2c9c77df191d61b2d350a62a8af5a814dd3c16296e6d2b371654d7cc2bf9d8419c2b81d9f1eeb258ee961b53530499b5aa159a9a12f95dac104c74bb414b958c05b3f95e7d47e56dddf08dc859637df643c895cecf43a566e79fd1047a2ce929fe79d7c125ded99e25cb75b64ba3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d78a7690d47e31851f267edaad9385bb9cc7843ae13fdc6570d64462b43dfd650dbe981996c3c72fa23ef85124b0716c4a9b2a54eb485aa889f384e7201e0d2e3198ba0b91f1c9b1ff639da76d44c40db835a66ec90baf90db5b2556d9befafc736e92be6e5dc95298b30751f428a87e4f85d24642d3575;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbda01c54d194abc8912fbd066e32f3680d641e915715223773c1585271d52b7894b6511fbaf344f35b6729a37875223755ec2f034c20112102da0425fd6c1b09ff67310fc7d2d9a6ea8438c24816883bafc95eff92242b5550d9d73c5181ec21071cfb3f4e426ea0fe6a2c8762d40161281923396f3cdebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135402b90496d7da5176fcc8041742037033173eae65c34c7125d7a6d3ba18632d9de44c53422b1f2204696565acf347422c0785895c281bb1e11f53ddc0a506810dc3fef11b6dc607042f2774795e71baf272efeb6a70ea99744c6503b3f932cb243102d208590572324e145a1cc65b2a41e9f9605bb355f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15aa6807b3c2fb416797eacc1d834097b2c39ccce0fb85dcefe748d87e8080ade0b05153ebf025da6d19250e7ec3b0c098c62f33cb8112a028dc762cf51dc560a60869127fca8becca7feffb5096e25864924b47d9aeb64b7ed9d1b57ec2cc254e199a78379e047b52e3dff420c47010045d4390340e4508a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9251d3848052da3da8a5954e1abfedfffb7634ef2a26aaf11a8c2cff2652168ef120ce2ecbadd5b03041ddffa8ae31a312f24d525d63789c5d6f3fc1d9df9813ab9f7f7bb5129f6b358e55e4c694ce84e53d458d170f2fcb40c5e021f63af7dd7a812e72ffe466eddc05d1c2cf5fdf9c08efb3d486cdde82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1184ebc68ccde9d072ca69543ce6f3f8a7fc6a639ee7babfce40290cee97884faf332a7181661afddd2d236d88acb740ae201020d4b58c7be9dfbafeb5de6c9bd963e3e6bc40531bd982dcea7413444f15d62d5569ecd22ea46dd9e6101f5b0ce1d21f6350f62dd84a41366426c3db5d554e646ffdacf56a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1481f98f3703e35beeed556564cc5359668d5c2c2230037bdd474774031a402aad48af67ad94c137cd43421745d09960791682a3ceb08a038cc9a85ee5686489ea79c97946530ae0766b4031c68b74b4d47fc9c1e2ae361f9d03fb4403e80185dedf0db1293d7cdbdbfd984e4a071e54d94272a27e039f4cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fa127670468b1ccd098172a6433be19a246ea290173cd7f8b87bc08988189149bbf1fd160c0fd1a9aa1d065493042e4bd39e23b596ee003998aca3a402e5bdc81d727e4a1f1b5c386632ac2e4c48e7da45982167e0c7dcfd8a397049d15c2edc859b6119b1884d186e9e201cbddde62559daf14ff965cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e3ba0315a27ed8c1b50f99136ee7132db79204011a17926a6fa7f813f845163631b85099f3491bd3bce59ee051ab0ca89ce50bf52ce96b9ec46dfbf9b95684a5f9a418b71382b1de3b0f0714a1d05d00ccb315c8a97e92dfc89640b267d08b2af07a1c5d68e140b2fa20a2da1a196eca0f8806f5281179c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfeeac08c7839305f8039f7e855ec841ec3b48ce3ae70144a5e4ac8899871278a43adfced60b0faec43b5a5ede9f3da3fe7f4c3ee27eb62c0e9f221c6ff5471f0e16e89264575978e318e0295f369bf01789f6198b340a0b2c9c497793dcc8d17b9368804029173443ace0c8397a89e41295cf1fd3ce9e5db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129be48b96afc494580e8d30e5b8a12c87135f451923fe452164faa9e2f2fcd70bc38744341a474f244bb83e1612f1d7058c4715dc4792d8766c59c854607bf8e770456fa05fe34552ec4e38755aee2f2eb4a8e92a7dc7b4a0df4a1d729785e13e186e0a477932ed33a8fd1b6f0102345cb08e3fe9cb79d63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa0db311b52fb6ae32e0cf182165235a96a8b5ec94e2680a6149e875c47015e468b9b500499af9db4d35e9319bef4d0ac1ed08381abbc92d9aa4874302e4de55b90473cfce284800009c0febb5f60beb8ad5f47bd4ee5d0c34061d96b8cc4a002a94d3ea3e64eb859a2b7a63727e115d14ae080e50035163;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bade2bb011863f50720bbff96f297038cdf538e39e7dd91ddd35fce5a918745962163b5812792349f17cbc4874305fef214797ff62ee29173e49b854593c4ae67f616191f42c9f8ae8395960487e206ac106a0aab3cc53c1343f0258f2481706507aa0840688a2434807789d61b84513c81beb9e0ff18077;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f05377547adb096bbf9bd1744df1edbe145c93ae29fffd6356c9d3383e21f3a1293933f4df8b1755f199ac8cdf8fb02ae4cac2ae3417829a63182ff372fae190342a7a602058fe965ae197752b666860c444096b6a684f207a5e6ddb70559b27fd5c97b8903bc9d486f7ca51b1ce76430d47e33a5f5ff20d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c241ec6afff80f7ed5eec37c1e554f16b580f40cf5f8b14e3f051851f8b0e6cf799c8d231ef8d80120d01cff0b173ac20b5dd49df346baeb4bcd764026dd13a41c56b8a0072faa0ee25fb93794ccc97acb37a03b8a997689096a36acc9880b612fcc86ca5292d372a17f9895e6b4f0a8662c9f71b9f4651;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4cbf0d38486c8fbf2438abfd5358b104a1d423053bd3a794a43f1c91a9be40b9063472afe6c347e19126a50ae96c24375887658f431a5ef10d107e3e23ab3a461a60d8961542d1fd3ce8f14eb20f968671710e03d90cd7b05c293fff00220e4683475280750433484761ac21eb55cf87594e94716b320ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a0aceab142695a817000f72a9839d16355820c86e73808c648057d622d8f50bff05eb85cb31d2399987971fc9dd091652c84f600e95cc47fcb171d3400bf8a03a6a279243d2a3efe9193382cdb4f5b8c63538042049862d994230e40906804ae644093d2a275f50a1957a6b1679687c2b329ac537f09523;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29c326388dc0a3d34d843438f22d4303e50b0d837184bf533cd6f37e3f2e24aea1b181044cb808238b9ffb09c2ea7ad7762def24032ab18ad1e18cad036cf1840c650a81a71511df780520ef224203611b25c7652d64cdc86856edc9ed9ce8dfee5c4d2d878794d8bde47f0740e5fdd9cde4acbebb7512a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9dd964c095df84863e483b1a5f2a649dc23e529da2e4ef9d593ea02a1c24d05471fa35fe98eed00c6b698e01ec7d7e553026ff513bc3e6465f869adad22c3810a979369a8a01d92185bfb79c68f30d1b7a193d304f3aff389f13534a6d471a9cac965ee110ccc51f90c2d6c0f5bad4221146964c868983d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fee2eaf6b48c8dcba6f531fe43f0b77279e35e756b0785ff98754dc6480f91dd2efe2f790c29d24c8a8b42066aece9eff593f0e57fff5e06d45782fdf3bcffe8e6ab6590e68e81192070898b195977e9bdbc083f4bbadc95dcdaecd9fc25f7c99beb4349e6e27944e9463e4d42cd23f9fdf49682ac7367b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14848929eddfb86d11e10e37439c91f9452fcbf0b0531cb24f0a5810809202bd35900df658cbf697abb1ede534cd1291fde7cfa304904b5b4f5250f05ac1744278ff23196395e44e32df0c5c411a55b7bcffa6ff89282f442aee13ddd4905446cb2ebb2f8ba3f5b0b538c2c2445084dcabf767a11a6b2a069;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab5ec7e50e75ab8ebf0010a7e9e0a3c5e9479aa3dac9f9abb7f33c70deeb2a0432a23e836aa743a563c6cf9c1585208864f954461c7a2fb46faafe1e4ab681b96736a1498b212b1cdfeb1f5ee996236d4be7df24f979412da00f82643ab71967575bc336be1b583fa87bea409261d5df8d4c9aa60c46505f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a643590891e9d583467ba8d78ddb90998ceb3a72edb54e5063bd9360fafe7f7c5290be5abe49839847989d44bcff1d9c14052c1b14895732ee0d9f3b062008758a35d6592549e1fa2bd10e6964568980a1f3220a4e70270092a323312f9c5b62e3421b4f596b85801f93cd2a74a2f826f546498ade9d8c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1600a2b6b81a99807757076d41c5c4b30cfa286b531a200dc5a4726f18d9ecf072208903243a90331d06f35fefe2724ec69269300b2c889e231b77ea624ff15dc536c573e37d3a6b2ef908e118ac40038e1a1ef7e6334bf9c8f80c97d222c56dd8764525d1afd755ec0c2d448e7400f0cc1cd1fed14b73268;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1781974b2bb064cbc83be8aa15acd365a05bcfc80e38607758029c08ddb57298f16889f563dd1e742fcfb2d3b2b5ea4e9b1ce92a54ec9e8cc109a88e17c0d535d4a5f82e7355f3a61bdea7740b8a6fef9000ee39e1f2ae4ac0301568fcfb058737bba9fcbd75924fd68a3ca92e7e0b2d4697320b743b8cc7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa2d16c222f042f6d10c8c91c2bbd57ece3c95ad55cd69ee4b6af8889bfacc4ef93bb413c18403d250714661ac47d4d0784d7027868430e38dd57e9747c8cb7e04ef33e50ddbe888aa3437ee16c51a2f8ad996b40a4adf0c5635bce0c2df5d7ebab5cf632a3fef045b5f39547db0756aeff72f99105dc066;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b0f27611cbed7e4acdf28a5c518c811a219669584516300c1ed0ba7d376f420ebe3abd206248897c48e95d2205eebf940daf9d26a87135df887d5b1e3792e37a0c7e691a5fd330c594309ff180752946040535d14e41db763c6155c5538cbd8ecf9501a5eb72f697272b9b2e9586fa5d344d90890d2556a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heee740eb56a75ceffc7b3d7115c35fdfa0f531b66dde7ac11b071f30a2390a00f44587003b33209d656d92f7f9ecbc02a6f742565252cf7b088b63374811a4887b7726613a7639110c5b4015b0e145c2076b3e3bb8cc73d7d85ce57a0e415b993b9d2f58a588d94be6e06bc68f6498c86b393e46339af208;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80b3410262979bcf3868075ac0533cdf129f7ad475686e598818ae77278d337fcc2811bf1d0fe254a04793b905189117c6792cdd71ba68af715c1fb4dc2c3f9876701ceb9143a4ed8c9078a0315a7a37deaa5d5b63a189cb518b53c2002885afbc05ddce80937c125684e6a1d8ab231488a6c630bc9f1dc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa8b92f66feb281ab15c843722706ce3b5c079378971e63f43b8dda0b34577800519e5a02f27970e83dd5db78bd2c7d61f86243e95ec154ca0c3780bb623de31eee064a434b429408642664cfd9c5dd2dcb6ece17b5025c904063c10f5275812ade84e8e0a39cab2a346aa5affa847f96f1f4507b89eb6f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154a6f29d5818cf7d9a58816532618d8aaec372a311c3d74349af51101aaf1f1dcf8e0974c83eae48438636f688cd5b6206f03cff09e16ecc63781a20b487426fc4e57dcb9acc82554fb8c2bbef9fa8b5363791d30f00f8f9d04189c6365b95a2e9e256cb2c95acbdc7a8e019b53b52deca305d8f092e6f8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h971e7927ad44bc5e1c8df0f8a184c149bb07a8ccc88e32e42495e2754547b26758df729e55a8b9cdd9d98a8ae634cbd2e9d0ad5f2ef2308598be0b76cb191737cf7e8a54a5e0a74cd3192b9dd5f01ebd3024a19873847c4bbd1f0786cd52d6170f28a274e6f8b4a912e2c56b60818af8cbc95a82409bbb43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108624f8e2421bb7b5a07d1a1637e41e6378afd7dd290dedce9110a5ed81154f3c9583e5452ad05e0c4789ccbccc71a2ac21825f65e9f788d5f9fb27108029bb4d903dba92631f1b82bff41cb7fd78940c7e23b2ce9fac205b4610bdc40806214312c66714417e776b0312c573f713fa5569686d6d786ac28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2e1e204aac61b390c94b020ff54347389967868c090c425881238da849f61e494c8e5c0de3c3506e94fdbf24d48a2e0140529ee04070361da62b88cd4d0b6e859fedb48b3c3ced83de34902f9828a7fea364c52ea4036255aab2c4ca0def458f02524b72375bcccfc486fb4e9b5b9eebe9fc6b4120581e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h467b1197339c67e51c42402da902ff50dd680ceb73d56cc8c458bf4447923113712f4ebe8a2f52688156585d548de3e7e13ac19984edebb4615ab7e167fa9282a63ee59e5b6ef215c15fd3d3aab76b6d9cafdea02e32e21af8023a4b79c96e57de0d1be25e02ef4389d3d72b57798c38da4fd97fc3f6316d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17799404f9c91e3a7426be7fbfc200ba24758a111f6c382fdadcc7256c2f80693d82f3b33a411134ca61a4fe8e41ad342223e8f7c4e7f76d1cbea120b4c9bf237e71f7c7e728a5c382e36065b38bf4953663d905bf2ec59d6b9b2f244346dd4a149fc235170803a6a7adb44459beadd8c7d90c4d983291103;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d7a9c54253ddcf928b644d63d4d2ab9d8ffa5d455a59ff584a9406d74cd5434365b708c65b783fc980f18ad784e35ba92da74b4b829453e068d9735eda3ce0619f79aea413e3000fedfa803ef3d0ea9319f26bd932dd1b8531969fe4050c514c98cbb76e7678328559bffbce2071aa79c14748b137bbb12b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50b5654e10cf713e9b98ae72bdbbd8462ae30d789d74f97d7cd407622aada05de1b1d39f05ce980850531461f8ff466178095c34c1bf5a532a3a425fd6400b44406d4a4e75c50538edd92c1495b66b6bbaf9783fec406058cec981556eafdd702197ce5b169dcc49a51202c324c3d3abc78a9e0822a98836;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha83a16405d6aee327b5307b70da60a546428c82c660dd3779684eed954c5715b1fdd15965729e88521974fe09d8cbc29b1716a1d42613dec6b7893d59313471d079aef37f2056295ea703764c141920cf0cf834aee8c73e930503f87e888b52f9301a79413b6907fc4de8bd60b2502497087525d67a8b48d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165a5942aabef8d9cc55704c1b8ee11a936921bfa56f8d1d8ca18fb398b8f8633901bfbdfd740953e733421dd33e187787273689015f4abdeb83715fc17bb0db218b89896731ccd46c33dc5b4fe02b4f52e66a0e3ff06b75831f784dbee54984d517fac5e6edc4ef302ce34e31347bb8ed28b54974c1f1b2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166d71510b2e52a61e45b6832132a185fec4ce6a44b4a1c76c7edd18d36ed20d1a7e366ef94ebb9e4658a56dbfe58b8434d2043ffca1ef284e1f48473f6a812b76ac849c01113b89a5d2ba33bdae57d1cf7d47f6b34898936bf3c6c29fd4e249119fb00f358c39be272a921ec6f36d2f2508f27748803645d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82d1de2bcac4a5bdf18ef52b1a97133ee2c7011b833b1feebaa4c17c81a513a4e480008126b7f10f3944281894122f44f12d3b36dc07661e3fc7a0f8be04d1e78f7533ba3ec3219fc0807546d90e3fd79be44da0db6f4f7912a05d8eef08dfec5a52a5fe2d81d511ff9ab919b85361cc5035fdd1f52ff1eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17011658707bc606019ce135eab6c7a74f13258e2299b4c01a57389cb82dc38e52edfeeb13d773e2ff43702d60648a9bbcadbf3329e5ebe96a09e16471f2d9fac0a201d10e55d5866e5d6ae9c351df5275d2ce13f955b1246cb2b6aaf807c8763b1cfc1393903672a428911862c5b6175c0e07cc3040cf96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a54e000f001469f4f7355253a82e884311fc5c9601591965de0ca64f2560030dd785f5aa4b79240f72e30ea0b920f8551aadfb48efe01f90b57a0dd952f024f6ff90a51331d3445b1fe35d0da1d396648be74bf257e6e840768ba6da1fd03ff049495a363436bdef070a6ad7750090b6fb223a5c89105dd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he17d161b071b67204a92433914f53cecb231d7716e15c995307d448e0722b039f6e44c36fc17ff0c08491844f2d53cf082dc085c391b78cac4e259ae1fde4ec7e4093fc21361a53fc9b357c5a3ff47ac0dffeba46ff99444bed1786c4c0d1adfb200266ca041ae1fbf6f8fd6a3fef6f28b6005ea3a88ebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb7af6491500d0bd19c36fef1538b66e782c97cd9380f6c6a93fce84e661d7abaea16bca90dd6381ee81cab9ba1feac16728f4bf5382210e11862034deee71432992dbfbd67abd9557ec184f23cb195e3668604c9b32bfc9019c7f06b5a0029d35627747651f6663f245a084b388ad695b9a22477185ea11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147c973a2587070463b962443d9c9459f4a629f37ef2edf3ea79c0ce862e6287c0416f2bd6e323c2db57406535121d6d141baa32133352ffcb4e2a3090267a876cf4765dfc0edd5c9d29bf72ee3a30d28d49d27ed8c4ee8727684229c5cbb9ea098ecab22b8735a744281574cd421c8a9a8eaa61f5e345f9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5c9bbd6b057d35e3db85d4a8b4c365b6cfe4fd4fcf4147fe93b8c6beeae3f7bf40cbee309f8571794ea56231b90e8cba68689b7585478a2f2bbf9212ce9ab812ebabd19b6089a9c88eb7e73ff863bb30843306d4874c4d2e32e232b33f1fc0cbdb71b39b205fca4144d1df89cfff8c35524941d0fe87456;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he07bae0b73cb602f5f7993145d494732c10dc104c149c9a0b3f123c6186c53d9a4f5d41072dbc207fd3d91b801c03eee462e018256a319f87a3c3039c07d93250a7d453944778951bc53af5f8473e5c1e192bce9ce8de5bdb2689360056b0d9ae3546e74f153fe6d212b3801eac0f855228de26eeff95f8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de26cbe0dda5560b7625ea81314f01612d08185fdae38f4ec52ce5867ee174d155f5cdac2d08485fb00d92335b697cca783a4cabe8a9817ea47bb2e7e1a32c8680b76bf5d516e5aa403c7d64ebf2ec8054de8b27a3cd1546d7bf4595ff829af0c282ceda7608c5f0c8a6277a3bf3528caa60a6dc22e3e244;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fab9dbe0327224fa3592544b9c9cc0d1ed76fa24bdc512d1c52d24a78b44d8f43ff1e8edf2ab753e5285ac045b9b8344b027b83fd8c82bec24945da47e4c7397f7fa81e8c41bf502644f27891ccc72ce7b11fd4603dfcae45f884a3d587eb9184861b5fa34548ac24d461320e4eca865ba8ee57f2030d16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c011cee95c7078ab6ec8209638294726e3d22fcce671b0dab5f72b6606a99efa1e6168b6be7bcdebab17d0f30191de679b0204071876c1cd2201b66efdc88c75968040f8d8f20561ff68d80a63b347273f8c2c01952ea7d28581d289ef363c448c60fae3f69fbcce77bbce4414846460cafe900c811e508;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1d1469b697cb0b63e4e1c2028fc73a7619872f6d672ec148b65fb0b9baae83b6f5f44ef05b003f0ddee2881b0c0d010534689665fc8769e7318a30bc98ea771dc580ddca7e6cc2601e80720dbcce8da5a74ac9c2fe34d6f9f2628f095c54fcecbb6e7d7aeca904efd57a15212eac6a28fbe3bf3ef37a47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8d203362465b090350a9fcbef80a94d99070677a0b3224eb7a74de1995528912888182e02d7f5f204c74e9cf8812a68b143d2f9d81ff10b44fc0dfa1eff557ff8daf73acfaa07392c1218c5ce65179018dbdb1a4f3c7a78c011f1c84d9de0e92efc482da818c4e4e91d1c2a5b43647f251ddb1d0a555d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd0d283e57190eb70c31db4425adc167799d249bea1f60831402875aebd5928587758c7d7cfbf4dfde3ea984f0110eb44676cc1ae3c5a5ad80208dbf7d7e82dd5d178bda14f8d8634d0dad1667cfe3fc110c4295b06f288bbc6cc670b974b7387930caa159d12ce9a323da683b596e81f4a4baa8cd0094ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1c2b5e841e44e936e16b74af2849448976a084149ae65e093ad43a1ebdac26be40758e4fb8b604bcc34065d063a801116671db2abbdd7c8b6be92dc8207b71cb624bc5cf12a7845c43546ecef335c09c694916733f2a723a545bebcc2b41897a7e4b2b2884fc26976beed6b9fef47f0eca8c6d52674ddb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151435153eee46f1a715c0a2b50728d0b758313cf37e4cfad7b3e3168b0b13a4c37d26961334942bdb0eb9bcf914019b1c8f55c08639ec774fc1b7978c4d0f9dc3d20160d5baca2b47958b44a0af5a767001771e981dbcca36e5d6c0110126326624be8158db36e266063156e1ce998cc8f0c79521902150;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e4946cc7a1d4dff164f15de8949dcf8020fa7f3ff2146763cd68f4b03cd8afd4ddf63e75d82b94b9c87a415a355e24ef1e2171f3c873945d57f356edbf5d53767f016691d69c1a24b010e00f013130c0045431fcae31951a185bb571ae3427f1abb86494832e0aab5ebf74ff21ec472452ebe9360ca95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf56f783db61aabdf6cbe3dfea8b69cf2682ca6d1baa9fa0cdac496a2bf05d6d5e33f13669e0b75cd59ed208622ae03da215ab591fafccd21407ec6a089874cc0a6d5a215d907dcb635392b7d1a9b8b2fe3e2dbb38ce210541901fd5ad90e31ac24e313e91b797c6736cf670f7a3a1f0a0d5a15818f5de91c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172a2389b6ebe2761db1de17370dad82c6f615548b6102099eb31b0aa88a84469a93052604e2b44d590770da758cd639562f2d2bfc2b44898e6159742149893415615456692228e0142733570adf939e380dc37994d555539b9b2b66571110efef4df0951b8493d907dace07a46cc31c2bf66f90921d6bdb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2aa4a613f2b43ed770047df677b9e60ad8beb6ed52920e9185de2ff2ee46120214084e9a9a45b8abb0d9f36a4a77f7d39260204127480311c603a24b400ef989c4532538cc666f259f545b2306d2fd48c4e1e2621bfcd6f0ed247e9d68bf5771d534e7a4d26ddce6857c12c638884053428096328b33f659;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7462f5579a3598648d8968a575e9b10697e184e072386c839261093d1cd114becf336ea0869134f50b2a7fc4bb0d161a4a7be7bb4bd2cd8285a511870f4e2a3ed7cb6d180d2480db86e818bdc85d3b31f67172bc082322ae32c3c5a81d00bf042af959627b7e59fe0ce8f0c8468385f50a00b43cbafc39e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd7d78b87d28cfdd13f51485b064b0b8b359c1f4c5d828932687223240ee9b00e0dcf6d49dd486a644fc28c4be3e86201cbcf954e66f92d43ca2346661b543ba99fc5be959622d065afa3444068f1bd6bc16b1504ec682c7ec65bbde8ab4279c26cae7026141111a14fafb5a546d8bab0510c702c08f941c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbdc759408ce67cd195c018ba6660cdbef9fb1691c41e688d9868f7f5547b9d98c655f026960502b7312210fe0498728890808fd4b28f30a52117a6a9491521ed3e9253cd4b56ee34505d9693be1304f6cadcf9d51e5be56ce0b087e23668f5027b5ee7fe4439e7e2bdcf186652fa67239862ec5f9f95192;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175ac935d0f5c662c38f53af2bbcfe001e749ce23b5bc0b318e351073588f44dcb18f7cee328aab5be0456534b7471a0ae54562f919e2be1424f0f27dc0f952c69730c4ac41283ca24681fd0406d186ce9914f327c86e850d2fe489bddf047c4d1d1a596b33ca2dcbb7a208f24647be49f587c5044601225a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c7a5b1e486821dcf69686afd56f18987c77cae96d6af8408d50c1d2f3b1b764da990bf27e2a94036f88edc948cf90935a60f4da7ef26be34365239fd497c78f5c08c2f2ca10d69c4e2f66947bab8438ec4fb2fe3171f43353adccd2e224178e79d548333c68d858bf76ce7898cf9cd728e7bc4d4225673b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0aa801169ebe60bfbc0eec630c6049d39c2e282f57190d3bc436318cc99b39dfa08e9e20947c9617563810e1f9327c46907f5b9ad6eb73f2794630d5a023a29f0b60d6049c3a38c1d80b2cf723097af63e729371b2dd947527b8eea938a410c2e50759b17e486bb7fd9fff7bafcf635c02369ba53871ab5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0f9041ce4b9f9af2d1b30b6481ee8063e0b3a2abd5840658be2648b34c30baaedfb8da596f476192de54fd4431d932c3d2d0af501b72c87dab96d59fa701e5bff75f0ceb823053aa17d8c9fe4f5c5fe3c1ac32b9c7c2a1f117be6da17a355b6fbeb684b0a81e76c44731acf87b19517d6b03658aff4e497;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1358fa1a2572d22c3d09eb131a19cc26e5ed0fba6dfa71f55b3001fa05c4fdf5d3e79ba0efb2660fc0fd31fc43aab4c4b45aa59081b928fe1e4a2283d44f499b05b0c95534fc4d201d782d7967052a741ef5d02fcecd16a55e15926d20d118fd26c41d7c7ce14792489c31b2064ce4a7407c902971949e232;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1181f163bcc30f13f2ba5ffbec48e7a6279ed3d76d7f8cfcfb46985e3a1406ae5e572af9a35d24d2ba8d54d21454fb5e1a3ec30e5e29ea8f0472030801c4f95252060b9da72ba43e5a9d4a6272075e31026f8a44f7a4a61d285ae1c131b61bb14e17d330c4b9b07cc0572e35c941d857fbaaf10be103968c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb54c5fb57f3040b6388f40f520a5ae1ef84dc6ec064afb6a365369803315e4c69671f025356cdcd4f3d9d2b35fad6edb8a3e521352e01690e9f6f1f2ebd64f164cb2e2a843ef062d2dc9978ae7b69c5c5dd7cd219685398af123789efb5e80f40171e4ba3a024421779991e91cbcd9245d323fac85dd3589;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1985bf61d39cd2e2b5ff32d3dfbe9aeefe0fa0fdb12e0b6acd9babc6524ad856d44f18bcd5caa9539691577efa87da5affbdff0db140177639c76c7b0502decf0a46147ddcd9d39b98d39b1b67fce9a63321de00d5305c93487a30ad7469b1c7562dee9c6d3536a469ea3e01e1218969e135d27095cd58d42;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7829b651597fe423b021346d7bc6c7ffb0779393041d5cd9329af8c852d949e712c602b1e826153c8046f1438bf6aaf47b65430dba1d44bbc65ba8daa10add7867e333804e796cab243cc6c0735fd12ba9ded954d779ce947195f0264eab052b0cf92f03e28b16fd757796154fba4bba2caa936e885325f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102353210352278e24d61f554b8efadbdc9e54cd41c8de47f8fbe9488349501bb9739d542959573b9db323f6eb6ae792f6e30791fc922eea0111c5d6f9f1f71b7e0720e565f23f61ce26ce3cb404d5604a9526427cdded941e6b4a6896601643f19980a8465a8289d8f6d1e08f7482ade38741ec5f500c493;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a719bfb4a2d72872285ad7798b760e5a403e875888e2d2d5961aacf8d4b0c08f43944eb0beadcf783a0ba6201dbf2d841f530a2a5ad139f6a27636ebdf76f3c236625f6b64305b93e6c18a4e8860aff78c654fcb6a6384b5c0da2620a26bbbff9031595c671c4869c7d5e152816257f4456cce1a58d7cc34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafb552c0ffb9a219fb1ada96ed53f53a7050f496da3d0ce88bd31fc07213913ee58b3687c7c2599764dc16ca39e69ca5003fb3c4badb69f6c0480893b1255fb5a50637d59138e8d7102405771667f199bea3ade96f7253de9f0a91ba17f8c26ba880c1dfba76f5b2fe920c018d47c52df0aab85c6675a92e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9b61cac482822704568aecb249b0437e7f7c1d894ea2d6b084c6db8ac6f0890d43d43713a3d9636178fb6099f16e0031c819f698a6dd4666dd38be770be4eefe838f9e88cb76243052bdfa08954d24c03f5d8f12d427fe01d4124f6c8922aff5e8fc731922d19066ea9d97625c0acf25826763260f382fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119e32de7dd5d935d99365baac021df7bedfd59b3aa7c2cb8cb81259950caf9c1074d6172eccac12bbed0e20a51c440178a212a196c15e31a7e88d7a49278365e7c2b494ec0d44ac4bfef2d0eea6ef01dac74bf65fbaf256e75c8f942ee3fd10ec9423bc9670dee7fcf33c6bbed8859be489f632884b4d3bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167974d07ec8c483a254de5d0041fc2160889fcc754b959ba9e295112a177b7d67fa25d8d9639598ffa7bde187362d39c25724292c54a1aed52d81404b206ff166f4dc8a139ee5621c448674aa33c015e89ee537f6bf7c0f707a9a53939fec7336f520467198d105e7c957dcecc45ca62ffc4feb6e22b964a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5841723d4b126dd299a76923c721cc430cb347caf6e8c275432381e543712cfdd99390e9d363af475db78e3066a8515958bef9974a176618cf09f4bd515c42ef54cfcb407bc04ea7431136c774d868f1779789d073d3badb6ecde08adb11a9a9d1a091f81bf6fce8a587fd4c1171daaebc36664be7752951;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b30407559f8f62bb253260147531724e59cf4418405ec35ce122f4a01574ed445c9a93c13ff190752d9b335c321c049387bfd6031f53b697266eb9e454aa6c64993dc62bf2ce8abeeca6f34a97de1e729255b17ca6e5742fd78c7c0993d338894d851d23fcb6057fae1f12c73e1c6a206f2959564f6711b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1927f964d61522342179a31a7d32c017e5eaf7e845ebae75850e7cec7a5eb45be1863f73e60761360f1f541b44ecdb392456db595bbd121b77b086ceac960a26eafd2038d98bb2fcfc86e3093c5b8eb1c08c588f7fe4adf3cee3166db9819b5db027436db368b6a27899f89ccf11f565230ad95c7af0df572;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be0f9d4c8bd98bbaf58a46efe13c2e910ee91004d3e7119444b733107b985d9a2a46094345fdacbf777055b436fb8f96144149516d5e48b1bfaa34917b9bc3c66bd0d04173253a11b62ec218ef9e69c96f6c0e67356e924a4ca098689cf22c789f2bab1eb1aafeff5e2aece1fa9c1630240c130981ffd719;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e00154443a0ec1c7f66b8d02936e35133e2fdf4d5497f21d4d2ba53f2940efe5fe60759f8081fa6113ee8887122316a1ad0dc9a78d31cbf5a9aa0b386f7e9551ded748df39d8b60b9c3d650091b2e786e5c739b3ff351bd1f20b91d67504853c97379a0c8471b588e87cb277d7c6cc29db1165eb5bf7218;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de7ee2083d67adc6590bee290d41dedf013835b395a56d1c2cedbc71fb7fd4e36dbdd38946bd37c9f1bbfe9a8a3b42311e1163521b5f7dbfb8da0b9df6c7d548efdb56a546f28693c0af31df671e4ebde1681246f5346e93e1d13d8cee989899c1822d6b8ba3ee8654c3221e34b6d5dcf545d16933e9fd44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6ab89156e402a5eb876156046dae985d9df7b1d8de41464c9bdb863be3346bf8a32a20186a029a0b844a36c3b9fa05228c366c60dc9fee3416a032e4b47bc28fa893256c53957c325f72d004b58a09f115e518952782527d528b1cb610f176d3d667a5ab38887ca1811849fd35683f330ab2f5f33da6ada;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8026b553d8c061e696bd8c767574323d563412340e36763fa6fdebb9d7e661a95d21ed5562e3b6c966ebe157a341bd1a623d3011b1d6812c69f5313af4c68b483bec77cf4223d1d780c4a706965c3ba86f171fd300092770f99fbdabd761af4f9786dfe802cc0ca0d2cfc4040e3739c730bf417afa775218;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd8c0fb3e251da8ce07e331bbe87f8ee8d4da2f067605a3102f3dd2892e0bffdb16c99cb78a696e1a28e12e317a6b26d518d382ce73ac321d856b15eac1330bf4def7384d353939f7991f999faff4406578315755b7ee277a896626a75f685df61742a3da79d04b7e86886dd3c9714991c209bff6eee6400;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31552b679e2d6078ede7692f7c50c8b725c8a2cef2d388df268377ec1f3f085e852c540e3a1cacdd21ad0812a3b35f844e837813d5897eb43b9c21f06e04851eaa0ab5b6aa7f63204db1d1766a9953523a89e9e96b9a9b7ccb6c7a3d4faa220d1928b164ddb37fe4016a902cba54e4153761f89d2db2c728;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9514bfb5657944d1ba6e2ee9faddb3dc8de26bc782ddacf50300c277853c2f7976625d49c601553e98dc824374c9f4d05e45e98793c99f687c1d5dee4f7e65b0fe130bda3391a04b8d1038a40bd907e0bbb52132a2cd3c75a6e5f98d1239eeb5680ec8f7dc102171ae8dc19a49d291bb63b333e506cfca2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14576f39ec0a781b72bfea9b900ef960f6b4238f2994597f5721c11d17dc21e6c47abbf319373d56ce5e42b0c452eee1a81399fabb837d2192de269851ebe95595b35d249224acd51ceecee3b62c6fbae601912b4d559bef322af532a769801691b74c11b5834cbca8c3037b97003cfa4c7000904b7877fba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62e411e2cdc62124cd0169b13b715496b3d2836bad2000ec268c818fd5b1d15bbe25b9956a0e331de5d6ac1a5b4532de9c28bc059e2c1202c4424603a3fb935ea8ffe8b49f8e42c444d3ba19686d7b205c1ebacbc817d7f50f601576d47993d0f05fc32790404412fcffcfa5f3128d4560669ef1d94ceaee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d9178b3767171377f033eef20569ee3a5160532306f927b762cff8338b3d251450633ac7bacc008f641d7e5c88b6a9dfe4bbdad73500d0d3b2d45e2bba79cf0ea74895a12df5be4ccbcac4aacf08185947196c2f339fe79058b31070f6bccb12b6685dae22df237af889fd93c27005ed1966309e451efa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd10c241c974c3cb63f405636b66c39a109876eba1939e546cdd2137b1ca280ee9fd8168b5e01540c702308ff968372ae7e50874f601aa06ba05c4b81b8467f49e83f11c63b8a859b22346c6250d21673d78d80f12c351b4093997e82ee09bf83344048603f8143f3c17e04d650794e123d56d760873748a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb40d6835b7a9bc3f49877d5a3ce9970f4a1d18840ecd5403bfb917b9931a63dd00174e7cb2122c31d95158099f3e661e5af54b9f940f85ee6f1d476410222f608e63c5818c455949462229e3358ff98738ffde31c89aa34d9ab5b499a2ece8acee436dcc91a12b2839cf21587a86bb11870f0096552aa5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15629cf486aabc6935f8931d9db8ca3c5df08dc71a0207dd1bb617397f02bee343f5823feed342f5abfd3f0e5bccf50bd08ef846a84f2485b81645ae62ec9d925448de5748f5cba4c6e90d609c0961ca159d9504b1acd5e6f3344dcc2e303295293b3a9043f54e0e98870cf7e2f61ab94a104cd35829b1fb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h724a086866d7b9f7816fa021a8b8679ce09fb429b5ebdeab1deddac9d464b128736bbdb87e5644a1d3437d716ecb65b0e9c45c5196eadccae9c8cb36f1d4fd5f1b85caa2a3013db233b6017633f9a2e3d495725c34e5fb8e2df3bcda3c548c4a30f385cb99a408b0e6ffbeda8fa1336ff8840fd0203ef171;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc453d4fabe839ccf4cc0a597d7d6aad396bf1d5a78b6556543dd492cd884ecbbe58322999ede653018cac725a40326b89b61cea8426388b5617005961eef5f738602e159b77b714578744ecbfe4bbe2a1baea572ce397ecce97d32357f150a507006fb846c19ac9e9671c05fb59269c8b6015b94bcfe5864;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3db7c205ab9762d4d391a401b2d006d6169e1edbb75203bf167c61d9a00c26c3253efdea74871c9ae2067dc1c1c582255a812cef1f3fa5c4170a1a0a656ba22b1e585cd9d54d6450496806d7a644901999b2cef9c793d6be22788c88f1a25c94cef9ef8814ae9b319cdb8f9296b29728339c06e06a6ce563;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ff0b693ce24099ec215f12744f4c76da4c07c7605a688692128ccb43af2d48ac632fd0aaa18dca845fc0063a47f8fafd713961360385599760248cc91c913c0d2312ed72eb184f360178880facfa45029f293a46c1da0fe7908698f131fe67f0c1be9e0ad1151243f729230d94f8bc593089f62f998d8bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48b52d77bc977adcef518ac477c495852f3e29f5c5fef863d6965b1e239900a7e99b432b9b296408fa8ef03f9c711c7fc60bae2194b07b196dcd9ca495c13d5bfc89e15b20ccb4db8345fdbb9af5abf8baf5380f8035260b813b4c12051628ab9e904610a897130e57fe76400c562af82f02a183fe26fae0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14649f28fd2ecc51407349bb0056e1621769f7d7cc413e399973c0a4a2183e41fce43cbfe619d81fa230bfe460f999f0cdc5da8a1329e3d6b4ee0eaf978d0f3522d0826dce3fb877dc66c789d96afdc14883287983ae9b1b16e59391d17ef4acc0097e191020c189e7b35d460f0dd5f7beed951ac12211b7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbdc6232d38cc373388674a00ec6370370e8a853e617e47a51b5d5d83b90b78684d2d7f7ce2834acd170fe51bd147f9e81279de84228c80cc9dfeca9ef81b28496403db188ae744dad20bea782b4fdeacf7e45b874992b2e9b4fc084465e7e69aee5d9f1b57d858f6e97b5586d0ef2841d9acb3d3dd1176;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a1fa4a6df511b0572b1d9b06db3d6c9812fef451de4d679edd5650354248e6526004039c2cec95adf305f607ee021bf746f687b8c613e225c28591d00bb4d830478c5e80abd584a2187ad9ce5a9f633d3f1867eee9f8a0967bdb14731ee3f0ff48ce8a2e3b478757b199eaf955ee4628a8b63aa7f366fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ab1b929f00564f988695bbe2b7e08287f8d6ea182a28a5ebf14e743ebf28ce8453dbb82c06b30f5aaed1b57f0197d327c2aee49e3061c4e7063be331c1e4868026c3ea57c8713e41be3869ea6e264e0744cab7865577c4823f480a44d6636621a49bc5bda2344f8f017b1f81aaf36320622073855e64ab0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16fd82d1265b6a8b9f3e116f6b68f1ce2853e78a5087fdffe88418e74e62c3a7825f9a1bd5ff63fdb1e547ad7a9107bf359f756c4e819ebbc476db68450e7259b83e5ddf3b752f21f50435e0754a2728fccd32d3d9cb324b73cb10fa52157e7c6bcfaed01c17f4aa36b7c69159ebe0cc13a95dd630ecc60fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4dd21878c9a3d8ca21522850914ba056083e59a61fb230609b5d964d2aa2fa2fc737c32f2841d9633bf34135a3475d7353a9dfc0c415b22e0f2576313cb990a5fde38d6a7f6399f027c084649b161649b6ff8412f06ef8a9e2c383aa11c74fd4d35acb080ca6c75abb1fdb2b3b513d0cab1c2f58e93544c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee6f0ecccdc0d501c45944423dac8fbb67fc6b43ee2ad71cd49f3b8852ea6d95bb7c346d1c5188fb68ba9f6ef59e5d4788cc98a3636a6140fb9856888dcd90e38ee4bcf9e605b5f13ef5799f045457e2ca60907c36246db145f9ec3527dff7a78b227a57e80c8fc2160b2795fbfc5e6256592e3d522f1fec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5fc8ee59bee0d3c2482104c2f239e2ade847eab4be8b2d62dd5e48923414ba3dc087668a53410002f75171d6b06facab28918c7539e0306951ae98ef9c80912266cbc24368896ea457b885d501c795f490016ce0f0db55f5b0175be05ba168fa4dc7c6b5deafed383330e8b0cc4e3a0ea979ab3f5c2065b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd10b3e344faa0b3016fd6b0535779f26677389478c3e676dbf52b728631d5ea270cddba9fdf0bf975e850df9f7ccdd29ce504eac6575887f052244572016d04b4a4ce502107c41cdb2d9ee159ab5d0f9104d1accd824fa677cac3ebac666080d1d46633ae5bcb78fc16f4dbf19ee9145331167a2f4091a84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9661d42e0237b714b012a98a836aca7b86be71da32d44111e519a04ad491809eefcce2915c78c8fa6101735f2f1c3ccdcbccafa30ff354dc73625cb95d5c8cd102050c5f6671c42c12dc05ff0e4ed222cb78b8b9f3ab5dde2861bbd080b4d9238183cf8626cb30e05421128ff0d672112ae8f8ba8bb5201;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13eea6c7a14a69780694beff9e350874ce7adf3fd9ff4a41a6f962fa03deccda5b7329ba4760ad946cfa6f74e1ef4f2649cbd278fde3d23d5a64681d114bed125798d9d1c8a4030efe84cbee927b4736747c0a202f1bd66ab39c4a7687fd4744c9b0ba0c2017d7dfe509cd0fd8db691f97bd7d092b73fc47b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacd71edc4211d86f164d63d609e20af26baf65e1efbbcc23cab8e6c8ab12e83a7af9de721f00b6270f6b8ac06f4ae0cea2272c79c24758489353ecb37a661743d2141428403f8ae23e8cc4067f5f5e54b6b993ac086cd4d73ae6760c7938430116f328673c61596750852e02cc6379ab3cf4f9c9bf03ef10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha680cfc376c9336874774a859cae938c8b20ced7fe5ace57e8b6934b06e5edf80a1b6de59c8b368c7bf5e05ff04b2e771087849dfaeff944f0e85b91b92d3dda409521e88eb6c71550e6c1ad459509781aa23a9bebca5ec5eb19ba1bfe4c7892ef8cd33e2c56682e386d7e8b6cc2ef55ec6ecb992e7d2fd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5dd56fcefaad9079bfcfaa46cd5cc9359e0b61ed59b153829431a358eaf403e40d0d0189ebca4ec35e08f847a06cff002a35228ee61a77415fb84bd4ebc0e0f4e9c6174a10bd77917fd0c5cc62e3fc32d7d7f5b48f190d9b233c0037d68d8b650ffcbf27500e83af31ab719df3da9c1c22039d6f43c39a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff02df4e8e955c026ede6fd29f75277f18f32bb6a981bad0371bdd3c35d35197b071b36645b9b71a79836aee4e4911c1a3e84135ddd51dcad2646a9c693f5c727b138f58d89fb4cecd6c6c59ff36c62ae89d04e77a376105e63a53b9cf1f32c0c8de81720759795cafc54059e94154d5d2c2198fde0334aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0a2872b9d7b82ff52cc7c9b18bd260f0c0ae41906750c5396dca6876ad46a46860bdc88b2e8661b7b4de708a8d62ec17682951d3b0e949dce08f39cb5a3996f743692edb1a15d685748abf19a5fc5afedfe0dfef64cef03fbf609ca0b3b435bf322d126ae170759a212f1c2016fc71c93320114619479bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ba65a01a1d43b4872a170a39d8e0a7944985202756405ec055f6d04737067c7b0950a1a0b3d9e64dbdb9b73afa504f08d22058aa14967820a8c6d1311e65efcad6a63d56435304ba0da090ccf5056215173b13cf3c492156f2b2c5b5250afc8b4ab0ebeca9702a28abddeeceacdc20130d9acb00ce32176;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h891a7c1a3e6d0328a7e45ac23b32cbe1d9342fd844a6eb26d45f9a903ee29bc157282974a5118c3003c84010edef149abd9509c814fd1bff9eddfa5f7ff224b09b85a9a08a089e1bfeb1275f207073f88eb8d5588b897675c97ab8ebca244b925342b7de2a6c1409ca39880c3f33b4bc0dde804249d542c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157b91e9273c68638c5cde182d9b6b47ce7bcbded2703d8434d8ea9c4440198fbfbef41da51f5f5393982cfed7d8a4a6e6b28f6f61ead7564679d00e3b600d219abf417f29c909eaedd37cf3f9bba3cee3ba33b4e7864efaf1986d6b0ede4c7c98c26df8889b5189c1c1c959a9ec4da0ec644ecbe9c91af9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64d20ab8065146bbba6213f6a25c4c64b321dffef5d26768ab4dc4a6cfc4f32e047a2c762b2c73befd5b75c1ba813a86fa5467b70399fbdf3644972c8d6eb8e1e320182c7e1f5c33599a30b87b225fcbb41f1a28c0fb2c760f9376e3179910014029f0efddb5cff2284d66d0236a0edd9e9e859a4fe24249;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5aecb560059e21edebe4c84594d810599b3d60d738a2fa476b364be55d9ec5a7bfcc352ee16dfc8bd56abadc4c08a5c1ae9e62280ead152c38b10a3aa0b7600050ec3ccc2f944b2731cc763c2560c663f41f8d3727ed038dcfb6c6b81bd713f4471000938c7c8e843f8eecc2f38b06f3bc6c5cb09ca3987;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b1ad463f3080176272485e797f5d3ea5baa256847555e44588b6d44b5ecf98747b71d3beefbb7c3a6e0250e14d88dac4af0b47d218ab0cce721971989ea0a63b9748875ae9e75ebbbb4e6a74b151eca89e103de82dc02b910e6d9afa9a61218eb19ab8c1248656ca231130978a8eb200a8c13fa13c9f7636;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h838f95fc650d2f66a65a358a7b54a4228cc5b1e2b7d091f554aa179792dbd44a1113585a2d4e022b73fdbf51c042f681781d3c5c2e81987aa610dce31dcf25395256403d787a3fc1c02819c10aa706916f93061b27c543ec4f187f8b5e226938db0bc88ed4dc4f698f861c5e56a26aeba2ce67bdad936fe6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7c24484f65aacb64cad59157fcf9d28a15881a1cc76bef97acfdd0fb1a2d869aa0ec9a9b0667bdb0ddc54580aa3c6b530a1f259b69e65e1c57a2134b90d1141b130e7368791908d27f198a08a06286e3e2ed208c94de3f2532cc51bde7abf21519bd90cba569bd91a485dafbfecc150e219b9b9dea15bd4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a33c969381a1085cca2da7d2a733b9437d4c2b45825919443255b07fb9479d390d32b98fac7748dd4f3a31d077fed317a243372943281dbd8ad25d346425fecd123c34411d587a46ede0de1b14254686dbd2704301d2e5ce5d10735cb2582e78eee767c00b7ef133acd6ae52cbcc9406e05916aaf87b770;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h941b149446048bed05ea3cd63d68ab5a02d5255f62aff5853cbb5338682e9158b3b52dc8c3f0189f1e349f7eae7faffa00f8a53b4fcf708d53c33dce153114e34af5cb4a72c3a14181fe1d5ed4358aad59a7967bc4a055c95fa16be1d9997e48ce9affee8deb84b65bb87fae579a7207ac3717dda5fd6d1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d660a226be57a77a939eb920c839f57984561a8ab8603cd447ed341037158eef98fee197cf03768aeaa471f7524c6142c6c40b98b28984e23c2fc6d8a8c134dc1a1e9883f55246f15c57b37430b093bd242e4b90119809b40a2ce5b357192014ec9eb1c16353af3b89b1df8c0897eefeb4e5eee80d4a107;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4ec5819d784d781bf843a44b9edd6c38f9451dfda2bd4196a5c7c413e1e85a20f03f6b2314dc70d22f9e7eb9c18da7ceae7accb1f00781fbf8bc9d900be5493bd55eeb6e193a2967e1d1e70752f28f3f4d1c9f1a177484872219d8d53ca00a2fefef6a08063c2a866e147dbfdcf49e535ecfda423e35e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d5583f932aa09adc9896a9885ac7df6d2f0aaa34a24811f7a8eb38fbc10fa51d21ec79ccbcefe1caae67cffb4e34b38393d35030d60b6f35e2051c478e30a793a678939e113f830da345ab6fd7ebfcd31c3de2f17ebeefe75cf99530a8f7a9e96fb753998afdc42ff3b3cd2b4fbad5bb3a17f60d6a8df52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14067e1ab14d5f8d6fad6306e16b46b3ae87846f90475f82029a8a6fd30d9460cd911432a2ce09d2bef8cdb7ab5e86917aba2465c8aebb37710e80f2cd75701443efd153e393967b84d9e5fc63ee283549098c5dbc6c1d69f3a17ffbc631b041cbc9f717340e0e4541f04ca51a83db347deea24497189021;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha191964daa90438dfa0c455ac5e475c3c40db316f77249efc0ae3c1807052ee6402823839ecc9026590834b13cf109d11674d42acdc619c7a31506b266028430f06273fc4af86b2c8a1bd48614f3249042e8e017087885c8cbb69d662eacf3b868d7b8eb3d80aaf36c3f15e92f4a5e7a4152753acf4f7efa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf2a093d7eb18e40dad4e46ed1c3bac28f8ed26495546ed938a065fb9892a25d1bd5260ed2f0c9669943b56cec2373811f53bf87addf1ac392d3ef69efc541cd49666107a82bf5e4d8b127e08ecd78f4cd56951cceb57ac03c2c5bdec03eb48bc439adeceaa77d6452ca50ea8c02e2db6dfcc64f6c6a5d13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd41465bea812253fd79272d122da0fc2486242fff91a5efdba6067146f5af4a69b85b2ad5e6bfc07ab50d5e8bf4d52eca2104267a59682e601d9c6b9b8b88591d18099f511e5cb3476d4bf208bf0e757ac75a25869e270af58fbb7993e6b49bbb80ea91b363e7d0312572f6f4dc79dc75c9bde8ed2e9235;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b3cdd997ec24a626388d4be8f09a3b95cd9ddd243f58855d47611fd6a0cb621a084dba83d3476695c8a3149fe062cea37955dd3325089852834555bcb25f4333d4ccc4aedc8952e29b3137dfd5fc4f358f54e6e98e55300590d955e7a8bf8133bd7a68484c3c99a53f2d6c742e4343ddb4be8bd877c6dad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e61bb516a85ef8cfa5d523ab9bc484db89df4b7c1aeded15790819728ea3296fb4d9d8620d0db4e8268abdb5802be2dbc3db3193f829ee5784a03033c5b581cb263a394cfc628d061c33e6232bf0faf762dabdb94a3bb1ea272e2f8b8cee258c192aff70490a3909d689d27a536c31992fc89c68f6b825e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5067c7a0b8d77e6f09a5c10cf1de4c779ec564a317993de6423c2e62a41bde028746e5332a012e7a65fa44fc71ae8c2cc18a74cb8aa713c7a0420c42b67c1a5a6cde538cf6d481a3c622dad126984e78466c002c1554a302743d7a1b021725ec910f8eef9bdd2ae79ea5a7ee0510dbfd190e182a15a9469d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f724f6ea411cf21697bcd7ac9a9f364a8873b0fa1f8844c80b418aa8d6fd78ec83f45af02a5ae3b03dee98932b893e44a2ddca969baa5fc7b4b197df58c32377546c14081528ae345a45863643662943c42f338e4c9af46a0518429288a37c154374defc54f328d86693a38c9bb47d7ffd3d0c7490bf8ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117e9b8e2312ef4ab68d9cde8be8eb9ec6bb15435f84e6019d612801009bc00ecad7c8d895a053bef356aadb51a77fb1e6bd4e0c6f8522f64fe7c6ecf734bd82adc0725cc3a4a8d4f49cfa85fc4817905ed35808d988cedeb2c0049a4f6a7c8d31be9e5ee23fbdd44c86c73e31f73267ed7d970488598793e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9af7863cee09e177bdae4c848c0d00e758e962b7ff6129383c3cb3450e436b8d4f8fd049a44103611d978575bf905e15d94f6a5f4a3dc8f287b41b21157663100a93429c6575f46905765bdd39d407ef9a523a060b7aceddb1781c072445a132ff70a08cbcfae9236cf4bcfbda652677d426ad453ca290ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83fc8ecd43dbdc76daa9da40ded30c1d57adbae82a7797e182f3f9b244aa9f4ea601dcd34679a9e979be483d0d596265ac9f4b5b8fa25d297b6c70cfba46002bedac8345db81b31dfbb04d39e71ea3d3a6182c192dcca72e0495f109839749322da488b3d5689a0ad94281ffa8392d057aaab33262f4a372;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h969ecb2bff49451e3c297f1ca123ec834974d6b4d174580913c99482fc7a427e200af3a2cf077fec4b212d997982bde996a686aa991b421a62a5cdbdf1de9c59c35858c741b882b9b0f45b8aae3e0ed8b688bdb56d3586fd8c35f064d1b31a5e204e18b5c538467db68101f9a87ecebcfec0f743176a0e8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1852c4978a1017045eb41a07b51b6b0987e2e8c7ecfea93d6aab2f9ee3ff6900357111829e31fa5497fe33e6dd369111145456a05a8ed6011a06ea72fa6cca9cf99dfca585c0757c4d59edb4e04ee41f92a0c70a94fddd1d64af3e1c1f3c5587a90f0cf9187ed2c465bbb64e5355969f99120c6ac82bb16ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f932b3dbbddf8e29b44f418f8584de08c5c815c8c618dce70e5e5dbc3cc86aa36d622233f4361525fe940b31a0656c560442034ad52062b69856e2a668f4e621f0807ea977999a519392c3b7e9fd182d5ba4dfd1069a8646490fcdab96e1f9401f450c1470eadae086e4ece3e046539356d0c69616b9e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4bf57fbff77fb7c896580734227a836c77502b7f4b53707714323d2080d645fef5f61b41b5cd7551b644b811aeea1ff594fb6f714a6c1a81ef4a9ff292b9b55d27c09f3444c5c33cfe69b9ffb49e6be1629c1b809c024f78535d706e2c22acc017fa67cba2407a69a6aa77074633581bf919390e7c4bc78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3ef39fae661059f1691f2c38b8fc6f674d7f05f9bfb360d1097f71a906a54c99851e59d3b8dca0584c2e64aa24e4dda0a677f743a68cf794c3d0bc3d6622ad6a5975ca3af54b5928a3c7a3e19f20013f61bebd049c89d3d5b70ea4d663b3564c46a0d8095fd2ec937398cff41992e7418b2a6dcd6b4c116;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a546f1afc35cdcfea93753ddb59d92b153f7a9187525998576ad2c02e9a1d88b52e448fa737436d948d11d0b9f5ce0287e0c6223b675e743924c981eec60c3598fe0c67b2cad381045660c18c1db52c92b0aec84117ae4767ad265ffe903a00280ebac1146990ed526b5c8293153f134947a81ae6c25b10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102b50768cae2cbb15f7d06c2eea38ea2ff43d372635cbb399f23895ded61e5c656a81fef5a7c0c1eedc8791f3996aaa0aa998b74967ca86b13a49dd7dffbe72092280242452d4dec5d4afdbcd58c923e458c610f070263753646f3906a99eaa6e129ff4bd86f85b661cd1c64031fe227f8137a8da9acf76e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d19e627e5c4ccc98684ec54ebf549fe7fe2a3b54b75dbb6f31645ea708fd66a84a0037a4025dfe77992fa75314c94df8a6a5e8d3d1ccc4199bdf3ca887a4195e87aed91dd92a01b250d45639190c200fd1289fa7a81be74a23366eda3358c3e537557a27762a521c9c08826e8efe4d5734191177ef1a7b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18309322ca3e2faf064f3f76f9dea4b9e195495e24b995688694b5b268c5782fbe2dcbc5f5920bd19c8ef1e04bc61925d753a0f4b2519a57214afa60fcc1054187c8e0351e3f041e1e1fc2ea84ccf169efe3f301b0a9d7cd5d29a559026cb3776f06ea681ccd3ee8f12c7ae2165a074863d120309f952f659;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cfc9b25714033e25e5835118bb535bd9ac83034af69bac83c7ede8d993c4c8d060692b2de33090a93eac7f143ea8fd3f66c4c22c8a726509c0d06a60be0d6112d5a64b648badc53cd35a1fb6ae76cbaf41b80bc643114f5a74446ff98bf2e6f8929c0f3333e1bc73a85b69a7c02e43acffa18b490a1f4a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101f2b86466a3584b9c9e1288cdc3e3310ed4809c09bf8e7b37f4176727217ddee5164d252f96bffef66c4d0ba0e1c57fc30630c305fc146f20a66ab0c51aa238f7623f721d773faaaf62c8b729926102274bd23731a4a7022fa445043a4d867ccf5948663f58179b98c94c988914231848e569b4ae43b9f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he84189f71b864dea5ec1615bc422467deac6c8970bfa9758dc3e7758fd46f8ca6155358ef14fc7709c9482d8df3d6db4f1499fc25aaa9d67ae5abe0e195dbd5511b631c3c979baf650a8d063f970ba58b60f5e0e38b9cc3f5f4c58c807b54c766a33fed07cc9e2521e605be8ae9ef5573dee5790755fe785;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9eebf0bf07ebe357d6606b9109a9cf546eada0a1aa7ecda89c2753fa3ad5a866fdd2bf02d9ffee373a13040411ef9276bed9c9db74b47f67b90f0bbf6d3ba8b07db04f6d728cd77fbff18a75c395b1e7deb45512de89ae8fe20a357affdd565eb1ba0c8857b9b04c0bbf800c515151a9a704db8f0f2c7f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b063d1c492912f7d520069f8607a45be311e94105d844a69d8e8320a0c1a766c1ddcf54b23594814b1137c42ed6343c0417d4b338c7173f113a38a47bc78caf338ea18156113cc60b0362bcf1e3a27066cdecaec86a4a54df1555ba46a762a62a86d650269e5ad3e335a5e3330fa056e989b0a76ef063ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4390eee7048fb40b7ac33774af9daa4d5053fe7ea0f5b1f0642930c6b99ed5437b9f28b9ba1db0c7d69795b459186f9b339a3c4de0edb5ce550ccd27841875bb67098e4912f4fcf1265d66db3dbfb861e6a6d716788e81bab9591f66c27fad9c490685cd26ed856a41e552e180898a11c22bc57b06a1c8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74fe0f0d4df787e6cf00829cc263ef5bd0a3a7b9dc1bd43ade06a8bb4ff338b362d5cfedfe87ddc02807e5c1b3e62dac204605b614b6ab00737a061617a8af0710ff52549db2187313d815349f3cb441bc4ce7b03a9f2e4564890992901103f7b30dbc30b6518a8a1635223a9575eed587a0b911de67ca90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1762f06a479423a2d015985c134b28af17b0022eef8d60859aa2d3c8ab684ee0e0bd7b26a76b4b627323b7cc9739fafb9f5101c666925e6a5ea177cddb855d013610e7e6efbe5dcaaecd80ed401db69414b5a9260059ad82f74f5b51b98145c6696ceba44d79840696756f9005bbda9d50c1abacfd588509;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10afa0b5b77822fbfe5f570a38b5796b88d4bf257a00392b6731bf3ec32eaba381affee76d9efbde64d192258c94080364827d3487f8d44685a54bd4ca0605dc46f1a13a4006030fc871d71cd902ecb01d4c382f349d6180b7ec7dcd043991985c73110c0abb675ba82964f60a2ceacc415a2349f349546a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9cd1700480fff4567fdef9023f423c88d98b295b21f1dd7995824a1afbcf013f533d155cd9722d74c972cb77d7d22bd230226e1bb7aa643cea216941843b501d28e30b8d24b2ebf9f184f85ffb797ddbff3e2dfb062b20d5949132f093a1c33e181a928d9a428fa09f6c84318d31a5885bb0b78a00a97e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d321cd9c2a9fb2590ddcc30284b8d804116b6ca91ae9308bb0e767a9a5d6f034fc1f8c4dcfe16c2c8808e59a1a734b2bb8a09fb3a27f3b3a06c83cf2332d3c6f4784baab07e0b1e6581960f8ee8c02c7c2b991c32205e4bed467dacfa7bc099e8dc100902e806135fab6c35f00bffe9de54dff22c4cb22e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71d39c8a7907a1bb23d20d47945d4d94b441c0a0a6833a2e583bc21e585e1ba30d4508cbccc519c429263236a5479243b79a9ed45bf9b41690f63b65fadf309a9efaa174eb1bf0888497388dd25492382c1e5fbd5e25ec834fee99d173a5b0ba1aa28428aa3cd90b384d529da7786549deeb23168ec34695;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116f825e3c16d877f672d189b04fa1e0c1e37f08f46fb784f03cf33132209219803b12c4182d66439e38fb1a8d97a9b5270de51b87d70e7a2e331bc82a41838eef43bccc6fc2f891f1d39270e12a714bae924f6a6356b9294bcabfe4877001fc62f321f95428cfb6b0b0b27f2fbfc5eaf0a09adf53b040da6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9ebb884d8c82f875e7ba421258347e6227c035977d77fe2891f586e00812273bacfa167b34a7734c094f3625f8dc40b7aae18bd88bd0cf1690c508a29960c22a08d5b1f73420eb71a20b9a52ea8ccec1714aa89e53250f684a1f7ec2a61558a6c59c8b315b3dac5f2b402d553187c05f4a5947a490846241;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1870d77b7e96ef544a52c7d6952cc1d2cb4adf479b8b51df1fba777a5e6203906d389857bb456a819dbedbb57f80d70651942297e97b2f69d9550059587bfa2dbd789d51995e6ca4f40550c9ce082f1eed9ce8fae9887cd44a088d877978fd82ce436751df311ed6568aa5198562d7650709730214f1b6252;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14222e7f4504d1f37c3d45c00c499eb6843467f4b58d11351f822529c9282d37fe78a9b78fddc6da409134985b2a5ef5c334b104045e5ab87fffbe4bc248562c6b641df293cd499a0d9a5ff9d9b4bb674644d8ac400f0c46c98eed18dcc1c3dbe989f648d80fd3f95b9c033fee79f87c7a753830426c27d23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a274764e6aadcb59f4a35c5f59fdcfed1291185291ac4d8dbefb1a0f453e1467a9015d9ff052db88fde4ca61208b75987436227c1b3fb75e985d14cba232310d8862e5aa1146ad502dfe4adae8f523ab8b392bb184b7f12e8563a06655a2a4e039b009b0dc1821607696f40dd761d2fdd37c0b9cd9bde768;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7b3733c5b621305c1dfddc6a085de856775f3cd606be2c2f3e5e7e8a1f75abcbbd6493aa9d8ba51f05c833ef067218443a3b27c0ed675a3074e5c7769b3a16db90330039cdf1939eaf679e2eeb8df89bec63ac8c9d6005ae4e349388bf3274673fc7c10df67701bd7ecee73d0d6a44f36b0c096db9fd6c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc97231a868d7bfc67c9fa74ebec2078af891bdde788689abc29fee1cf5b27a9220e27327a91e83a00fcf8ecd25b806d501d599a84832f6be11f05486fd7ceb5e5487fb150a12ceb438e83e418a2884225943d8fc542415c2dadb92eafe9ca90d53f8ca8ea757f93af88db0adbd6ada45b84baf6eca2a2c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c81675d0d21b9dd76d62a453efc0e8c8727dd694849e7521ce99f14c048c59632a8d42c89a9c68f83d101ff682a62021e6527b073e58666857128d9c9cc96d1743d133fd36c74337e9ee8b94b82b0da29367ed17737efcc20ef4ad7ab1c2327827b74d2cbc4306c4136f2fdf2d3b94edbf94795ba4c46ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fba009bfd74af20bd53c7ca9791a62116ce86208686cac7ec20e7c817a7859cba58f3785c61603856653e98e1df1dbe73fde6defc7084ee434726abec05a689deaa9d42413661e1dcfcc35c39a96158209cb64d052aeb90ac25377003793b27df3ecdd67a55a135bc4c9d27da72dec2e3027362509912b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf1fe5b75378f108d61482d6fae5440614691dbb492d1067f6c3e9d69f1dd29bb031e440a71f996fe7705cc97d383c31a5267090942e4cb06a4aee469be80e6726e680d2c4e312ab63dc71f4261a49c742a33cd6ab108e7ec07f08e64cf2d57b8c5a3fd3214d647e70f7e5eaae03f02585684b1a07d4e25c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22272c8415c6dbb32337ccdf0b1352d108ba4420868f53ff83bb147899554cb4f8c1004b9b68242a7d66b4097dd8424bfd161b7fe4c20c70e800dcfcc247190b43b14be963721ec133de71c7f5ba03c772b07fec259587b9a94e4b35965c1539ee9ccb6f214b7378e19554d025d018b6eb0ae7731a884ba4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0625e0a98c1e5394aa6da3851b26f03c2ac3c6aa8a8c4d761ff15098959d6dbe888dabac01ef53a7f56ffffcbc61357b344cb80ce1e67ca73c996b48750a369b32eb7fb778532e597083f871ae9def6ac47a4264d2dcd59b22597580f657d16f1ac7eded31ba6bcca0479a1a4b9faea9f0162f277e7d0eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192ad8c82a31a3c6982adefc2bad28fe9f9ccbfd25405b21fd4647c8d064cdb00ed0d0cfdc127dd6f98077748d3620b0ba26a17b933ac1d743af83059ddacc33c82f5d95b2d242c8aff264e31e87a89211bded01678ed0ee31e8102b62d67d578a67864754cfdf9ad0d97e7ab2580d8986b22f0a4f0f37ebd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb791ec4e38f76fcf3de5c89aaf163e8f2b43cf70920b65976f34218f29165a8fd1e3dbe94703b4a8949ce9d5f076612600dac60e06a12e06a563c4b8245c2b86c7df7afe563eb53fb88d8503f227442bb68442605a8d15e24e439d42ee0aa7f18f360d41c91c6fcf139dfabb1c103b37274c0bc39b731c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ff6c639ab148d67a53535ee7da8586d5b55b2bc17d627cc6c2b68da642916e7a7478f2e3a25a945f375865c5b2275fbf88bbc8931c652eb1054dde357c61e714170baaf8745bb77ebdadca5c65deade7bf7174750176c944c5dffc9a33356d048e14074e61a4ba9f78da47fcfb77e891ea879902efbbdac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b844a3553f78d8d4f452c636738c2cb7ef5402a01b63c7855ef19cda6ce77d8e3abf7d4fa57a707e723164589e0b611a4fe0a86ed90d79f5faf74d8d2585e0b12d420109dd9223b98f12d1bafc60887e8956ddbe092f817cb68651488253240b7f356e34bba6e52d7d955a298b005286cd7c9c7dde398138;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h915b8338f8e564408f6a94b02873c29fe87e27a14e5a77c5749aa77dd3bd3cfad23e06cb1054a562347f68e3db43a4b526a58497b6703bc39115ad63861937fb08161f302662260ee33bc0c285c0d5f25fb54955ca9453392e729b3ccb5b1a1eb8ce7300b13193e4b29e70c635f478ad4298213ca51fb351;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d0b2d16fd40ff87885f3495e618a30c3bad995e05ba647d5eedb95be803aef99ff30040342e3bed877ab85a13be03a8019e80683bb2b93146f7735e69b1f1747016199e8f3c68429eb6bccd556568a335640104b64b9d767920527fd218aef99aca6b57ac87ea9eb5c27bbc3d0909322522aeb0b916e610;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105f0e90a4a3f845740c752dd601709d3c2066b82787d35f111fd28fff02d085f67cafc61f12b8b356ea7107200d7d1f6379edfcaf99c578ccd90c60252b09d992088633ea2b3ca164b2ffc0443351407211f416ca3aeb9f94897de84594027533119b043b0a2f4d0f113ac35c199f13bac32ee50d487a19f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18dfaaec2fe6839c9657d299fb3336bf6cc6f4fd9e9f7a4efafbd64a619caf6bc34466e9cb33faee276d730bd1c647fe8a33cdc47f2c98b15b9cb5b07a13a4a4a7e37e7e6e9ee92fde3a69ee80eddb108ac0cfa7477ca8f94dc42aa05fcf66d343f894e6deaf226e91c0e2a8349f035d3fb30e3c8da303012;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114342600a264f88d6fc3267d8dadc1d150753dc7c6ba012580e0c5715f9dad8ebd6d2d784e50fb11dc793d988f2c79d028295ae11ed26bffa4078fb3ff91b5fb062643f211590c2fc88fbc2cd98db5c2814aa932bad7b235811f038d7225a5a49ab8b2dc58efb7cba17856afeb43acb6ef01d2effb4b83cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d925fbdc05d980d28a3336320a4fcc5c27bf72b35466f73c4dc5a17640420b0eba60dd78ad7e016afccfd048fd7a66c82457cb91ba09acf644eb536a64e1613771f85f4116d4f4d95c7a911b648fe9c3fbbdf98dd0bcba4e0b1364a82fb184da19516cf076e93d2a45976eb0c76d1d2e4794d27b2b38ad4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c410a18d04cfb0eda4996438838e942932d7b62683598e83da8f1dc5a9659ec543bde27f34b814030f2473caceaceac314cf0c3e453c70fb2228fc8759cc858a913f36a03b159638459e1b96dfdfccd1203d5a8afc3e20927727b0083f56a8481e8d8c5cf6dd00349b54cce9f72c8ac733864d7c211f6e80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d80b5d754faf51962d883fc741a31982825d22a2bc2bbac27062974d6fba50914c9b8f182e4db4c3b40a580ec9bf35f75b9a52de9758087af6dd950e23c195387123a923a795289f6d5e248d7c228a7bc68af28014ff9eb9fa17b4938c9a666133a89b5c835befb1dd7d415bab2a2bdc8df7f691367f1d04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1067f54e7eb56b4e6d66ddda77b9048eb033c451e43e1f6d3a319f483d6f291de8497300d07185ce758f414bf624a57d4694a251f831366ced5df81c522a3bce6e7ccb70449e272492a8209fbf57e931525aa21d34e1243145e9c62dbbba6a637f0106a222210ca46e5be5366d11b1d81d757f9cadd7b71f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadfaae950720d38c9f608c0c236ff57a486605c2ea5265893f6daff0b6d8703958a5fcf149aafc2721d08a7a30d006e471e21602ee43e6daad89e5de7d09e6330888de9a329d95c132e8551914267265a9ee72be9ae846d73ca9dd79dac34d73e59867030d4b8a27a5e500a853bec869591730bfc4e13d13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8108c769a6d96b99a13466dbfd7eea75424d58985927caf669267a79f8c37a0cdc333fddc63fde98672581bed3d2dda6a91d3fe77284113586ffc6410c92c81d129c0608ea43b3c59197bcb8512f67403cc3104d0df9442db9fa2f26ded261c2c3d2b64f3a067798e5085bdf3647d7748d648067c7ee3d27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d02125a854d685bd857b4fe1ee6d9f9401e0a1b1ff956d06eb01715ccbe4126e7af01eea446e7bfc167fd68e7f8a2f08d040fe6268bbf1d648c3175e2c0140ea36ab3ac631d318e3a5d3d1a43e791eb2f1200328e8e68110bf8d97616ca4c4ba952c0806ca8ff94afee4901cd02e683f99d052802d36637;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117541d1c216c89599f1ce0ff46ab063f995058d1058d627506524345fb2cc73af5cfa583848300ddaed6e639deebd0c40a66ec4a827d23d5ad9a0d1f5a3d1911fe365ebd5418f237504b208c5ba00da8c0aeb8e69318cc3e0dc8d15aaa9d3997399f96881c85341a219820793dea727de1660b9cfd3b2585;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199bd9693038f72ee60390c1931a52cd892fa3f455307aebd0c654d69347f9942af577e3232880c072d7c01d1528dabf53d6a9a7878b471079177f186c074db57bfed09e72d03b8f73e901efad6cdb78147f2327ff84544b891f7a64597caaf174019ad00e1c21805ac5b469d7b9235a5a59c69a42f96cd32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h993f40506d7b17db216c04d839464cc12a70b8551a99999563425369ff5082756d9f88360e716415baaa57d9dbe7e8fce8e6cb29d7563e323c00f3ec50076c45328bb127909dde85515929e8fd43eab21f505473cb1e1b74764286b1306401fd04fe3e2a4d83f507d5d6035d1f8967fa64a019ba81fe9e12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfd7b702b08758b3a0b7af1d710625df6a11aaf553ef8b8df4d367f8925339ed2eb8bcf3780f6b5c2c37461078907ab4e46b76734f66be6a5eb6a2202316701a7b5458cad191901f5161c5b7d77542fb2b099eea9eec88a73663e5deb50f18c5a0de924c6660f141d9789a746b3e8544afc2e038c00f962d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2f5abcc00cf2bf0934ff55156d2068ca7f04c0b6644808a619df9ed385eac5a16ea14051cdbb07e75de463514bdb340ce5023dc6aa8d6c7cb0788de916cfdbdee3129a81a891b9d100a2df4e69d60a18df8bbea76ca28fe6278accdd67aa0729afad7f5feda0c9ca2f56fdba177693b351738e08789285;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d812313d92786e6a93fb3371908bf7c14be7fb184a0c60876cc08e71d4f969c84ef16f7cc143d06f6aaed55fd454fd9ee797b576ff76a9951bc6f82d898e9ef8c5afe1d43e370b4777e594d4126360b71dffe982dc2e714c8dae64a2dcef1a76993bc819cde0cc83da69fee4a528f3bf774ae69cc5d9b355;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fed1edd72d0c6a8eb1ba315b026532377853af9dfc9ebb57f6e50d2c418daa2150a54fa9f0a87245ea9c63ba03c11b6f7123e950cbd8ee0f06338bada163a22d8c8f076f74ab5ca22408691c4304dfcd08835ee442df4cb5397ed6e5400c672fa0cc1f072612b84e1dba3e8d00df7578bbc3beffab1a567;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160819d26c9d4402a31f492c02e4fe5d7f11298d748327c9e138b32cf73019de4ffad30d00312fb3a4258e9ae3f7efe70b72fdd47d39a4e3ebb70cdf4e64561d27ba4cbf10c344a04b49354bcc0859b8ec13d00c918a8be3f4f0a515e52079edb93c6598c9e150346169069552eaf06c27dbcbafe6d24c036;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d8c4ef789bc47e16ad0edae0926636ea9ee495d3eca7c816dd647a965a02a2d5d789f4bb7cbba74d7383e91cd41420714f1b780183efcbb98b776aebe85735ddef34441e437f3d7dd1ddf70b94b9118faee803bf56679d50eac8b86cc312acbdcb765d7b8a38a675a4af67b8a44086ce49a4cfc6e52c1f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a8335828edc5964cb417aa3490979ddc6f21c2eea346da48400ab6944bbe940684034f1360ccdec0dc04ddb3666ef9976b85091488f3e0b97199b079c5857d2addeeafefe4b6fff23ed162d66f5ab9fa69a0e192763145ec59c11e3780a5fcb98fdb43da088c71c329a461f9bd450e62c0645070b6a911;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h936a15cc601678459edfb668a69e559c0e897ab7164c7ce45986539bf19d9a901edb986156dfb2403e1947c85d10f451be6dee0bd7444f55604e956c790fec400222ac4d49751c472c964c33ace27baed9da69914c435d556e2d762a4a8da5f651a0f7852b8c207e7fe20f4df2ee049eb389b1e262ecc2c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120d2d716b25af542b98ee8f2952afa3b97ac7bc59be05d02c6e382a716daa59b6e7439f9995ec104e6014dcd4ee21234b80a2d18fb67edc276814a30c887a477f323062e30d473ba72092842f3f289a903732f03c7abf95cfa271e3036935e66635874100be4643a9981a22f2fb66196cb3ebf5208e5b8c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb669a6bb72054e26a73a014621c2f321a0c1b1d1ea3cc0322cc7d91fb7ec25eb6c53afb214380f97531d93e7493d6e74994e97ab160858b88474bdfe84f17c5797216a91e3e71b438e29b9a41fa7846a1024f554e8ae20f9f6984a2c105d1d5027ca7714881668f0618fd1af1a697203635e35952b7d9fe9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79c717993d0f19abbfc48d251e03c417ab8f2aaf5766e82b2a2106688ac9e839a774842396244d0c9f9e57feebdeb18958187c1deb2f9ed157f41dd65fab0acb219977d0c6c07f753224522e074fb9eb65d791e19bfbbae287e60f6b9e7f1ebc63435d04fdfd22cb795dfec8ebb2ac08670d8dccd4c13034;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f652ed810b3d608ab7d7974091931ed6d6eb19177f11458727faa7ca8e1e7ec64659d0e0cc2591b52a751571d9952a540ce8174b5629cc20283d8f940fa5edd439e2708e442c32145d09efaf82601d96349e2ba6ca6982f89c38df1b86a74084a5252614993c4100645a674e283f42f17dac28f956e8145;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a2675bac3a6529ce764b429cc30d3502fb1614360eb76e8f733098b137d4d559f428a1c2dea423f4a452082bd7842b77cfe38ce0804c42247a751b19ba2f1c462ba4d1eeb57fc556876418554487e07d7c9b652e972846fadd589b1b21ce862dcceefd57c6415537cc0bc8f0cf5c702caada6d476e0a6cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75d55c471009f127ba29ae627aa5441f38ebdbf0d8c348b8e7b08330bc89387dbf5735b9663a14d4f58cfe2bdbd71c063e6d775830191f793a4c13a3e983e03f0ed9c7de5e3f2348c93e7a4fc7fd52b23f469879fb09b69a48a74b490b97576bf0f173c7bf822fc8d7b9873f4359b15d00e6b2bc80d759a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a53fa97286f2c3f2fb934acfaf454803da2bae81eb7ae8f5aadc35ec50b0fe8b0c1bffc822a6cec2547d19f145031891783b80cbc2427dd9a9eb29e4914d62a55127afea4c015dd8917b50c96a44dfbd3768c1c0b27906607239a29fe0f36baf9409cbbd50ca36024cf2ff2e0f2eaa246c169e5df7d7062;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had5100d090c07f8a158324adb0a5a086fade2da2675971c60458d5d7c4a35df40a0ca7a79bf146e084ae41b8a8587c2eec3e544c2d14fcf4c25de2507cc7811d26bd1ce69a5505bdc763bbb8bb5c5260672236b7570fcdd85e3ff1ef979cde4431ea754726b36b24921eb75c216a968e9f6403c24a950981;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8763038904ab6b7b7ab4260155f3c2381d673e320e0146556a457b71ea261850ad6add058fe2d1f74d50a7e7f433aa5115209bcce4163cbb43d5bdb81340eb09cdb82b7c71b4c8616426dfb6c7a72ea787bccad5bbf8106f3363df7121587d48e3b9b40ab016f1b67a500c436d487c6daef453bf0b3dac18;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4e60eac22315c6ecea64b4dfce9c15779b107d2e5e9193af3e536af17e6ac11034bc065ef5e9452f4d74539f937618198fe334c1201ef431f72665313c7b1b1a71dcc40b396b89f3f43f7a1e111f66ed100b4292a2285868eee66680431a3dea98d8f3c48db2bae7a65555514abb17baeb81781892e8347;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc086407afc4daf284693723d0ecc0726314cceebfbf44af01a8632e798b7edd39c444eb19269db7c806f98115dd5112951c16dc4c1a1923bc87dc21c2a0e721d3ec211e5e4612c897cac6318843e6ef0e5fff3857c8edcc66ebaf730acfb6981c32e0e63db35a5839153407aea3e1a75106b2b259709bfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c870bc09fe0e7757f642437a2bae574ad09013150f29c73dcff0fb2cb70051fb30f686dfc7422e767e593c7145340f50e261acb6a63f136b5c1a13c92464d7363451c0b795a64b451f973776e39f3635af92586600ff702a2bc41276277777abac50716712a45786c9abc555cef57621a2cc9aaf50877dfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h278ca93c719ad053fe879053146a88b0db54511051d503965a67ed0fc8cd9ca8f540fc0f67584cd106fcaec874ade99792145d96aae3131cea19692afb2a238c3b9c2972389b1f61c35d88f3c71513342320c61c93074bb50f41edc939fa988528039181f045927f704b467d3e88c49728fe6648c87574b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19bb24d7195d4de9aef6752218cbf67a60c210478c00c6dc5532cee2a1b1334e2c9a53da9274bc6a1702d182f070dd39445fa91dde3a2a1870e138bfb6781d9fcbc4ca56d9ae302539e6e72f4fbdf18135189431917978683b99bdb64fd70ea1b8c40aa3eafb4062df9a6bfc6d0e82d059faa8329bbc59829;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41f20d5e1a0b309047f2522f91deb11e1b39764d8662667760f47d114fe83a4995c5b3b4425d444cfcf521cc13653ffbf68e5ae62f5f3a9449ae747433d1a9e907d9cfb9db5f2b563f6095675ad557db6b7e75a3368babe589cbcf061242555efb1c80424f9884ae8e23c5211bd3a43d7c6f07483cc598f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he521eb690a3a45fecbfb81d85f8c4dc9b2a865866550d0d7ae931605a9c63c43380718e369e164b66fb8a069c85dd66d5cc0754eed3ba78494ba31e63a04dbcfcf282a15aac97020fc010e0b3e446597aa238e3678aebdab546aa903ab87019ae4b5e5e6418da283003c5a5119c060d2162940e1b84ce26a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95e69440ce4bd62541b5de3075153ad9f65d232672b15163b6657e6904f9d5c218f74b33925c653bce3b81a8d5269f337fa8b5eaaad9fd150fbc6af08aeb9164f7731162b33572cc006e26eff05ec398945e5e23d319ee5ccb12f6052e3b3897fec1a4d759574cb89d3824bd0aaf64d665acf4c34c521251;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33f3861cfff31d61c336f5b1aa505cc89bd4600fc5c30668dc5078a2ad58149a275a55b5c2c9685c06484c8c7ae6ead0d684c4c931386fed6cbd5e15e8412545ffda4bcf38eb91a6e0ec6ac41dc9bbcc2dbe395adcb13d3315e05ebbd2a77f85fd351e8ee0f717aa650b01a07bd66aadbc64a375c1a600d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5a32f9289f79ce0bf481f79870917c4aae521a8cba6e967043eeb3611481430b5c98a48fb025f45e81f5ae4917f8ad31653368038a9f4c0c1f5b58e93a7d4197c7fad2b83ae53aba7cb45fc01625db03ac4362fad610f1095fcad47c944808e71df3efe8ab273a4ea033cb8ad89a01aea3d9e32d8b7efb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdc4a191639c159d0d8ad041de185cdf83d5b311309d98a9d01a3b585ec2c37fc1cf94d63fbf6d2931fac5633177b440f34341f22501392bed75d8a627f8a8b9b002023c6635a2be892ba3397a80623a11aeaa8e223f35908876b9dce9ebc01b27b34e47d4488d18ede590c4181ddda3776c245140515c21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18afa7c21afce0c480f7342b7f16d94d535766a834b82ef92c4fe4f4c8c69357e616804a2858b6d19af229c9c910eb7ea0ee3b76d61d4fe69f1a5295161ee02a986c00d717707fea1c828288365e046a53e1f2e0ef6b449120694f4b86c643341f5fd74e518b36f9aa1dbc70d135bbf993e22eeb060c3aa03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12adf796b1bd04927c83854735f147d84130b788cfe48f7b06553bde2f25ef2d170f3aed430c927a3680152f6a5b6a96b9528f29b759b1cbaa6f05d8828224e31f26e007f30a62a6c25507ea798a35cdda67cd917b9dfd6b18bbf2df77db8dbbd1c2e4a7602d37199ebfd1c61a23a29d6e6290878cd0a5240;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d60b074d1ea497abbfa8e1689923989f2be306b860de8b08cf2fe57a6c7742f0f8b1e289cfe738e8847f1b207a1efb6305ba887b520027ad7e59f7dd1ece0c5d8d92ef74d7b3feee660d8037b1c25f9a009883b61547e8b8bb83f7e3e1ea36fec441cd1159743f8664db51235ca058a95fe499242058fc0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b5a529eb702098231f6bed00eb7a8b35c8dd196f42332b5152d62c93c91137604ec19a5d0ac33bf38420f025a0e77a3a85d556088875cf37bfe7b4f6736a5691375669e8dc4ca54f9a1e0a393da90c0f75ae56ce0d8fe1f0cd5c0f885fbb3e3f67b5e1deff276aa42c60ee87b1878e5245f2140dcd8d267;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d45e683a057f01b616c5e9cdb5086c32f2d9b1599d12861b135788c1ae17189112edf197ac2521a2e1b92f5cdf550ea479dc189003f51e4cf90b923fca946db82d58a3b98841a63cebdfc56ae293dd9e1cb6c1d334c7b28ecb16e59cd64a4a8f9abb0436d6607ebed369eaddbe7ea1ca36da08cf73a10af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4456caf74bb7af4aaaea336efadc1a43d577e9e968d27ed2b2eb9a736586621474f2e67c901f59a06049b30e0d981b9e38e65e5398646f36a3965dddf155aead90f0b59fdac3aceff6cd3915d7d22a4a50666afd778a15e781cb6cb4c1730dedcccad4d9b396354e467862e0c5cabee4946d11700e2f5a52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd37973545bb1a3e136c636b4aff921621164f6c76537066391f5cb85fe1ae39aedd84814ddf5e6a1d7efd48f475bac25f406a8ca22b4789f62f61a96eec2a71b7aecae75303f4d5e4cf544cccfd7b36f27dde36f0253b598a9769ea0977a6fd4ce299fd6b268492c991982dfbbbc66e2cc461534496f4aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cc8f789a7e9776c826736f817c3226edd3916fef06a71062dd50ff314af9ae197629a7d2cdc31fa3b5dee1c07aafdb3f0c504b01002252fc4f23b8bca3d4dc88adfcb8e3f68c73c7c6a95bef9e270671cb6600fc48de54e120e2cf118af54f22cc85a859e995941df1a6cb67283484b820629c0b965ccbc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dfc9998eee59598086b81d556610af70d442368b08bc71a3e1ba784523a40b4da1ff6d5a735a3cc0ed8965215070fe4a3ec998614068df90af9f3b27addd80acb3012acd0efcd46d66de357654e15a243b0a4041e7789855a76086d3b42cee7651cea11fce09dcadd9933979306b04d27dd8fc4c0d2d7c52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0c7d28e81919ef8273424e417fdda4af18ce077a5746401cca8a8257c5d8d4ba4653414c70030ee22cf254354c93a164654325f14effc20af8d17adf1750e55736744c3abc6f525a50252651507a8acecfc326a70659697c55cea3d8e0e976af723d9895a4e038fa8ff27edfeec33f5ccae64ffaaa1823e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1441d2269168d18d7171c775f1c08a21e10f19941a334ae0f939cb7e6da2c534f3dc4d1bff246d67915c80c82aacb97ce92e7ba082b29a3cc1781b4b0eab7889f2bb3045dbdaa94012f7cdf063edd109c5be81ae40f5de865e83d24b44f1a51a426369cda7dc46cef95edc322dc685eae4672906518ae2eb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e34b262a938c49f5d76a63b5f53f0182652b4a367119f0483ac1efa99f9a8f91b6989bcdc8fd1b56de45729f048fb20bbaa079e351434c8811ce9b4ac1449f6453419f1e0dd4dcb9150100aff0aeb6f16eb07fcda3a669c164838ca6392ccd0913784518271c2efed6bb28d2839df97404553f309a3d7e29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h823bc7496cc2477c5194234bd3ce227d92299451c8537940d4086f095737a714c28bf27ccd98f099cac6aea7535b3eee2fdfd721ea2712f126baec851831e668df6e6cebb232f78dc9916753376114b231649b7e35877b9764935465cd38e4c81f07fda024e3b178476d420f61971d88fa715e62da758bdc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f36c6bf4844400c33f3f4ca42cac80ffa543cdba07e81a5dfdd5af7ec8d0efe9ef56d25bc475a8c74bbc9f0e99c7eea7cb4b123cb913d8d5b7e634340b95faf000a2c51f9d490bcfad5d576df80b37def45e6febe3d138060bd3aae19f5917cefac292f10f9354baf6b34d05d6e69112703600468f9f2db3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4b0166909355f073b6049efa0b530e522a9f7232a585b9e60e7421bc6bf344f430ec5d3d7542e1e41429cfaf349889da49f539e67f28e9bde1a4ace73d42d2b76c9b68ff0b5e09b2d09c1db8d8c76c0c32b0ec7bbc5805ba52c37a73be6fc67018e8e1b08b225b00425d07c5bd35f7ffdad59208354925f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcee8a12c9c588a1d7309f3394b70c0bda9e256e2cba1e1e40aa8f426d6700c927c495a8f515b379ff8f8091bea41e8c3237ccedb9e9fc3e180f59bbc3010093ea11283c8db5489869f62254e8df11173773e2067d4023b50584bacb07cc23733dbf3e595751b5011209a502f8eefed8f1d2c0cd0aaf633cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf19be407f045053957b02f8fc5eb28918f1e4738c51e3305235edd3073b12a69feae6c1224a4fe987c67d7a4ae8b922c6cc8a0a3b76b06359053cb44e94a3839861b4d0a250b1e8b05d32df8092f8c791eb46062d0fa5efb48d526b2755ba517c30d4a0a3c307f921bc531a06833108eb4e6a795f19ef249;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f5206b2535ee3a492a2fd8557b65340cd814a43822e4a3deb96dd775355b0582b153827008b40487911968e8367cb799772c137e29c94bd7e3d3e4978f8bffd4e4eef9c19d041cb3a186e655a55851ceebeae9e889d16dc248611ddf2162cc6430833f995adc51a6d93c015bb623f2a0af0fdf2b03a5023;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b860f5b209a8495ce28bdc7da6deb18445f59b5d395376509910702956aef25802c1714a1efc5dff73f1f1a00b332abe5090eab6323b3db4e8d244a21654604e64f4708f77b336e1520e53641e6f0ceee5c3777e6c279b62179b34bb9294a018899be55922e4bc24deff91787a23a08a7fed34cab9fe9bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac92e721e2e0854baf67ee158911462ae7b3cf96ceeddef5f2f39d6c8cad138709febe0c30fb8cf960732a7716024959e29b19daabd7731c433d704c69b0b1e1a6c58deeaac074cd2c5de4eb72319f690621e8c7068db99113378adfa8db87af55156f03e8c187736acc3ca5d11a2a2870afbcfaa33e9408;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbd9165d2691bd40952145e4ccfe2bf0b455003f8b26ac5d312c3ffa041913e4fea8be82060cf094f35e41353fee8d0322fc6784422a66d827d4ffe9822ec6b9b63147997754d06e5a5b511df51972e237e94a2d34c1dc578bb223e9f1babc358b31b697928312dc447e85d736e6f0d6729ba005f6304871;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e81ec1128ac9089b29e046c1a14349a17b5c0431f407d4fbb5ff13b40209576b646f87ff761db1a516e9b41cf8c6b97bfff3cfc6a1183fc8dc290e4e4494d15442cfe5998dbb514f23896d56c8cb74f05f955f01a97aa04d3488b5cb43c7f753bcb2f9a51f8baf5a4109016fbc9907b6163ffcb6659f5a09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0e9f9bb307094a277b69f820aed69feaf8e43037186ecc481bdfdb608dc44c759ffced00d5495e45e1fb1a94b1289efa0861f19bfc1026cb55bada929d6fdab7acb77b20e91f852f314d388c0d1994172f3280bab61163d25c4b15c09f7185a02b2048707727dd40154481a53f15f9f5f2a202408e21262;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12cb2d9898c673c074b12d4e110d83ce0f60f75be9a5b31e9a5b5ecdf68346bfcd2ffc5c8c6da2c13a02ef01f4f53d1bac68cc6cc097a7333c076d889a04c1355c81a989a20adc6e06db38cb68a3520aa9248298b60ccf0951e00e18efd7f54ed064d2fcd96411a718ff55e79ceee3863e3bad076b4bedf37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d6d0bf78852a260a92dfb9d919170487c22b2a77bafb4c06b5482b59b4c33255b7e603f8586ac26c82b863052a76387c9165565e7f2f5fd7ba6696f44dbbe67c936c06ebcd9130b571ee6a4e8f5501abfd36f5e20afdce1e14178c396bb7709500f12362802cf5d360a75abd0081ae51eafadba01ac9dbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b242232b2604074d560d7bcd7385a4d36a7fe851bb62cf7cf458275f801f9fbcfea0ab17308550368d9324be75b436d302aac32a661652626cf7efb39d61a679b354e1d65f0a325f459cfb05ad36e2e9e202138a69af63b7ae60e0a7ace98d0e74338c35e95dde5cfe25bae8a1e6bf42e8c1bef60ddc5945;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he98dbe93ccb8451691113b5a703df4aa684e5c543e5faf7e3641e076772b5ec7fbe42a1b9a70cf0c6f529deb101f655be8010fe67d28d4696e730c9d9fa20a02a4da36b7358993865684eb01dc6aed03856287e96fcc9aa3b5f2de42b4dd42703d5459f91908f55decd3feeb63cdd58092666fa44430333b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84ffb5ea944dc97f3207a0236edae64fd495fc653bd62f1ffd352c857b6eebe3cd0e58925bd313154b18e21459d21ad6c87a3b826e4e4132749d9085ebcd442592a9c3a40fbfca1b4aa97d88daece85f20101f05c6ad4f030e6c650a055f332c15c9e1eb984f7016c05987d06c77a900a8e0f6cc3cc9593e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25bbec24e02f80a19bffe959953866406ad53034f55da0c1b8acc8e5febc7140ea5a141c80e5fd55a76d8ad24ed75aff1805088ffea959cbf34cc4c6e546d8c7efa3fb0610255c3a81bf4c1f5cc4aa79df7ec98ace9b986d02b8a23ffb36761ac4e667cff9c1a8731809071e0eb6f88e4d83827ea20acd3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b06e0a02125022b7e3c8086ad740f30cab824f8501fa84bc28bf65402755636b3eb6fdafbe9dcad211e19169329d9ab0d9578fdc49d2b922189c1cd06e154d8d5d5309846c03e0b34da39a190ac5db3d6a099035b6b17fde1f2249c5aecd68d94c36c6daf90766647e7d9ff025fb637fe6d46a651bf8183;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db138150a1d246f3d2273457bc0d4367764db0bf6b62c79c48e11151823702411cbb8018e98cf638f364b9ff891b2c59bbc529f3112903ac23f181abf4f53da8a07ee34226dca0295ab5175edb88a2887f3cd39017f3d66c76182f12d30e7907d228cce28420ed4edbeef26b54dd3a167707217bb886ec9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f9c37471e631b439258d7739b80b3f04fbd29f440da666d582e183e67e58711cac6c04a1e3e5fc34dc200d56eeb0276200b9dd32fecac91f20131c4aae67da87d6a44bd67be323d85b1ecd1a3662c48bae046da78729052f1747caba6f5d284d24ac7d4586cac46fb435b71828317c1e4a73a1ad39c2c56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h350f62bab2d946c02257769a06169e8056a13aad3010a892ce2b23ba835048db031963d5f171204bcb4d4cc176cb607c3a6fe109006f3ff83f8dc60c8cd2ec892601db0bc7b13c73052c03024411598d75e27d4e2d38fef7b3b6fe09e4c78d29652b3a9238c4dd90635ccd90ef09aa32afc841f18afac10d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1932348afdcd5f4e9de37720b9c0dc4e6c5ed0a0c89a1d9a7b52a81d3bc3cd2c02e0d7c341a85b6edb0ee822759e9be9dcfb810c420e4f69162e3a6883adf0cf3001dca22182a9b3cc58da21f3efe1e1e5720b7aa8fd89e20601ff95f7a6c681dcb965c860e379513725d704f6541e68bb0ff2f90f1e2c3ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19872423753d7d55b040c5e003e1a0acf8fd73d5e79854aa15517e0916ef59bc3bb4fdb68527d6b3d4c44d13418fb90453585d09b75f9d10e2046e52179e1b5a02de051ed69c97d0685806b246e55071c0c4acfb4fefe33ed25b42c02337deada5d81f86076c55b006baa279d956903a67da5426a78fbf38a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1522f053669a0d276397ce437693eee9f8b289794a9c6b6e62a43243931b6891476462140a8cc8724c77e2a6554967213fa5df7fffea8ddd46c2a02607c0c9ed0017c0e1a6dcc17512e0422447c1b7b548dc9029432b5db89c0eafe3c23dea36260b857777c6bf9aeba1a2f69d08bc0a72ab7ab4325c58e43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44f9074b8b1df3ec8333accff34573967157574502f310327167cc75a41420f3061cb4653a2cde93998fe77bd4c060b98dfccb5925a22159c06a94d2904f26b68f534ba761d7af58f7d7f7281a54c332490d8863ebcbf5c9157140c6a5bc2a12b91c3ae36d96742b3d8ac7f92ffbf8bcb4a91d361cb0a323;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce3559249f9243a1473c40cf5a7b6393a2865916774ef06d87474eee6b30ea1a2881124b71a1992ccccfef30b2b9ca93512d4e587a8d0e84908efe040f03f5f86139f1e355322a0c788891a21b99cc8dbd9df406351727b35315c118a173b9df3a97d4851d9ea0eb10089bcb4567a684de2ae27f04ffc5a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cb64f83da242aae017c87b8ba523dda50113e3eb07457415bdfcb859aeeb28494a8dcfbba04d28f107f4139a3247321aea0a6ee16ea03a58c73993eda55cf6c6ebe4dd3e386179883b4ddba6e6f1a696d92c30badd1fea798fb7a78323a2535de96957c31bcdfb947560d097bf106bd38660aa36d34a9e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16504859026a570de9471c07300fe34845acabc42abf3d96908de503458a740eb0beb46e0e19e816ba55a0cfc86aa784491c6ec93bb55ab2c9f386e38e9eca7935b1d4cb3e3e81b2bd1befd51d7ecce0bd6de5fc6baf66e4b5b5a2c4be629627e5c3240232605b5ffef644da496ece210f0355e61480c9e26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5895a7b6e27e4c982742f5b9a1a809af3d100eda2e4da93c8233094176f6845a5ab0d6234ed7e9c0ba72d70f6d9b468c798c5c5a53a723c37f673b4aa577daa2d62f20a6b0d8ddcd81502cbd9715c8df3d47fd0d25e47ba9bd47053ee90da0ce05ab11728cfbb09a43557b0a8dd0fd754e5b05484ec8fd3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h931150565aec8a3cc5b243fdaa8b01fe383c7220bdb6a7c9144403443ea53b21953a79e08170baa4a5913ade504b2c1ba91a8de253e2cc095dc0a30081891a25e998d33ec96715f4a23ab73903c3776a67b6fd2d22fd4e5084950545244bdd880dd40138950400cefd68fa8e5e9c09eccbb4ab3e93651141;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he09bdc88d6792b584dd5a40765b1779ec2777ca5c3b3dd0ce3f7023edd91a7178018133447d3f8c1394f7bd635d21ae22453840a7cafc12fe2a0d7279f0136babe90afd02eaa669dd9d2db7c039bc21c11e484b8a1f27a243b168497bbc38b65d1f192ed830f55ac19231de8fab432db3946fa043b66229b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adbf0fa5ec42c8342f29d58a8744e5942ff505d29385771ca5b02caac028aabe57d4ef3bd865c8ccff6ea26f5e4d95e1581ae3e124887d6c0b0b10779f304811a767979cff7800a44f761c6086ca16e41b1c84a118fb65c1e0ad506da6ae0e68a31436f0d3dc6f155a577ee24b93efd551026de8c1000971;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cd965f8fe9981920f328d8dafae0e8743cecef832dfed500ed498116454c51a0317bf93d24abef08b1497e6487b3c8314f99145e234b68d72bcb905b074e5bd69de93d31f158a28e9dade1b44d97cd2ce2ce72b157fcf6b37dff12cc1fc26ca19b62510e1b0d1fd7a39d730aae8eb44af2f5f196f3c02a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a125e035aef566af57ed7c49c319e721d28a1870999ba8d4f96944a0557d297aded4a3157d1be115e336a8973c590d2a18a0d554465badd3ba50b6305a5214db28ce12127a789525c5c0005856f29f8a9abb33831bb54c899ef4d6853c2d23f44ba3c63fe8493bd1f329920f2dea122e99b87a969bf313f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176c93f21e0fdf7ea185ea66e069a5934b590050a9359132f94ab33bb0545c2862bbf50460786d11244022dc20d16b4e7f73d2a65542daf6e17bc8b57b5f0f19ff6a1bcbf5ffc9124047e480e01c1ef36a9decbc4eed60a0b57e0405d153199faf6fe7fca60fb4acc132ddc792cf5abf92c1a57d330e586bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf438581e1be93c837a0e935bd08f8873b84afc6a1bf4ad11d6b4fe151ff031d3464b5662b2d4189deddfc8385012a635e657e7670c5dcd7bab618dd26b88097384cc10269c2ca37bdd0c6da9c641355bd175862d193d02f9a81a82176d22798fc50ea805c5595c855739704964b5850df4ddb7241c4dfec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h714f9c6932015db5f63dafd463e0ec209513d9a1640ae76c7195f346b3b9670a5d4fa21394367537565b7b9aac2e6cd851547c4bcca9128abecc9e6c58ef0c488f0eb3c5fc6771e1e2cceeb515def7c8e150a4b4dd7552994b5500673078b2466893d0fe0d65ea3287de56593c3b17ce8d8a3c70a10dda0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f8aa49807593bca0f8ac41e3ee9ba7794d200dfb7fc885e6c21354e13a73a6a344c54ed95fa51e2cdc7c642ecbf99710000557501160e05aad65aef55fa00be5b99a67d7d2460f338e14eba8300df5c067b37482ceea3fd88a671df39f43012f81160480725b1095474c4ed187ec6cde3dddc4a1b1cdb98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19753c254df719f08700720f37af132e540dcb74329a8eb031c979c471784e42786a22221294be47d49f87b52f3a452f57f0ed1bfa0f027edfada07e185a443baea25be5f700a978ace8e9cdfd812f12e9acb1d69e31cc15b22086d35beec30e3a30ce6399c715291447533a83474f1f65b69c3c6027db3a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd0654c5e458237216fc834eec578e7accb133911e630ea2761e120664b1f99caf70f5a7f5bb4c304c02f08c6a831cb661118a30ffb435ae2a5c6bff95b3459f7c9a7b0781eb6901714848d5dc8e16006e4c1aafee24dd350bcc069d963489c516af0ae17bb0d90e43fc5249ecbe2d66e70069049a873c99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c84101c9788c0b80a44dcd084793ecfd7e21bf04c4e206a7a17b4835ac9c178c8e8ec9bb1c8cee5b84591a99ef23028e5a20bdd1844a23944a923a9806a2c27aa832fbdead2e10b9e8b784cea35ba88bd160e7183febd042acf0688feea3ffeaf9d9ad3158cd454ba5c605baa2e2233cb931913a2ad8a22b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f44b42cb35ce5b78c6156ecb7f27ec2ceef0a64963973d479ac3a657ee7988a9ff7ca5ffaa55e89d6153f4eb5615b7c84e25a20c6973d29bf7e88ed37e2a9b1e7156981be38bc51d330dbecf0b7a387b4c5400206e30135b32a6b9160694cd06de58d6ed9d0a7aa28e3e7449dc5873500c45c2ce05f0b73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23a0696eec86ebba135a225d7770478a9d095cfec6516bb426881e2e1bf7ce5c35a14c6e59569951b05d3591978e4c2aa59805ba5568b0286df9ec81979885498cc869e23a4efb28b441005bd9092ced94edf9be56d409e69891638efdf58d6e7d5426855b75aba931a2b5d918d2d4cd9de9a2d5025eec0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f28255b5128194fceaf93115cb4b7f3c8548f55d95248e444061b2b2d88a98261743299ae921c54377904502e8a46c528412208470ca803484c45d906bfe13d3fc31f2e34e51d4728831391e29f611d9de94f38d2a43599d636c39dede5533ea61cef101ea2e45cc933b761e8b0a48206e9b568114200b09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a143692dabf3c65492cb23d05f71eacb30a03194e811c12fd7da3803685d6ed07baa63c423b761ba7b6ae1a0b97ac1cf23859623ce829ff167f3c5146894c08dc53bc6890344378c0cccb7342c66d2d02836803a070f078dd07819471a91f45f3cdd2aed9d51850891248f23d1db2a3e59d84c1c215d73cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd6b1673251089d7163ca751370b102469559eb2f156790459d22d77708308cec4ea1a3f7513af6b52415ab800e322dfe75274f599f17764af8435cc314899381a37066b3ba518a23ea62d33ff0622ca811a21f4763ccdc9f008a6a062d0485794a3576f262fcccd481977752a357630bff88b9a613a01d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d90e45ed5543bd34ef4f0e6791d148d6b7fa3d82aa330148d97a3a06afd557eee96e420e5d969eb7a652ea27bb2601198eb02bced488ef299d5040b0f8b842b71b6cd998c582d231a60bd6eb2f0c43c67a9f60bc67aed754efe197b39ceaa67903cd95083e517baf9e44cea3b5c51cb1037d2417d9c0dc3;
        #1
        $finish();
    end
endmodule
