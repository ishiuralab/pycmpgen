module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    compressor_CLA64_16 compressor_CLA64_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA64_16(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [0:0] comp_out20;
    wire [0:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [19:0] stage1_0;
   wire [29:0] stage1_1;
   wire [23:0] stage1_2;
   wire [26:0] stage1_3;
   wire [39:0] stage1_4;
   wire [28:0] stage1_5;
   wire [26:0] stage1_6;
   wire [22:0] stage1_7;
   wire [28:0] stage1_8;
   wire [29:0] stage1_9;
   wire [27:0] stage1_10;
   wire [23:0] stage1_11;
   wire [29:0] stage1_12;
   wire [32:0] stage1_13;
   wire [24:0] stage1_14;
   wire [23:0] stage1_15;
   wire [18:0] stage1_16;
   wire [9:0] stage1_17;
   wire [3:0] stage2_0;
   wire [21:0] stage2_1;
   wire [7:0] stage2_2;
   wire [10:0] stage2_3;
   wire [15:0] stage2_4;
   wire [17:0] stage2_5;
   wire [11:0] stage2_6;
   wire [11:0] stage2_7;
   wire [15:0] stage2_8;
   wire [7:0] stage2_9;
   wire [12:0] stage2_10;
   wire [17:0] stage2_11;
   wire [7:0] stage2_12;
   wire [18:0] stage2_13;
   wire [23:0] stage2_14;
   wire [7:0] stage2_15;
   wire [12:0] stage2_16;
   wire [5:0] stage2_17;
   wire [3:0] stage2_18;
   wire [1:0] stage2_19;
   wire [1:0] stage3_0;
   wire [6:0] stage3_1;
   wire [3:0] stage3_2;
   wire [6:0] stage3_3;
   wire [5:0] stage3_4;
   wire [9:0] stage3_5;
   wire [4:0] stage3_6;
   wire [3:0] stage3_7;
   wire [7:0] stage3_8;
   wire [6:0] stage3_9;
   wire [2:0] stage3_10;
   wire [6:0] stage3_11;
   wire [6:0] stage3_12;
   wire [4:0] stage3_13;
   wire [13:0] stage3_14;
   wire [6:0] stage3_15;
   wire [4:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [2:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [5:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [3:0] stage4_8;
   wire [3:0] stage4_9;
   wire [3:0] stage4_10;
   wire [1:0] stage4_11;
   wire [2:0] stage4_12;
   wire [2:0] stage4_13;
   wire [8:0] stage4_14;
   wire [2:0] stage4_15;
   wire [2:0] stage4_16;
   wire [3:0] stage4_17;
   wire [1:0] stage4_18;
   wire [3:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [0:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[50]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc615_5 gpc18 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[51]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[9],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[13],stage1_4[22]}
   );
   gpc615_5 gpc23 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_5[6]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[14],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[7]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[15],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_5[8]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[16],stage1_4[25]}
   );
   gpc615_5 gpc26 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50]},
      {stage0_5[9]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[12],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[13],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[14],stage1_5[22]}
   );
   gpc606_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[15],stage1_5[23]}
   );
   gpc606_5 gpc33 (
      {stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc34 (
      {stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[17],stage1_5[25]}
   );
   gpc615_5 gpc35 (
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_6[43]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[18],stage1_5[26]}
   );
   gpc615_5 gpc36 (
      {stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[19]}
   );
   gpc615_5 gpc37 (
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[17],stage1_7[18],stage1_6[20]}
   );
   gpc615_5 gpc38 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[18],stage1_7[19],stage1_6[21]}
   );
   gpc615_5 gpc39 (
      {stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[12],stage1_8[19],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[4],stage1_9[13],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[5],stage1_9[14],stage1_8[21]}
   );
   gpc606_5 gpc42 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[6],stage1_9[15],stage1_8[22]}
   );
   gpc606_5 gpc43 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[7],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc44 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_9[6]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[8],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc45 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_9[7]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[9],stage1_9[18],stage1_8[25]}
   );
   gpc615_5 gpc46 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_9[8]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[10],stage1_9[19],stage1_8[26]}
   );
   gpc615_5 gpc47 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62]},
      {stage0_9[9]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[11],stage1_9[20],stage1_8[27]}
   );
   gpc606_5 gpc48 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc52 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc53 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[17],stage1_9[26]}
   );
   gpc606_5 gpc54 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[18],stage1_9[27]}
   );
   gpc606_5 gpc55 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[19],stage1_9[28]}
   );
   gpc606_5 gpc56 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[16],stage1_11[17],stage1_10[20],stage1_9[29]}
   );
   gpc606_5 gpc57 (
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[17],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc58 (
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58]},
      {stage0_11[54]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[18],stage1_11[19],stage1_10[22]}
   );
   gpc606_5 gpc59 (
      {stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[11],stage1_12[19],stage1_11[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[3],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc61 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[4],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc62 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[5],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc63 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[6],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc64 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[7],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc65 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[8],stage1_13[17],stage1_12[25]}
   );
   gpc615_5 gpc66 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_13[6]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[9],stage1_13[18],stage1_12[26]}
   );
   gpc615_5 gpc67 (
      {stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage0_13[7]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[10],stage1_13[19],stage1_12[27]}
   );
   gpc615_5 gpc68 (
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_13[8]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[11],stage1_13[20],stage1_12[28]}
   );
   gpc606_5 gpc69 (
      {stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[12],stage1_13[21]}
   );
   gpc606_5 gpc70 (
      {stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[13],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[14],stage1_13[23]}
   );
   gpc615_5 gpc72 (
      {stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage0_14[54]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[15],stage1_13[24]}
   );
   gpc615_5 gpc73 (
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36]},
      {stage0_14[55]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[16],stage1_13[25]}
   );
   gpc615_5 gpc74 (
      {stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_14[56]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[17],stage1_13[26]}
   );
   gpc615_5 gpc75 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_14[57]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[18],stage1_13[27]}
   );
   gpc615_5 gpc76 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage0_14[58]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[19],stage1_13[28]}
   );
   gpc615_5 gpc77 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56]},
      {stage0_14[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[17],stage1_15[18],stage1_14[20],stage1_13[29]}
   );
   gpc615_5 gpc78 (
      {stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_14[60]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[18],stage1_15[19],stage1_14[21],stage1_13[30]}
   );
   gpc1_1 gpc79 (
      {stage0_0[53]},
      {stage1_0[9]}
   );
   gpc1_1 gpc80 (
      {stage0_0[54]},
      {stage1_0[10]}
   );
   gpc1_1 gpc81 (
      {stage0_0[55]},
      {stage1_0[11]}
   );
   gpc1_1 gpc82 (
      {stage0_0[56]},
      {stage1_0[12]}
   );
   gpc1_1 gpc83 (
      {stage0_0[57]},
      {stage1_0[13]}
   );
   gpc1_1 gpc84 (
      {stage0_0[58]},
      {stage1_0[14]}
   );
   gpc1_1 gpc85 (
      {stage0_0[59]},
      {stage1_0[15]}
   );
   gpc1_1 gpc86 (
      {stage0_0[60]},
      {stage1_0[16]}
   );
   gpc1_1 gpc87 (
      {stage0_0[61]},
      {stage1_0[17]}
   );
   gpc1_1 gpc88 (
      {stage0_0[62]},
      {stage1_0[18]}
   );
   gpc1_1 gpc89 (
      {stage0_0[63]},
      {stage1_0[19]}
   );
   gpc1_1 gpc90 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc91 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc92 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc93 (
      {stage0_1[54]},
      {stage1_1[20]}
   );
   gpc1_1 gpc94 (
      {stage0_1[55]},
      {stage1_1[21]}
   );
   gpc1_1 gpc95 (
      {stage0_1[56]},
      {stage1_1[22]}
   );
   gpc1_1 gpc96 (
      {stage0_1[57]},
      {stage1_1[23]}
   );
   gpc1_1 gpc97 (
      {stage0_1[58]},
      {stage1_1[24]}
   );
   gpc1_1 gpc98 (
      {stage0_1[59]},
      {stage1_1[25]}
   );
   gpc1_1 gpc99 (
      {stage0_1[60]},
      {stage1_1[26]}
   );
   gpc1_1 gpc100 (
      {stage0_1[61]},
      {stage1_1[27]}
   );
   gpc1_1 gpc101 (
      {stage0_1[62]},
      {stage1_1[28]}
   );
   gpc1_1 gpc102 (
      {stage0_1[63]},
      {stage1_1[29]}
   );
   gpc1_1 gpc103 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc104 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc105 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc106 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc107 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc108 (
      {stage0_3[57]},
      {stage1_3[20]}
   );
   gpc1_1 gpc109 (
      {stage0_3[58]},
      {stage1_3[21]}
   );
   gpc1_1 gpc110 (
      {stage0_3[59]},
      {stage1_3[22]}
   );
   gpc1_1 gpc111 (
      {stage0_3[60]},
      {stage1_3[23]}
   );
   gpc1_1 gpc112 (
      {stage0_3[61]},
      {stage1_3[24]}
   );
   gpc1_1 gpc113 (
      {stage0_3[62]},
      {stage1_3[25]}
   );
   gpc1_1 gpc114 (
      {stage0_3[63]},
      {stage1_3[26]}
   );
   gpc1_1 gpc115 (
      {stage0_4[51]},
      {stage1_4[27]}
   );
   gpc1_1 gpc116 (
      {stage0_4[52]},
      {stage1_4[28]}
   );
   gpc1_1 gpc117 (
      {stage0_4[53]},
      {stage1_4[29]}
   );
   gpc1_1 gpc118 (
      {stage0_4[54]},
      {stage1_4[30]}
   );
   gpc1_1 gpc119 (
      {stage0_4[55]},
      {stage1_4[31]}
   );
   gpc1_1 gpc120 (
      {stage0_4[56]},
      {stage1_4[32]}
   );
   gpc1_1 gpc121 (
      {stage0_4[57]},
      {stage1_4[33]}
   );
   gpc1_1 gpc122 (
      {stage0_4[58]},
      {stage1_4[34]}
   );
   gpc1_1 gpc123 (
      {stage0_4[59]},
      {stage1_4[35]}
   );
   gpc1_1 gpc124 (
      {stage0_4[60]},
      {stage1_4[36]}
   );
   gpc1_1 gpc125 (
      {stage0_4[61]},
      {stage1_4[37]}
   );
   gpc1_1 gpc126 (
      {stage0_4[62]},
      {stage1_4[38]}
   );
   gpc1_1 gpc127 (
      {stage0_4[63]},
      {stage1_4[39]}
   );
   gpc1_1 gpc128 (
      {stage0_5[62]},
      {stage1_5[27]}
   );
   gpc1_1 gpc129 (
      {stage0_5[63]},
      {stage1_5[28]}
   );
   gpc1_1 gpc130 (
      {stage0_6[59]},
      {stage1_6[22]}
   );
   gpc1_1 gpc131 (
      {stage0_6[60]},
      {stage1_6[23]}
   );
   gpc1_1 gpc132 (
      {stage0_6[61]},
      {stage1_6[24]}
   );
   gpc1_1 gpc133 (
      {stage0_6[62]},
      {stage1_6[25]}
   );
   gpc1_1 gpc134 (
      {stage0_6[63]},
      {stage1_6[26]}
   );
   gpc1_1 gpc135 (
      {stage0_7[62]},
      {stage1_7[21]}
   );
   gpc1_1 gpc136 (
      {stage0_7[63]},
      {stage1_7[22]}
   );
   gpc1_1 gpc137 (
      {stage0_8[63]},
      {stage1_8[28]}
   );
   gpc1_1 gpc138 (
      {stage0_10[59]},
      {stage1_10[23]}
   );
   gpc1_1 gpc139 (
      {stage0_10[60]},
      {stage1_10[24]}
   );
   gpc1_1 gpc140 (
      {stage0_10[61]},
      {stage1_10[25]}
   );
   gpc1_1 gpc141 (
      {stage0_10[62]},
      {stage1_10[26]}
   );
   gpc1_1 gpc142 (
      {stage0_10[63]},
      {stage1_10[27]}
   );
   gpc1_1 gpc143 (
      {stage0_11[61]},
      {stage1_11[21]}
   );
   gpc1_1 gpc144 (
      {stage0_11[62]},
      {stage1_11[22]}
   );
   gpc1_1 gpc145 (
      {stage0_11[63]},
      {stage1_11[23]}
   );
   gpc1_1 gpc146 (
      {stage0_12[63]},
      {stage1_12[29]}
   );
   gpc1_1 gpc147 (
      {stage0_13[62]},
      {stage1_13[31]}
   );
   gpc1_1 gpc148 (
      {stage0_13[63]},
      {stage1_13[32]}
   );
   gpc1_1 gpc149 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc150 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc151 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc152 (
      {stage0_15[60]},
      {stage1_15[20]}
   );
   gpc1_1 gpc153 (
      {stage0_15[61]},
      {stage1_15[21]}
   );
   gpc1_1 gpc154 (
      {stage0_15[62]},
      {stage1_15[22]}
   );
   gpc1_1 gpc155 (
      {stage0_15[63]},
      {stage1_15[23]}
   );
   gpc2135_5 gpc156 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc157 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc158 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc159 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc160 (
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_3[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc161 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage1_3[9]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc162 (
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_3[10]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc163 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[11]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc164 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[4],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc165 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[25]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[5],stage2_5[5],stage2_4[9],stage2_3[9]}
   );
   gpc615_5 gpc166 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[26]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[6],stage2_5[6],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc167 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31]},
      {stage1_5[18]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[7],stage2_5[7],stage2_4[11]}
   );
   gpc615_5 gpc168 (
      {stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36]},
      {stage1_5[19]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[8],stage2_5[8],stage2_4[12]}
   );
   gpc615_5 gpc169 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[0]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[5],stage2_6[9]}
   );
   gpc615_5 gpc170 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[1]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[6],stage2_6[10]}
   );
   gpc615_5 gpc171 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[2]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[4],stage2_7[7],stage2_6[11]}
   );
   gpc615_5 gpc172 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[3],stage2_8[5],stage2_7[8]}
   );
   gpc615_5 gpc173 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[4],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc174 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[5],stage2_8[7],stage2_7[10]}
   );
   gpc615_5 gpc175 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[6],stage2_8[8],stage2_7[11]}
   );
   gpc606_5 gpc176 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[4],stage2_10[7],stage2_9[7]}
   );
   gpc606_5 gpc177 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc178 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc179 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[7],stage2_10[10]}
   );
   gpc606_5 gpc180 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[8],stage2_10[11]}
   );
   gpc606_5 gpc181 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], 1'b0, 1'b0},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[9],stage2_10[12]}
   );
   gpc606_5 gpc182 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[10]}
   );
   gpc606_5 gpc183 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[11]}
   );
   gpc606_5 gpc184 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[2],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc185 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[3],stage2_14[8],stage2_13[9]}
   );
   gpc606_5 gpc186 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[4],stage2_14[9]}
   );
   gpc606_5 gpc187 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[5],stage2_14[10]}
   );
   gpc606_5 gpc188 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[6]}
   );
   gpc606_5 gpc189 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], 1'b0, 1'b0},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[7]}
   );
   gpc1_1 gpc190 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc191 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc192 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc193 (
      {stage1_1[15]},
      {stage2_1[7]}
   );
   gpc1_1 gpc194 (
      {stage1_1[16]},
      {stage2_1[8]}
   );
   gpc1_1 gpc195 (
      {stage1_1[17]},
      {stage2_1[9]}
   );
   gpc1_1 gpc196 (
      {stage1_1[18]},
      {stage2_1[10]}
   );
   gpc1_1 gpc197 (
      {stage1_1[19]},
      {stage2_1[11]}
   );
   gpc1_1 gpc198 (
      {stage1_1[20]},
      {stage2_1[12]}
   );
   gpc1_1 gpc199 (
      {stage1_1[21]},
      {stage2_1[13]}
   );
   gpc1_1 gpc200 (
      {stage1_1[22]},
      {stage2_1[14]}
   );
   gpc1_1 gpc201 (
      {stage1_1[23]},
      {stage2_1[15]}
   );
   gpc1_1 gpc202 (
      {stage1_1[24]},
      {stage2_1[16]}
   );
   gpc1_1 gpc203 (
      {stage1_1[25]},
      {stage2_1[17]}
   );
   gpc1_1 gpc204 (
      {stage1_1[26]},
      {stage2_1[18]}
   );
   gpc1_1 gpc205 (
      {stage1_1[27]},
      {stage2_1[19]}
   );
   gpc1_1 gpc206 (
      {stage1_1[28]},
      {stage2_1[20]}
   );
   gpc1_1 gpc207 (
      {stage1_1[29]},
      {stage2_1[21]}
   );
   gpc1_1 gpc208 (
      {stage1_4[37]},
      {stage2_4[13]}
   );
   gpc1_1 gpc209 (
      {stage1_4[38]},
      {stage2_4[14]}
   );
   gpc1_1 gpc210 (
      {stage1_4[39]},
      {stage2_4[15]}
   );
   gpc1_1 gpc211 (
      {stage1_5[20]},
      {stage2_5[9]}
   );
   gpc1_1 gpc212 (
      {stage1_5[21]},
      {stage2_5[10]}
   );
   gpc1_1 gpc213 (
      {stage1_5[22]},
      {stage2_5[11]}
   );
   gpc1_1 gpc214 (
      {stage1_5[23]},
      {stage2_5[12]}
   );
   gpc1_1 gpc215 (
      {stage1_5[24]},
      {stage2_5[13]}
   );
   gpc1_1 gpc216 (
      {stage1_5[25]},
      {stage2_5[14]}
   );
   gpc1_1 gpc217 (
      {stage1_5[26]},
      {stage2_5[15]}
   );
   gpc1_1 gpc218 (
      {stage1_5[27]},
      {stage2_5[16]}
   );
   gpc1_1 gpc219 (
      {stage1_5[28]},
      {stage2_5[17]}
   );
   gpc1_1 gpc220 (
      {stage1_8[22]},
      {stage2_8[9]}
   );
   gpc1_1 gpc221 (
      {stage1_8[23]},
      {stage2_8[10]}
   );
   gpc1_1 gpc222 (
      {stage1_8[24]},
      {stage2_8[11]}
   );
   gpc1_1 gpc223 (
      {stage1_8[25]},
      {stage2_8[12]}
   );
   gpc1_1 gpc224 (
      {stage1_8[26]},
      {stage2_8[13]}
   );
   gpc1_1 gpc225 (
      {stage1_8[27]},
      {stage2_8[14]}
   );
   gpc1_1 gpc226 (
      {stage1_8[28]},
      {stage2_8[15]}
   );
   gpc1_1 gpc227 (
      {stage1_11[18]},
      {stage2_11[12]}
   );
   gpc1_1 gpc228 (
      {stage1_11[19]},
      {stage2_11[13]}
   );
   gpc1_1 gpc229 (
      {stage1_11[20]},
      {stage2_11[14]}
   );
   gpc1_1 gpc230 (
      {stage1_11[21]},
      {stage2_11[15]}
   );
   gpc1_1 gpc231 (
      {stage1_11[22]},
      {stage2_11[16]}
   );
   gpc1_1 gpc232 (
      {stage1_11[23]},
      {stage2_11[17]}
   );
   gpc1_1 gpc233 (
      {stage1_13[24]},
      {stage2_13[10]}
   );
   gpc1_1 gpc234 (
      {stage1_13[25]},
      {stage2_13[11]}
   );
   gpc1_1 gpc235 (
      {stage1_13[26]},
      {stage2_13[12]}
   );
   gpc1_1 gpc236 (
      {stage1_13[27]},
      {stage2_13[13]}
   );
   gpc1_1 gpc237 (
      {stage1_13[28]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[29]},
      {stage2_13[15]}
   );
   gpc1_1 gpc239 (
      {stage1_13[30]},
      {stage2_13[16]}
   );
   gpc1_1 gpc240 (
      {stage1_13[31]},
      {stage2_13[17]}
   );
   gpc1_1 gpc241 (
      {stage1_13[32]},
      {stage2_13[18]}
   );
   gpc1_1 gpc242 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc243 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc244 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc245 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc246 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc247 (
      {stage1_14[17]},
      {stage2_14[16]}
   );
   gpc1_1 gpc248 (
      {stage1_14[18]},
      {stage2_14[17]}
   );
   gpc1_1 gpc249 (
      {stage1_14[19]},
      {stage2_14[18]}
   );
   gpc1_1 gpc250 (
      {stage1_14[20]},
      {stage2_14[19]}
   );
   gpc1_1 gpc251 (
      {stage1_14[21]},
      {stage2_14[20]}
   );
   gpc1_1 gpc252 (
      {stage1_14[22]},
      {stage2_14[21]}
   );
   gpc1_1 gpc253 (
      {stage1_14[23]},
      {stage2_14[22]}
   );
   gpc1_1 gpc254 (
      {stage1_14[24]},
      {stage2_14[23]}
   );
   gpc1_1 gpc255 (
      {stage1_16[12]},
      {stage2_16[6]}
   );
   gpc1_1 gpc256 (
      {stage1_16[13]},
      {stage2_16[7]}
   );
   gpc1_1 gpc257 (
      {stage1_16[14]},
      {stage2_16[8]}
   );
   gpc1_1 gpc258 (
      {stage1_16[15]},
      {stage2_16[9]}
   );
   gpc1_1 gpc259 (
      {stage1_16[16]},
      {stage2_16[10]}
   );
   gpc1_1 gpc260 (
      {stage1_16[17]},
      {stage2_16[11]}
   );
   gpc1_1 gpc261 (
      {stage1_16[18]},
      {stage2_16[12]}
   );
   gpc1163_5 gpc262 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc263 (
      {stage2_0[3], 1'b0, 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc264 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc265 (
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc266 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[0]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4]}
   );
   gpc615_5 gpc267 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[1]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5]}
   );
   gpc606_5 gpc268 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[4]}
   );
   gpc606_5 gpc269 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12], stage2_5[13]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[5]}
   );
   gpc1163_5 gpc270 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[0]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[2],stage3_8[4]}
   );
   gpc606_5 gpc271 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7], stage2_8[8]},
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc272 (
      {stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14]},
      {stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc273 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[3]}
   );
   gpc615_5 gpc274 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[4]}
   );
   gpc615_5 gpc275 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[5]}
   );
   gpc606_5 gpc276 (
      {stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6]}
   );
   gpc615_5 gpc277 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[4],stage3_14[4]}
   );
   gpc615_5 gpc278 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[5],stage3_14[5]}
   );
   gpc606_5 gpc279 (
      {stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[6]}
   );
   gpc1_1 gpc280 (
      {stage2_1[18]},
      {stage3_1[3]}
   );
   gpc1_1 gpc281 (
      {stage2_1[19]},
      {stage3_1[4]}
   );
   gpc1_1 gpc282 (
      {stage2_1[20]},
      {stage3_1[5]}
   );
   gpc1_1 gpc283 (
      {stage2_1[21]},
      {stage3_1[6]}
   );
   gpc1_1 gpc284 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc285 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc286 (
      {stage2_3[10]},
      {stage3_3[6]}
   );
   gpc1_1 gpc287 (
      {stage2_5[14]},
      {stage3_5[6]}
   );
   gpc1_1 gpc288 (
      {stage2_5[15]},
      {stage3_5[7]}
   );
   gpc1_1 gpc289 (
      {stage2_5[16]},
      {stage3_5[8]}
   );
   gpc1_1 gpc290 (
      {stage2_5[17]},
      {stage3_5[9]}
   );
   gpc1_1 gpc291 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc292 (
      {stage2_9[6]},
      {stage3_9[5]}
   );
   gpc1_1 gpc293 (
      {stage2_9[7]},
      {stage3_9[6]}
   );
   gpc1_1 gpc294 (
      {stage2_11[17]},
      {stage3_11[6]}
   );
   gpc1_1 gpc295 (
      {stage2_13[18]},
      {stage3_13[4]}
   );
   gpc1_1 gpc296 (
      {stage2_14[16]},
      {stage3_14[6]}
   );
   gpc1_1 gpc297 (
      {stage2_14[17]},
      {stage3_14[7]}
   );
   gpc1_1 gpc298 (
      {stage2_14[18]},
      {stage3_14[8]}
   );
   gpc1_1 gpc299 (
      {stage2_14[19]},
      {stage3_14[9]}
   );
   gpc1_1 gpc300 (
      {stage2_14[20]},
      {stage3_14[10]}
   );
   gpc1_1 gpc301 (
      {stage2_14[21]},
      {stage3_14[11]}
   );
   gpc1_1 gpc302 (
      {stage2_14[22]},
      {stage3_14[12]}
   );
   gpc1_1 gpc303 (
      {stage2_14[23]},
      {stage3_14[13]}
   );
   gpc1_1 gpc304 (
      {stage2_16[12]},
      {stage3_16[4]}
   );
   gpc1_1 gpc305 (
      {stage2_18[0]},
      {stage3_18[3]}
   );
   gpc1_1 gpc306 (
      {stage2_18[1]},
      {stage3_18[4]}
   );
   gpc1_1 gpc307 (
      {stage2_18[2]},
      {stage3_18[5]}
   );
   gpc1_1 gpc308 (
      {stage2_18[3]},
      {stage3_18[6]}
   );
   gpc1_1 gpc309 (
      {stage2_19[0]},
      {stage3_19[1]}
   );
   gpc1_1 gpc310 (
      {stage2_19[1]},
      {stage3_19[2]}
   );
   gpc606_5 gpc311 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc312 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], 1'b0},
      {stage3_3[6]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc207_4 gpc313 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[2]}
   );
   gpc615_5 gpc314 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2]}
   );
   gpc615_5 gpc315 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc606_5 gpc316 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc615_5 gpc317 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4]},
      {stage3_14[6]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc318 (
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[2]}
   );
   gpc1_1 gpc319 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc320 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc321 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc322 (
      {stage3_5[7]},
      {stage4_5[3]}
   );
   gpc1_1 gpc323 (
      {stage3_5[8]},
      {stage4_5[4]}
   );
   gpc1_1 gpc324 (
      {stage3_5[9]},
      {stage4_5[5]}
   );
   gpc1_1 gpc325 (
      {stage3_7[3]},
      {stage4_7[2]}
   );
   gpc1_1 gpc326 (
      {stage3_8[6]},
      {stage4_8[2]}
   );
   gpc1_1 gpc327 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc328 (
      {stage3_9[5]},
      {stage4_9[2]}
   );
   gpc1_1 gpc329 (
      {stage3_9[6]},
      {stage4_9[3]}
   );
   gpc1_1 gpc330 (
      {stage3_10[1]},
      {stage4_10[2]}
   );
   gpc1_1 gpc331 (
      {stage3_10[2]},
      {stage4_10[3]}
   );
   gpc1_1 gpc332 (
      {stage3_11[6]},
      {stage4_11[1]}
   );
   gpc1_1 gpc333 (
      {stage3_12[6]},
      {stage4_12[2]}
   );
   gpc1_1 gpc334 (
      {stage3_14[7]},
      {stage4_14[2]}
   );
   gpc1_1 gpc335 (
      {stage3_14[8]},
      {stage4_14[3]}
   );
   gpc1_1 gpc336 (
      {stage3_14[9]},
      {stage4_14[4]}
   );
   gpc1_1 gpc337 (
      {stage3_14[10]},
      {stage4_14[5]}
   );
   gpc1_1 gpc338 (
      {stage3_14[11]},
      {stage4_14[6]}
   );
   gpc1_1 gpc339 (
      {stage3_14[12]},
      {stage4_14[7]}
   );
   gpc1_1 gpc340 (
      {stage3_14[13]},
      {stage4_14[8]}
   );
   gpc1_1 gpc341 (
      {stage3_15[6]},
      {stage4_15[2]}
   );
   gpc1_1 gpc342 (
      {stage3_17[1]},
      {stage4_17[2]}
   );
   gpc1_1 gpc343 (
      {stage3_17[2]},
      {stage4_17[3]}
   );
   gpc1_1 gpc344 (
      {stage3_18[6]},
      {stage4_18[1]}
   );
   gpc1_1 gpc345 (
      {stage3_19[0]},
      {stage4_19[1]}
   );
   gpc1_1 gpc346 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc347 (
      {stage3_19[2]},
      {stage4_19[3]}
   );
   gpc1325_5 gpc348 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0], stage4_6[1]},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0]}
   );
   gpc1343_5 gpc349 (
      {stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc623_5 gpc350 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc1343_5 gpc351 (
      {stage4_14[6], stage4_14[7], stage4_14[8]},
      {stage4_15[0], stage4_15[1], stage4_15[2], 1'b0},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc352 (
      {stage4_17[1], stage4_17[2], stage4_17[3]},
      {stage4_18[0], stage4_18[1]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3]},
      {stage4_20[0]},
      {stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1]}
   );
   gpc1_1 gpc353 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc354 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc355 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc356 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc357 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc358 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc359 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc360 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc361 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc362 (
      {stage4_4[1]},
      {stage5_4[1]}
   );
   gpc1_1 gpc363 (
      {stage4_5[5]},
      {stage5_5[1]}
   );
   gpc1_1 gpc364 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc365 (
      {stage4_10[3]},
      {stage5_10[1]}
   );
   gpc1_1 gpc366 (
      {stage4_11[1]},
      {stage5_11[1]}
   );
   gpc1_1 gpc367 (
      {stage4_13[2]},
      {stage5_13[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor_CLA64_16 compressor_CLA64_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43b9102242ea3457c2af7664dcb9ea089e847a327c4574cec8df0c563386e86c465764dea296a98ab23e37036669e12e5a8778d0d4afd909371f4119f37f55603e3aad8eb36c4ad35f643c63abee9c0eba3c8b88e91ce73e8aa40a5fc3f632ff2c6947b6ad52c1a34409f3b91e8bf5023f1b2d3d1f969cbe87c2c65885b2b83f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h174cc21130bd69e3bbf0c19b288b6a55e68422af5d4e09917edb13b68cf620e42920729ef4b07a3749f419b6d388b1339cb74c5c34e118817b9483d450fca95446098deeb254cb3edef102f618f5d18f2ee5dee0de375db8ce5dd030a92bd5a4611b3a66e1cdf817af3f4604e8c1d8d02c8c778ebbc1c2e24e24d8e04ab2bbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5732efa7f53290d0ecadaba9871b58b0f145567cdf747b70acdccf2b066d2a0a1e5026b6a6ee16df1532eac1374ff667ca9a290659281d32b4eb505b13dfe4c8637e1a81eb6739dcecf575ee5308c5559fa1141a0f14588c71ce019e96a110c4029b493e69404a772fefeec11e49d97f1936764af2cf0ebefbe87585b9a9abd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bd3a9c88639f856fe53a13c9c3aaa5db0711cf5ba12289a954746740977a62bb0da1e14f12c94b9e12981579965d3407142d886a609a61cbd5238b73a069df9d52c952692cc15db65af0a8ed2242c6d4e069010027c0bb25ce5e57623212d2a7a36b0136d214c70ec9aff851ddefbe3220aa8d9918194c728348d9eabe1e7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha63d822d1a0f94c7da32b68915635b763311c106da1054f7fdba7e8e0a95502a296d2a4c8ac72d68a588a7ad6f153a3915d3b9932478afdaa146c24e23810471490b2ff60146b17ee1b8a3b588b92ccab4e22d188ebf5c84e0eb5989d84c8554454ed8f25f919103f1d5ce6d71ac715b4b55437de7ef32a0f321cfa6357f92f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab3955127d62ba4dcda09035caeebcec9209aaf561e1b525dacb3b6d20bb413cf82149bd5994bcd133907344a279b27802cb40da5b106e0987988dfd6be8a2ad1930c5b90277d666de2512872c812b5f9c639b5addf7ee565c59317eb2e7511eb9e174526fb6cbc1e0da6d714762bc3d8167100b1f92c4d63325e34531af9f32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb2d28ac8ae26d1545990ddba20e79ef42445a3baa06e269401584687a73a732a34172c89a2189b2ce97188a936dcb5a39835b86249695c3c4003677a94b29890781a5fa0617c4be77244187a6b7d359fd78beeee69dfa2b3876b2b1f57062d6a9e13f5423331aadd9cc82f4322c2c77940c83d15ab7394e51716ff520999911;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2068773b976c59003cb4564d1c2b5c1bf0ee3f0816cb74bccab84d8ac3c263a80a22fd171bcab992c1091fbd109a1ce86b37b3403a8d5308947146b919789ca077f7f3de24c3f648f504b6f1f442b442e30408700664be146baa025e0c6e54853fed21f3e3a2f0efd3a532b67084e650cd353b4add6f289a4a4ea4e0754653c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdadf109b70378f0b2808d82e788417b7900f1f18bfc2f7c6db54973398d511d9635ece250d2c09db1ca5f1177bd379843db8529a64ed68bf43de880eeb22a021bc4d99ac5de23b0f299aa50a0483019d674520a0cb37bd2b639903786d914dfe8e9564225b4abd26e16e18a59a0f147146cf00ab1d34dcf3fa5c49bf1ae7cd46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had410524aba027ab9d669f3f1c890812f2a841f318d2b5b739247b46be3112231d5c0b2557701f8b4ef36db1bd0cd2fab5a13df6c285e8aa3577a52c945b62b03899eb5b31e5f4f21c35271aa10bb3f2767d59af65d97bf0755481b15623e448618adc38060ba4d6b17a636fc2ee4d4e0089cc9f83445133c8ad938b2ab6f18f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b1c6fff6649919bfd95ebc9364c09698f91088c93ef9a333730fafdb5e97ad023058d048a08ae98e30b906c95f69ca1e2b51cfed1f3f638ae6b8e94820b8b547a9e9ac265a1119fbd0a94922cd5d65c68a507aec4beab77a12c16e76890daef7750fc7ec4418ca38814ce0327c9e0fbc7253bc36ea540c7bebf697d26f0e6ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c78a591cb738425c969b3d37dcb46d38e65d5465a388a1abad5f31d5cef77bd8cd74f3bb7be85f2cdd0bf5a5702280504ca3e302c4f5e9afb86823ee30fa74eb7f88eda49a6efa481600eeda121dda4b292d8bfbe84b18276538f684d4f0f2cd4da172e77a7f2e22e01c83ec3c9ea0a504a55a84e68ac3eedbd57b2e55aca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec5dd493952394be300c93ca2b69ce020eac264eb391ef057ce82ced1b0822cc32713e520f3a613ace6dda983319fbafb6a0d734c9ab42548285791cacdcf170cd49d4992ebcb55284082ff92cd3ea0ff730580c82df5075a740bbb51cff4c16761bf9c90174cce1525d592e8194f227e20879269acb1cd770edb39611bcc496;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8645a0c28e0913cf044af948d2a1350d66e4ca83b5be12aaab9e32754990a56bdfae6dda17d52afd0aa2d74c35d753c1070e4c5d29337e81d2b1017e5558cb2ddc69dbb57134a2cb8bcffdd33e48cbacc5554022cd6b10356a563fb0f8a222b90a57b5a78560d04207d90a39794980db92b428c200d78bd9826de90d549e065;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41de715386549eadcaf96ac8b7fd4354046eb894bdf5c12eb98710e70e94fec6d145ae01c21448e11019433c8d40b63571d29ed900993ab18f5f184d9f601bf23bd7a2dc62a8fab7283af1441d5a06f0e29653c0f477948413513937e0cb8805be67648940dd8be343b05ea5af9866ca6a291ed4f518b1610cf6580487f71a72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5e631334a3f8378facbf786ada1272aa36cf430c92ea4383bf251010eccea50e58d35225ce799a6f37a33f83574df955ee653eab4b38883ac174cc8cfe4c3baeae97b62ca45bd82f70acd99d80d4e68e59b781aa02fa397fbf34e2873d9d7252c4b0164ed122552faffc9072af50ef2a8b2a4d0364c74a678a5413e89c15577;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69a27e6b468794c5c82371eeec610e4789cd800f47d56ff8b4308e5d78b337a5bb06163d81208eec9bd08dc5861ba105e0154bb38930e210188d4446e7dcc4f07d37f091856428723f3f043214a2699570c91fc0dadd4d6ccd74c5d93f170703094173f557e8a3d362e79dd6711deaca35a1d3c61b8c71e94952af0a0aa513d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha664c48ae5973cd702805e7f57fcc309c605b1bfe2e9e7daf870f782c4ff84514273ede5a910b5d1aa4c3f7b3075480da7cfb231d0d3189402f515e940b550c4b817d2a3033b07033247fe1eab02f0e385e5103f27c4ec189e56c380fd0f1e02ef9872fe2d072e0c8c7f13656ebaca8be97dc8cfe6e2913dc965f12a7420377d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b995f8c9504dc8b3d6dc063612de3b147969af1af7cb041fff1a0c1850f9639cd0fc015f4f809ac159949d07a95881c5325006c3508861466c1db7c2a42e17a76251668949ed4946ba763a792ff52cb541deb96067468f2b3ecef2cdcdf259b41c43e51f37d19f30dcc2695459166e64a1802e6bfe75124acae6a103e6520a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5228fc7e6ebcb545a316e2e80c9ce73840a3b694b656045c0da58b35f50bdca5df6af80dc67f530d1cbfb3bf5c9e0563db697c45e262e16631e51a8db163c8146215d5922d9cbfc5d03fec0d8574092ce5fdac13a0d872f0422eb5264b428394e8c06220d528a296e2a3ed35abb0fbd42bbaedea34b40d844e69675bdd8f345a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0ba5d40e27ab059cef225279a6193efe49db8e1255a41562f7630f7dfc5c6a7f950d3314f8e826e82ac5bfb1aad0c891f3aa378d749d1d21a7f8a2708841571e5c50b9c423ee1fa3dac66be99e8ea53e8ab27ab5d0ccff5ae1ddc10cacbb7c984312f56f279078acacf101f822a9e789629c4cb02e8c2f808172688daa7bed3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80853fb0ad4b17335c00292e3487dbf566d7a55f8b972e0cc62dea487f858bcedc417cc70e31019a5c0fb1b1fa4403ca153efd8f7265f5881c945940208728cf09100ab80386775cbe0ec89ec4634274cd0d7706fc0f0be7d1549f1a2ea9d9e669682f001ee2700d2030e2d2da771437a98fd51ee514c72e8f96585da1a61405;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h391fa3d6577da5c732b758d09ad16454baf5de861d6ebcac211762aca6552b2864c852f563f271552bef8bad4daf8b144d3c9c5bbceb62b1c4c6aadba26aab0b7a90a1069333544bad0ec515499fde0fbd651a6872435776a9fb8c1c28b44db2d3f0c4ee1242a812a1df886c69748a68923c79c83e78e85bf1aeada59b0bde71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h398ad4f33d060d4dfe49f27611c58ad21753cc619a76bdc6a2d18f94dce53ddbcf61af1907595f76e94ebfbaece5cc1e89d41638840840f439fc9a32243430dd9acd1f5ab2fd857d8cb183905f761618dd0b2eb294d0554623d4994cb7bc88952b635bab88b16a16c2df0111a6535934bd9cc0b5c29f6610b71d180fdb6a32f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f650c8f7a3f1c01e4a590c43d4bfc4efcc9026dd4220e02816425659131097e688aac1925dc4386a0706613a53a48a7081cff214e0bf857b436c0a2d2ba7b83a8ee981be9e2361d78abf5d1200fc6d32263c63f4991401e101a6baa484f278f0878f1ad651b08a132f72372218c0218cac5c81c69ccd98ad529cdad6f07f31a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cd3dfadad118798c3981bdda3671db8e153c0c48a24f9503c020584d4d2af8094f8c45f04f4348611ef933013c3185346a4d48922475aaf74d391125eb537b30f865a48afa2ef4a7bcdd2249e62526f689454e71a905763d6c3074edf9b6a1312cc4184f358c57a73bb03da10e93af598bf1abfb9a3458a3a566b14f71d9bd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4d6d078c9cc774f0f11bffe0c21789e6bb48858d791b9a0291d951ceb0610dcbf36b25f6a6650bb46351fb15cd715cb3e5096bf626fe9fdba708a6c6f5bfbe461a0e4abd671f63eae9cc8e382b53d14b217ceb39c911162bd555969164bb0d5cb084a35364cbaa9106399bad0cae6e429c27b3317437cc4805353b28314e4ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87d53ca22be4132810b2dbd3ae196841c3a598e88570ec270952488a8e5fcb04403701258f003826082039f75e7462924f42192bfeca01761d7919832ee839b38953b08b48836ec554064f67a2e596f21c074f893e4529f0875ec173bcc8aa23c6030d5414fd4a5a9cccf1ad7a34f48960dd4f43937600b7c724e3aff6ae48fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cd9b2c2e06cdec0fd482f6d3597136b2b5d3bed88e297fe622dda73eda0dde7730c98f93c01da1eac2d48c97a80c5832ce63ef32e245fee91753a8938ea6ad8d235130a42e230e59e09a0e3333f58da7dc0c6706f3b6ce852efbc51e0e38177e0790d966b5d08719a6ebbf794d6407ef209c9e2df73453bd51398f9a9ff856d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1079050e8d2d2842ffa3933f8d69d94a25f240f63933628cb32c17eb0e8f9ce2f74511caee850f44b6adce86eb3af31783c97641898397d83928c724dd1825e573ec67f75f21a3c10376370e0e3924619632df6b4d282810674286899f483bc097be3949d6946ab08947fbcfe94a6b72d55fbb208cfe4fe0ae1821ba2faa49d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf49354bb2b0237c50dffc77f0d62db9ea6e7894fc6642b0eb876f2f6f748dbf330a5d47830304918321a02964139290ef9f7d220115de6811ac5fc96486520e2100e7889deda125ef6ac25eb7f865364add8a557a602fb8acaa0b504447fc50c227a7fa50247eb71d3685d26e76eb34bbeeb836f816d6bc42bbf3adbb8a992d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbfcdbecb9a4da41505ad3bfe94aceaaba6cced69ef5ccad0c8bc0a799d1ca4db2198ee3a2268132e7125c060b9fe9e8e3d7441990b682c5940d7e496d8d2302a7899c4b00e3928790df1b18f88b885c630deb70e5a69cd1c075085c34d18dba3674f3c98db1b061a46714a38c2d47455a6ebe091cfff0bebde2635f5a523666;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dd65ada39d25ed4474d3d35f01784cdb1d136532223eb43ac7e9d6503d8b303696a64d1b48ca7a25eb4d992275e300bc3832b2328caacb3b1483209e3569839c32947d2927b71a2e9857baaf29e80ff085b540291fc5e0a3fd00e483fddc69050a31ef76f4cb1380cba3f62f252c310ace0a3ec659efc0e7f0b3309aeed93d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d4f44fc1319642947035b013c503e4534ed29b7204f8b5d602b2472d03e147fd4057ea62f485032f57defd865b97aa2c6944c544a98e4d68088c6a8f99a8d74bfb43b752800c1d8dbf01d07feba76c2634a82762de8bc90dd49253bb47ae263f271528356c304198b66c747e84e9ef9c4814fe0449811fcbbac2d47664b857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ed6d64775df9e136ccacaf23325b050d048af3022ee3d68347c25be34fb44760c51b837b743b2ef6d9bdf0f39605fca54e6b8247c5c7d65cc4bda8194d2d846d03b7b297db25e5a00157fbeb3463e30e160d77563f5519de52f1214d46cc4064212d355043348b1cb978f13923074233ee2acc6010225c37321450f00b9b782;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he89a2552eab24671d49020322560ec7652f94450aa54dcc5d460a84f814a144bf813559aa2a9bdbaa825fb8558b0e256a3c123fe41c3ead38fc0d7e4040a5f2e3a8279125145e5df0899e8eaa237412b4d9ef0c167f5a3bcb7632eb48476420ec7f44942c847db6ed3545c9d62ff85158a40a9e4c2e4b466fbc1a571d224e30c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3a82c0907c3fd680bd835a3f961d2f6ca14f3da81c509b5d37fe8f955ea6a1d2cfd5fabe850604da74c2854763596ce935b27dfed01536e87e1f993c282ca19279dfb0e55a8d00d8f9d37aaaeb08d3b752bf4c3e5c7957e2e75dd893d3857611d211d89b5c28ae901178201818ef59f0b6742e67957831c84bb5607c957f77a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61a54798b151acdd84211e653ca4d0c3e7146b8cc1beda18b434063f5f68775997067bfc7a57ff35138609f6fdc4bccac22f6449c36597c9423681e545c09453d246de4e4093c2dfe86c4a3824908018ce34ff7d0f03dfadc9fa53173e7da412c8a598a699f5d6abd1f0569704016304cecfcd9eb29944199fce68a7c0f29353;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40dd404e1bb011fc2ca82f8f065cefd647f6ca253ce5f19fc861c5c22ab0fd9abeae1da3224d239372d35ed576fa073039dba6585807ffcc27b749b34328fdb1032656ab84e04574689b166005fdb30abc0877ad0ded69bd05f8c23bc77cb3e5e9951f8b2ae432b7d7fafd8a111fa2780991b3efed860dc0809d24b1e13a6f4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3877b7be248fca684f545c65e09cb3c144a76b216f2a2a4a873bd5d110b2e37b8335babb804e3ea335f92dea4f7a281137bbf8509c3e173fa672f9ddf1426893206dcf634898b6ee32518a249847d19200489d368b56468d99be376d43c35812bcb2ec812eb9b0dd77150f266871932f9b161fd032e4e5d7fd0b9502b8933cee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd510d513cf3b86fc50894276e27febc5bf4924fe1748de69f34339795c181252571a41489b4611d51d48fbec6986a23b8fcf4e7fde64669bdba2321081c1fc65d5a01e7b3ed354ac777922f38fc7d5c00755871c238a0cb008121a0d4139ff8cfe6d12fb2a55a8f09bfaab82d0fc0bad0939a33f525b9957a350c40bbae4c1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c9e5e615ce9f509bb92fcbe7d93628c1c9fc2a18ac0dfaa645dd659e7b171ab05e1058e17acc8d10bfab9ae04e1f1db0b1a4893f27e31ecda3ef84a89eff9f2745804c0df87ea88def1878aafd75fc4077a7f007d3032bef74e1770b63f2bb4503d7e25d41565031c686f455d6061c87f8a71ccb95bce368bdffcc407bd466f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf9ca840dea64773d1460a62871c7ba76b7a0c75f0835328941c2e586c7f1e6a2e8f2d769506fa837795e3fc917938d774b38478cfe350682a0e3713acef62a6395f643dad2a266f7dbf6a4e7dac2961fc0f54f604489e0858cc1ce274e24bb31071f6b4371ca664d04dfa3f5728bef7e6a0d2500a687eb6683ae50c2adbc4cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e51d07bece7848e75afbe039a4c942a8e44362250d7ec77d377fc0cf5c128060c656fcde527b0762a799353b1e6d9ef73e733396c34c180973cb9e62ac967c05fc73bf74638ca9d7a3f77b22e71dad9920e14ac34b6f085cbeebbf10c01250cc480fc33bfb7c26233364570cdc2e761c55e48d46e9d69fb32983cb67f373b50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a33eb59c2faad483e9a34e4347e5dc3a76945a034413eff24d7b88d671777ea9f6c0bad04ac09b464bc4b10d7ed29ccb51f4e8a443d7a418c92a4844281469f1b4505ff8260550e37f8e7a3f72c415cd89ffa0d767e5c32d42592f6a82956fc516e0a973f63f624cf346aad051981622472854d0541d20d0f11f841e4848da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9e1241e9c324d629753674edebebc7d541bdc1e90a8c649e2d89056d602a40c6fb3aff0ba0972bdd8196bbc7cc786852da6301ae17f652cf5cfccfc0a664eddaba668d4560c9eb9a25308f53eddbd482ed0edee09b0edd2864b6181eba1d1bc3f550a480f56fb14899b651b3f2d41cadc1c18cb66f9040d6429ab3aa155954e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9defb1fdd57600538c5522f21b47e5b17e46fdf37a3f1e3c766fdcca10630c41340193c8d9eeca3ba7c83bcd55eea5bcc0e3d1088e22f4d1db12eb8ac27117fc02ca7e61cb72b97c7e7c9b6d29ce31019aedeb71b51255d664455c7f10fe82f035a50c59ec6055fd8b4a2bac05ae5d45b1cc3f9a44ce8eb4d57e0db8b5d0d135;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2debb450a3aba593af01360457c806259cc9276611df8acadb4b47ea4442a52e1d6780051a02d3e93dc4ea0c374636e87c61e982a27e79d57b19bc506e5561a11118591576d08bb51b449102c2e68a7b306de4613fc19b92bff09ebb825ccbce4d96b58a1f17a0f6066306b69d15248728fcc9088847d58478fdf4373b1ad6e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f5d52b24751d14eb6d5b8d9b99cdc39818adc47f9d7bcaf3010e15adf2bc859db8e6c02590235d5990986caa5d8f8aeecad5ea656fb2d128c13626d9a1e4225b5640aa1f607abeb69cc37b5d560946e206a851c1004f162963ffd05f267a1dba31185cb82e8d22e01d26948a655a38d6a3b830bf804df5b01d185c082844e14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd16ce78be7beff185568f7be3e31f777f58d3f99bca255aec6282b7fa4d4587cdaac186c8691228da71b67faff4e019127d68e3976ca34729021af4714ff4c76c4ed0d9c3925a9ff56147d64958b087f9a816bc27284616e7b6dd8c3fe0de08bfc0d0217db101ffc8c9876aa5fbb09f5cd890c6ce6514af66b086a86394379e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf08d6dc2403983c1c4a1af9c052148170de936fd7f1c0cf61b48b98b5083763dcd56fa5f057c71b9e92926f6c2056f429f02522cac6306f978093e2464712c1499ed96b487e1715837d764c41295647aec674c3e0d108126844dedb15310945e591ea75e7ac65d5f87822b6fc63a20b561df05b1296b66635f061e1f59f933ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3ec91d8151ce3798a1bf83bf45c6a843e3c25c4df311cb73a68b60487b38fb85fefa5a7b79657da60a8343b0ff3bedb970a96bd08986792e8e4591361d71a32f0ca09c5b94a327cb1f5626720a3b73e573efceb63f0964810a1818243f1f318e58cc90f94f65b1782c535d6c3474bce73cfe90c759407aa445875378abd086d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69765e29dc70ad10e6d0b5b1e351295c8347420d688ae638eee06f79e4b0c6d5ab1a8384e478ae490f72b2db23643a5e8ed19d837abc3c82b670a8d95bc2a485b459f0c84ef2ef8e1c1d455a9b10db5085ee67968ea72878b29245328cd163a7d37cfe19cb8c18ed436794c6dc47977d9345f9be549795bc780e7556a4d30180;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b3ea093be896716ef8b66847f50b31cdbf6d32b9c8d26f71ade11b73e94c6afd730931b958ddaf368655568eab15ac323d497dc5610cc3d9416a41f633b5846b8dc6972e7fdad5130ad4a591243dba1aacd0dff579b4c0ff14f8cbc2b84f3dcd52ea6f27ac18a06d258fc315c19059a8838915eb2510d3485399716a07f776c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8562abfbd2c17a2e5437779842708f4fa84ff4cb3b788d1301b0c215bbdfb119d68496aefc408f48be882d51bd4b0c5c51a94a35cdba8cb440cb6b1f8e586c63b56f492bddbeb6b508e6991ef8aa89438458b09e93c1f52ec54cf7e6dc321ef9c750c3af793a53b1dc9f857f0d07ee613e9cd87335fcf4e9f5e0443fcedba2f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8999e62c326020f2ff53f94fd8d757b114c290077f84ea13b6fb633af6bc9d9be2cc9ffc7c8ab1f07baad6c011881b227b7866e4d8385a76b378adc2a29152cad60c93610c5a8ebc6055d0855e0ef2b9be020f71addf5ca449b1a9420972fa96f5f1e2a7c40a6ba5390503a55264e627e35f1a860f9f4b0260022258dc35fbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf301e78174ac68dd45e753b49cbfc1fffa7b8d8e9cc7905788f0eddc159b645d5e39fcf350420d45519e321548cbecfacf2b60337f9e07e4c3f1552ec86703e4918e7174f6566ec352da7138773b0c9652dc3b9a347a83ed22f53024ce0c4107b07eca0f0691129b1f7117b4de09255efa3c72f18d83921ac0374b5852bc0813;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b1472e56f5c94d2b1ff0b514f7f9e5ab78610b8a6d38d4c71e93edd1da055a9a64aa5295734f826acf63384db5b49fcfb7c097b5a560b9dc3f45b67334fa025d4e922da3d749e29e75d682bcb1445d2a7aeaf4328de986586814d4e35ec4bdc82657251e3be5e1efa7a0d3d7e16ba0aef54a841db9b7b939a7d9f3a1adcc48e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ee45b067150dca767ec5cc8f0e19721586d96bf63c5dda55efe617ef58531bd414eb6f3da0491d05c3d68b66aec6809a722679ba3991574690dff90d51d6e7c1da3f7cb1eb687de8f61553470c94fe8e619b61a1401c72187f8dcd8ab0d08c0975c3c0364d47be1d7039212dc4be246b3f758aba975af81ccc749569e92139a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3881378dddeba3b89a6a9882f830ac333cad9978d74ff6d0a93bbf6b99ef433a2080b11736ff0683a636e4433379a8ea2eba567d1f7dd45f51b635973b1fbc27ddfc27499586d57660fd4047cc1bfb8a0a155b43d5f3d6918fc1332b2f936739c377590aefb4ad5e302f31ae9f6710be4f0fc0a133a4abd6893cf623f80b87f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc11f10c69973cf2eb0f53190d98151114d349864729125137ec3865a6f71b02f82efe758fbcccbf2b3a30430690c63575335f6c9ae6849c1b25af02491b31b208fca277c6ccac4dbeb5d56360c50a1e49d22dae3982b10705a56577ed07c75235a83815848c30c471bad5a0835ee644a0b03a0ea1f26bc5a3b2bbee4f866e178;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a66fd26c5843ef43ba45f7551b64697260dfddcae0f4d254001aeb88116ccc18122ce0b8638ef054b1e978909f02439f61d1faa133d1bfeb9b40ad0bbd382e1267b2a97c6041ef99b07d351f9cdef914757c1c85a6b0ae6eb0948ad1140bb6afebbcae5550f9801b7ff79ae29131c1c1d77a2b2928f5d347b86a7946ba78b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86ed093243b84355e58cdc0189e88be350f57f73d44f8dbcec66c04dbbb031050b041d749072debfeb8e9becc11b18fb9d61b89bccc9e0762ee688d2ab60d1634a0b5dba1ba82781af68a928672cfcfa541e469b8ce491a86cf958709063576250ea681b499802ef53bab9736b37aee0789458acb51a0464b16561b5a9e4f295;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86e2cd925e6c0609eac23785b0f9aecbac5de7ec286a798128e39b2371a93a28d510299cea521b54dd573377caf8e1d38954fae71900537acd29993f97d86e03e274fde7e1b5605e1802741c5999836e1bba4ca247fe932d75650a6506f36350519e1d72a39280982eb373534403a06a699b007049e62465d09a0bd2fadffb4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h298a615fea1876c026970932cf86b71d1ea8600fa49be989c80b12a918e230b406fcf7fea16c018f3c7701f6276f8eb359a5882d7f81ee6886030c4eb54ad4536b4a0cbf3454e7b0c92b35e4510c40a37cb5e9149d7470a11f80b189eee556858cd00e90ec3223248af4a27cedf0bd3e244a06508a5f0fa17efd4ebdc4983b35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88c3a34a5971dbc506eca52ccc07a8ecbdf25b40d87bf55abfc425e3f446b407c993aa121b6d00374a500f84514c122c9d2c7b72e36caa822716d9b2a8828b5a5c29d0360b7efa32a5c70914870ce9993a4865d5bd1a3e75eeea92d8696124692d217a4aa55657d700edabb38ab2d28227b325c68741191598c4d6b81dc15bce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd88d275d10cc60f96a8e31ab1842207e34e75e5b9df4fd6daa6a0ca35581ea1209fa01fc9b052959b26fb5c0d5f5b257f777cee2b9ee400ff194d8e3b17affb3fc5231c3fcc8a9aac109c04d01a17d908c7752f963bebf56ac645e0cbb8d079c46e80daff7f4748efc9be2a14ba20ac0794e30ab05e30aeffcbe4dc8c19c320;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h103fa910a1f1ad7a1185ffd3674044ca52566bc524adac780058f77b8054257f740f69669a59bc93b0ba12f8954cba5a943161d29584d1bfccb6b9b8d091faf3c6e795d31d33241c21234b02edd2e7e6393105824dc37a230d1f3b53ca95771bccdc68f1ace53e00bf0349bfc77129a008769fbeb9bd23a7034d33303dc04340;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h754bef99b047d4b9c551bfac84492c350047b578e214f90c6551995938acb593adfb08f1d55ada83ed830a8df0262af4563f82c43b5b58d6848d8f950b633048d3485eadb7dcd272797a5b5c1769ee960f9ed6dd77c195f9f9e4efcc333d35523efcf7bcdd17de6df4ade66900dbbe47fffee19fd71a14597f95f705e191e56e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bacfb0df3af968d759d95c783ab9788a5a17a1a9330aa8f21dc43e9c182eba3eaae732c419f3d7c3cca7cb5b18675801d7aee62ae5bc479a46e9fdf9138f33626554d5f69db7fd8d31c062691d6332ace1754d5612107b5344b0d0f162030e30fb437a6ea865726106b69c2baccf15f2f44188c05f2d8e4c2d408939c88a02a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47018bdc4825940c6ad5c23bcac646ba39e5010a216eea42f0633e73b1cd29045600b397fa97a34222e9d47b7549023004fb577b1c0dddbf0882061e0d8727195fdbbd96c7a92a54ad220539723f69c822383e04bebdb76f5789b2003bc910f8626aeccb72ea1688f04ea4d8b7e3b0ce8e84b3d051f9933ac7f9cd5943c1b29d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2553c624f7484e308742c88948e00cdbca877c81dee275d0ffe8ab1f2db60794f237c3005e91083fa402eadac1fd2c1044c3b89edb84170ea10232797aa263a3b0a52ff8f546fd7f26d222bb652bfbc6f7bfbb35faf6e20a94f573ae86a57d6b84b593e5fa1fa6348cfb7b38d39a4009e0ce52068b80fe7131d4bfa63643dbfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2cd233f79a50ea48cfb82ccca1fd871197fff06b558dc0f57db94b3536cf83a6e950c1b07e907571b43d79613e7f7f04830072ddfa87842424680eaa9635c967f07d3087ba4c69bc635039f6717fa82036840bbbd1d8c810ace386ad3ea2deeafcf35a345c72b5b4d4d452f511f2e1293fd8ceba72c493bb97f26c295e4940f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ead11f56911bb31ca2ffceded58d5b3af78c930063fb6797a207d2f18d9ef32d52c41929d3dfea7963908c7ed03cd46f160759d5b9bf359aec991032f1161745b5e6276e254c4e484138df3e471cd3c89a306f3d1279d4a8c3677b64d502ff72ca1385147994f6ec80e1c6a77062426ba3f8ecded616dba300a716cdac4ce4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedbdad1ea3aa91b0a115e2d0fffe11cf230da847e0e7258558c148b3755361589c0e2cfddad6d4c301f26f479adb9ab9a5f874c0d0372ed0d436986c8b359f74bd3825902200b5c7630338f9a88db9ca447c876f498aaa1842717cb0cde049086a807929a421e4bdca677946f9c9c5047ce553dc05737e9b6d7fbbbee9292809;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0b9f794ed044c90a9aa52ab22be84940ad8566753bf341ee035027a61ccf69b086eeba025c756d47d2e1472df464c5435273685d848d8cbdabbd98bda294fb1f56f0ea292701e446741044ec2001e275307da591eebed73f6e35646e131274d99c76f99840f9be6206ae999b791a2803c085ab182f78cb4e553e6ca0b4cc574;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcadc9d1b2ba71faadedb26e82206da3646f1b7e6edb9ff064d91f73385aadf0362511e5d63d37a9528a4412487b44a14d81ed50d0cd6af4cb398e5a169bea03e1492d3c06b599282c342b314c4ff6a92365a47e2f44f7c5e5df3c672565c2a267b96a3f964c63873ab845b3418220adfb5c9dd1232755a1123c3e05eb4bb32d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ab138a94a9dd93f79365521fdc9bd20b1b74ae6bce193d25efed5dd21635e8a5e1b8f34dd5ad446d3eac7af63f59bee350c0446d22e35634028fadebaf0154ec070cd8aa855101640e269de669e84ca1d077aad661a0f4d3dc4ae74a9cabe3b05c21cf4013e2edfe732d78ab6eccc1ff7948f2fc5aa85494b8ea263e8f9ca65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h251b53abbd0ae4a494b2c893c088b6d6829ab5d8f3fcf106b8b954029a4ceadfc904062a01cff671e027b07e22ed8d9bea59543747b67beb815f2b4d35393837a2706430a5dc97d601f9caec049d2c94aca9fdb06a22047e6f5e8dfe77873f2aa69822f66c423777643412930a9ef9d8164bbdfd5267f618634155d33c234c15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0152b869e0b035c8c9e4793f80001f045517da137022c5b8f26ca513540eb66c7650ea05a0a45538338184f613179d81f7fb85f874f477db2840d73da45b799cacd4bd928587e6910f07e5a03a95e33fa6b129f7e65e0e9ca08de391fb0b6cbf3e40606215bf7bf007c27a29e8922b5fd55ff976469452394b19f198e263dd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81b1d6eaaf79245b0f88ca6a607a517f2de07049894c547fb401d176f2a2967939c540a417e084fe459610006ed99d3462d109ba9700205b011dda8aabc728a8169450d3f6fe1aab1e78af64c9e26f9bebb4171f59c57ae0e09a7133e3daab5634190fbc77ac39b8513665e7d51e2be0f732899e41b57bf913567d774a0b16f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8b75f5d3308f3bff899e98d49007dd3a27de60d0a250446a3a0847cbb144d2f50d610350486cd057db5389a9fef33cb49a659ebaa516cc4692df42aa0ab7578fd7ea9e7a358be2c93296e4f2b11794b7a29a8f7a4d6a4d08496f7b8851f6d61d2527b5f23d74b952d8916364712edeb53666469d1f783c442f9e1b56998641c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb03e42b1086a9796dd48437d67f76c6ce16019ea13a7fd53a49c78d01d7923b6f55175aa1e51109870345a14c572686cf6957aa34803f8235590a3f18e3868948773084a0c6c28d2fa2d31a95a4ed04e082e4b8eda236d94d27a27ed29efc516bfee818f20d962b261234be57e5e8f882f9c409ce8cbbb089eb8f03c431ab5ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e79293c5c706d87700275c1221a4ccfe3c961779985ae05264a730674a33412ee83ff0678c4575099f3f29bf740926206f09a580cc834894a89545b6568dc61f3511796c919ef85eb8e41137cfc09f4578d89db6d251f7ad205de61fe5b77213a4a9d5d38e1f64edf3f9fe1430a49b05967988997771a021b4edbcdf524cff1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9082fdbb573aab71b311218ccfa41211e114689b2ffbe9f0ec3759b276828e81baaf284eea9f4c9937ef25ad1d9f9e766795fabb2a9d5bdbd907ee4c27a4e8d41621d059cadc8b620c4b88a6acbd5161d57f98100f065544777caa903912361793b50171a436af111297fdf73ac9b8a030678e3c7e0d4be106c569163a7ba82e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h644759ec2a17246310cc8ff4f5e8587dd448440f31fcf6d6a155ce9bc13f415027908ace9fd50bc3b0d71b66185bd9c1c663546e9434132d8d134d722c5306d4d28adaa060c481ab0c0fd6fdaa8f7b6e7a5e9e53b6dfdb6c32f958d29756f6f2475925f6d409f51d98bc7c9628775cc6d65ffeae4b6cb0397cc291b83e4aa196;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f462b879f5f340b7fa712ca4697c9258e74cc076ab3c18cfb6782ab9500fba97b771cb8fabb48808654268032a11ec0750a5484475058bbc8177d934a85f5de553d8d08c63d75f7f438b88bc2cfc92ab715bb803ba00771c32c4ede7c278965c7ed3f018c8b5fedf2261a93c0e90dd49b7ff3fceedc6940854d5f31f2ad1b1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80b43e7d7dedd6b2d6ff36bd666600ade5ddd113d0736ace6aff4855675647897f3246db80d3e4ecbf7c11d137e3a364ad81382677efeaa477ccd8d5844dd847b28d7a37b9909e05f415c20e69622727a2b26bfd470a3341f4f8693e8484c24b41c3f4368dc5ea162facd0bcb2d370fbeab94f20df0ef8b6251b493a07139020;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13a2afc9b5003c7fbf6d469239a0c2e4fba49051704c05889095e1cb36452ec1c7f671d89e80306b6f72d374fecf6b9f964bcae31f8b50bc747c7a7914aa8002cc633db6b75f7f80bc25206d0c897c7377053990e10c55d11be4548ef7ae19a589b4ef7ca0b197bde07f3cf0fc1ebdbc4067d8ebf8f8ee689cdb4ab62c69c31a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd53b9007c8aaca47573ca990f9d9fd74d1c4710ccf7877d9e54b7d1cb0b90eb91eae926c714179a1ca1c24804dce1e73b79dcfc0bff560beeaf66049ae12b611262889d1736f16f8a04c3d661e128741fe6b01d39b946354960e6bee7746f55cd2c4985cb08d1f81e0fa7b84d59ef54df6723a84da5a33b112c714e563be9455;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8199524eb71422556e04de310bd8af4e7a336095da6d89f4bd696bc592b9527471a2636086c94691f1039df699313a7066fd3b611da3ec5a0723f9be3c6a62187703876bdec4e2fea2855d83999b9542811fa6cc2983c75ffe3adea2e92e5b42c55aa1e65330971b354cdc81877b931e776ff9236ab19d811249d0d407bc7d9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f9e3fd07b92675db44e05bd9b35ca6de481e5ce72f40d9fa0b3861a73f6623d719be57cf7c0747731a8c352907566c8b803fb2c90dce842cde3fa56524d55aab13b20c9a6fb02b068ab9accdb99fef92b1ef5dc9ac515344400e5cef8363f93f1ab9918834036fb05fa116514ece98d523e6d50486f422d317224a5fb8354d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he610afa5b29cb6db4b3798bf74c6c85e6418c185d131beac4c7eefd6b00a156a9f7ca9b5bc7064c1be2c929f7dd433da4a17b7e2c2634d2bd8f7ef6ba3d9b58d2e89c874a046906a6ce12b9b0259416f97d2758af6f97c235069175fc70348472ea85dbbf21dbde06c8f7b0526efc811f98f318c05d30bc88004c528c2ae3d7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61dc411bb5bff5132c4cf0becdef5861744015e9c41c51fb7123d1156be275abd19bb7bb266e216d5c412a0acd2df1c23621d79c26deb8cabf5c6f6b6c4e3b52392f9a1cc04198f41018b6c89986f76e45c4b81dc8cc2e613d6e1a6a64fb78b3e89fc38241b1642a111093dc3479804089bac5af815b6697e8424601f093642;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf22ec2bd8a80787fb3ff4d35b74db63b51cc07a72410c0258788b2d330039fe71da51e56e8735b8432cf51f2971f1921eb3b579ec6a7ae9bfd30fa7db1be1f3de9b47001c31b8a992faa4f39f28089c30884999b8eb3114a82b6f5d3800765f321d3021e3126215c02feaf01fedc81e652cef5d40c0145d7a1182b9fa3696dc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h255c206d330281be1590bd04fdcf3b0836b59eccda68aff057c1b9f803a7ab18fa8d31459d5460b7714f8f572a7b189bcb9eb6cb9e5bdb0dfbb4c0a2c0ee1c6f3b6f4fc3fb56d8978842825f5cbf66bc44fb88581c3a8d57d23bbea22e52f56d12def6a000309f2de6624fd7dd8400500ee0481bb8f82bfcc133219a336148e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cedca025cef28bd4ce5b16a2850235b56c848b0d4a1acbb13f957a5b5bf05e301a5c502100df764fa06fb712881a607abcf89f4d92c0b7c23108a9ba5279d66a77f6bc32bc5b250c05ad2357e9460385e5b901b9950741fdbcfc95e476ae2c214e5a12c14fdeb35d5ce8a61767339063ac370fe6df83f7d5f011cd805ec1aa5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b8fca70ee54f5b30caf8eeebbc5f4951f52da119f088008d89e9bfc18a148138269f96b5d225b4036eed125b767803e80a2970b81283176be968a23b691c65ae20b56e0f3df1d1048fbd4c5914728f844d1170144d020cd1629e4bc0d81b971985aab6b40da831c99d3bd72216c35e6da22106b62717fde4474795ab260bd14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h685fee71b809904830c8b67514c144e0dde1305efce42ec9b43fddea0f00f002299b4773b0d0d41b2168572e6f466fdcf3494c3480875f64d6e50d2fae7ee277a95c42251904a2b96835cfbf4a8f4b92ea3c3ee104e738b1fe99423528292546e00b0917c6dac0da01ff3be942614b9cc7f4b99e345feb06a7e9959b223d4fd7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6c435cd5c0a1318fb139ad8c67da72af89ef70fdfdfc1791ec68794999f769d023af0e6ed5f2ffbcacbec98dbaa99fa38f55fa32894d524e31b0b6b8d91325bea1d9cc6e58ae9fa5fc696bca9fddbe419aaf9956cf132e8c4fc2b2646dde0a3077a4bbcc39f4806056fdf2b5d80c5886f2eb1d68dc8ed32611a11bcae3241c;
        #1
        $finish();
    end
endmodule
