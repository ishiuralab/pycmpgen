module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [22:0] src24;
    reg [21:0] src25;
    reg [20:0] src26;
    reg [19:0] src27;
    reg [18:0] src28;
    reg [17:0] src29;
    reg [16:0] src30;
    reg [15:0] src31;
    reg [14:0] src32;
    reg [13:0] src33;
    reg [12:0] src34;
    reg [11:0] src35;
    reg [10:0] src36;
    reg [9:0] src37;
    reg [8:0] src38;
    reg [7:0] src39;
    reg [6:0] src40;
    reg [5:0] src41;
    reg [4:0] src42;
    reg [3:0] src43;
    reg [2:0] src44;
    reg [1:0] src45;
    reg [0:0] src46;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [47:0] srcsum;
    wire [47:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3])<<43) + ((src44[0] + src44[1] + src44[2])<<44) + ((src45[0] + src45[1])<<45) + ((src46[0])<<46);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h406de03406084417b4e94479a181532abff724915b158200b7930dccd967e5e0a804c607ede5f39d5dceb709335baa5bdd54100584a89c2d7e62696690674d26efe16e14399eef4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27fdc8860415506c68e26b29a5402ddf93f6c2b0106009d3e254adf6383b32dab2a3a543ab6585b63cc969f58d5a00228bddfe53846b86b2da40608dda49d42d3740f031561a1f7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9724397823b989e5ea6f8d40616f2d8b57017a4a897a74b29c6090411845fa1861ae6f51823d0009939037e06d33b7f3ba74029f55cd4b290db51e2b8a52cff81499ce5473611270;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c0b9ba7f59ab813c07cc35ec03a134ab5052ea4e0db935a55e563a3c0f462cc95af89a7f07ab2c0a25798a594f1ababccc0c30c13802212f60ce40d53a6f944663f2e1c4d3c64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcbb778b2ec12dd4c5e52f12faabba7b8dea1f7e67ea1170830b3e663bf24656013c3a3f31ab34e9c02cec335cff0a0c14b6914ffc0b507e42a5915dad7c78cab463414c77d79b64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6b40edb3b134b7b659c2aac55784ebdc20c5eb27755afd98972b90bd4e9ed1d6e39529055040c53fdd1008716a4e519a2740b8337c19196fee2743a0bef03a09a4508c610fbf058;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4450b282f71ff97cab7ad0996273b4d1d5da17b52a250165b1cca14880365e9f0fb23268161131cb3d25fb59be0abaf0705c4c93b2e7a3c89267a6ad504269fb880f620540dd45d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7677c71430541d5ce1ea3eca9b42d0b31701d1f5ba2f90ec3dd86ffdd46b24096aeeb26507932aedad7521459a056c6ffba12c4f46660add19f0517a5f560678d5c0f600aca9f64e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ad70ea006dd5d05b6188a450f66c49558331b50e372f54a24418eaa7199b543d31c795cde0a5570d7b211820caff10d255e7d7500574a7230137195711a384cc9554477afccd560;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h302ce5a56292affcd1c728e06d26a8c55f8dea9f1b2803b92cef6743c6944d6aee3ec20e0a8db306e539fae1417517a0803e55655d9b49798a94a36da1ebca2c2edebb0b86cae7c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h381976ef07ea333a92c7aa67a6579e588cc2528785b1d3a2ad62b7aa1e1d0e20da4dd6f03facf684c73bed80f84da4584e6b1d519fe233f1249517c8898d877ff3533e3bad125fae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a3ca360f4a568eb065825dfc1822026f4e66c984bd3d56da02d6cf6eea684c30d7f893aa11027c4bcb25286ac65bfb46474bdc02f6caff8b6d1d73f129406e1fb5ddd46b3441a75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7c7c6915f66f3f58a68c1b606de2f03d645361eb88e75d14067beeef51ff81bda380509a8d62a5078fffb64b41b3512dcd86d3b2c6ccf3830cc0f9467666fbd846722da69c9e307;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h889b3e07d9c4983390b1120cd13f18fbbe0dc979afeac0042567805dcc75c4d1eaa41323a72bd195caea2469c8176fdda914662ccf7e9708aa3cab6a7c739dd0c0cbb2ef6bbad7b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he24ff2715e86fdf86506eda6312bc219e3c2e1c78e1e96c6735a00f24b48ae47a288791425d25f6020a305c96c9b278d06f0e1fd4ba342b3235872a18f4eb4893829dc8beb662230;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9319a1cc2451aef5f699b5efc3b4a8cd7c107e01ab5a72b61298283cbdca84e872f376bbbffde3335502f0ee5e71fc63bf12b4ea9a5aab8c000c5aded4e9475dd4eab5308db2d1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha05eddf33f16dbe641346c6135e6317dd75857638e373019b2ba65988a9a5b8458d6a054221bc9222090d160eaec8020b1a6411e5fe052bffed7d35c98330b86525e3645e8dff073;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bc53f7200478b6b1d9e65bf1462d478150e91c90aa5ef7f2c7cb5ef2c48bcfd8fa752acbe041169dea359f3a924713955bbaf4c8b21c233e7e697468f9c56e3e9f49750c7392655;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd5e78c112ab5af3325107281a5eca6d1ed423b15878aff70ef96166ce5b411115d208e2c6e98175da731333d466be79058ce3e0c70aafba76fb6ecbaf5ec6bf1639bac0540dcc87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfb46674f1856f91c7d477a9199a500e5fdc09ada7e401cd5ea34ec536c54c4f6f52fa4452c30ba53d23b7d0160ee0ef810510d7c20218f07a58d48600515702216686025d7b11b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a2781e288e0d18b9d2abc3a6e6da8318434f7fdf5fa6e889da680b2cdecda30b7a989e51a46c8948e92e8e61c28c525a1b4e21d497d20a9058d3d63eaf52f0005aca0827a3c0552;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40a7f415dbb18db0c51098701bd78e8701f7390b65ccdff3264ce95f2581ac099ca31ed67534a6de6c8e7b90999dffe78e65668d554cd63ab175a1501b589f9bf334c18119834345;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6cdc4a1dc885feae0e818516e4cd99b5a1389cd82cfd81e0e3f83945842d441e70baffe620f96d0a8f02a4796dd4e68cee97b07ba48b3e56d70bdc0063272a03b1b648f0c8de0d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h137330e03e2751a8345cb09722ae5d0a63ef9c1e1aec1822bea75a47f9c4b66f6cb705033d1eacb6a8bc8d256a2dad9037468e3c6d75930c1580edef3aeb9b0be1b5fd2c109df6eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff174eed15d0389e59495db8a48d5e5118a8174ddc0b1d1b5b16f53aea601a30721d610a56c24a6993340717826a24daa7cacd85e851aef7b2923ca5f7064b5ee1aeba473dfd70ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb17c27e2e9d6b94c77d0a0c7a7e745fa5c127f80c36c3f54b9c3f8935569801943df2b7d7a1bc5bb2ac0add5dc02f3f146c914d837431fa391614cb2404c2bb814e33c553a9d7b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3f411ce65ea9f18abb82bb4b054bed2285fc65d54d9fafbe3ef6cb48f72a50f83e9484b628d945d1fc2f7cfd3cf038dc4c68988474a7accfce770f8ef542801ed7747c9eb685c42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87c810106c24300fa4924f7c87256a607abdb9a3c5db4ca78d2b9018b6cdbff85f383b2aa25325de4f50ad82500573e0d987be84aeeca0120d4f40ddfb45d5ee6cf4e3e5743362f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f12ebdac2cb1fe6f851f0acef80dc2b10a71214aa570f555b33ef39bcb5f9d74de3b820429b5a4bf07679327b2da9981621c58472f89720c4e30afc963864de9db5710c80441f38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eaa9ce9dad04d90c63080a07a757126fbfe803e180491b43cc21fed1782cd77d1961ebd37285919bf1e1045395eff5f530530251e54b4b73ae39c72e90d843c7bacd5890182ff4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b6e9cea0df492b3827d049f9bf0208411dafcae3db32076232fdd81696f7a1b3839e2f2085e955b1c520873d276e0959c84f9eb71ccba04630ca1eff3cf1329ecbd463a01706566;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14add217436904b6053ff4ace07daec25c66d0c2eff5112dbe66333247a9a7ea9646f648aba76d6921745d5eb57cd4495c575de5de8182e985f787e8f6d16d993a824ad8791bfbe8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb849171c12215cf9d442cd46008680bd32560c2460147dc97e653460742ccac0f9f2086cdb1b515688df3967239e97e78a1841a917cd05e86091d18fb2013a26b565ec5369bbaf8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h712e04dcb47e2493602dfde9846d9f62f6056860dc7479704c77148d402dc24a8adf194c874438c1549e3b2b454145c1cf8315fab0b31a4b12011e0a80571b36d1d857156f61b739;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc18392a3c96333d702a5b22379ae8b1abbbbd042cd30aaf6d90209b3e7718549ecee937a6023c6ced07b96653bc9a2de0513656b102cdb621b63991ce84dfd09dbaf82adf36ae21f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc2c8d3e23f4f20dc2de7bfb9ee50dc891e756a0a63268f508697857dd07d7ce734fec905c4d750d3873bc53a50e5de25a307244a425c28dbae81f9a132632b370f5acf6d612c197;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6efbd1a8587fb1a8b41b1f7d587dbbdd7a9041667cc90d6bcf7b3eeb50b259947f0676df931f7a89fbe7459056f305fb4905630cafd018117fdca894fafae555e373d0928779918d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18a2d9a92527b46e7a8a4d0030b7241a96de085b3467348810af78178e2d51c6d16bf2b6dbce1727f60d7f6e14937b297059bec0fe0e16dfa062883f9b1ede09a2b85b2ee9b7d42e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89da99261a34260347d187d00d28f145e7665f904c6367ff01a42285197cfdcd1f3315f670dd7ea266f972019f744a8a9bdef52e8b8813be9ff82293e0d559c9e3d927203c7d4c9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e722d2920d04dfa1e462c73f28860acab33f43939eb74854c4027aec5a48e41680405bda79a9c231b8a6c83e3fb0343a3a90627a8c066bc8a6b470e2ba740dcf4dc8ca77869cb1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbe04137d2084c407443adc838018a635c42db79a86b3bd6d9798d667e4f49d3ba011d26926bb5ad5a230cad9e5be662a3ba08caba005d1fb7dc22e0d2e99659cf5342fb6e6ab2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e049f865e655344cbed2cf6aa64d2e29056f7432dd659f514e8c2b0805e4756c150b1e67ece0161435ddc984848d3b9d8e1e63d04e006abb94ea38cd762ef71d73eb147409c7a45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1380b26a4ede50332e447451ed0d4ad4cbdc77444b92edef46844d45936e32a202976a37e7debb58ad3c31d56580c82ce662b8914bb1c75199a8913db19f6d0ef563ddfcc3f85f1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3b94ce7d4ac8b2f3171f632862db66ab8d103fef1e9f69502fa13edf35eac0ef402a4dfc9e60952616dd925d59e8fb4c31b4b2be18e0a18c54c6878b3ff6fcc9299b919974eb2cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h945494b94c6b096ec355f1fee10a3f743dc04c34bb9d74190123a11ecd9ccbe3a48425bf9acf766e8e9e1f6d56157e5ef89b42963478dd02495eaa4d2e6df8b72fd011eaf4acd690;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a034c0b149e34c0b0503bdcd3eb6bba38377ac8773aa09408fe387f464f58d888191bd4be8301ec811daba59b7e6aee8491d64fc81a8944770262d7d466371ee3b9e8f4e71c3c15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e8226b705cf2bc2f3f84e9dba1ee6064991b46c549c2a9b6f91ddbabf44e8560d8bccfbe1f0e1725b3af1929d20869543f13870b8cac4664797ae57410c308a7c7073fe2a58e68a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7968ed10c7f4e3fc96b405c5a8942f06a74ca0c553a40259e51382cdd517a4ac562b5c7fb882fa9c4c477268862200acf940d3a5f31997fa2b77b3b33e27eb6f343e58b674f5a7d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19783b82ab1507bde01e4833fcc26dcc7f317608f3bf25048c2a4a3ea5866a4d1983ef361dfa937f11743e200f778df1739a211d6ff7c123bda94b792fec7a875e4229893d67ae45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fd26c3e3d2eed14f4c86b99b81029865349d9f6eb6cdb90d4121bc86abaf297e0ba3ff62c4d9b2916f515165e908aac02804ac013a02be1c543deac82d37226b1ea4ab0c0abccb9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7f728dd528be5eb517bf21fb79800b6c6d7163b5685d76a1f3ea7efe85ffdc6a9b7071fb0a6d4960e9ff1aba4dc144751253f753fb210305082efb4044406ce9d67f7b65df84369;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bd65b8103e5f567ba0cacd95316c3fe60c2801abc76d94da5e19b4474699263142c401997b551918d028f918b733a03792c623cff3173e1dec83d434399c0e6f5418f0c3a2dc808;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd1520b9fcc9d4389b5a921ce2e2818bee0234b98a4df8e284ea8fb2b2936de33586bbfb5e21fec2d1dfd7143920adec851762bf9e0cc1d4ef5e9d9bb22d457b0747b658ceeab40c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb265740dcca07dede03ec39e85a7ff710900866b3b269ee7591ad00743eacd17a157c4a306deac3def52ea584bd34e0ca762ae5566ac96189494794f8b36eb9cf8c4257278c4c26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e2fb6fb6eeebb26e5679d3d41ee72c65a9c6a1f4bd4a21b7f3aeef96e67cb4fb607e2535c31e41e90e8203d0f2c2de8a598751f4002c6480a5aa720c3d40b1e6e79499dff43bbbe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97e234c88957853b5464c55e708e81d95ff4eaa97edbffc3e084dda212955cb6e381a12eca140d63abcb479865bbbafe9d836865c8e1a774a3bce2b457697798cf7dab8ff0c8bf22;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfab427940c91437cd39601543c9613071f10247074b87286ed44cd46766faa4bb9697773c82cccbd09dd989fc34f1fd06a106f3add14074405fa4ee480cc0d90c34445fedf2c79e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ae71ff4b4f2fc3bd853707a18d98f17020eaf0376d57102e1a25fa404a2520f36317e4b4bc2eaf29c8e431ff8daf57a974d205301c5acb90c5ee7f7a7421a9693f81cf26fdd748e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e208a0be5bdf686f7c8b0b8dc3ac4a14988920e9e8d496ebe303ae1dcb8d3f0717df076f25accdd35fd45b8d07742fbc2b4a559e2954718b409b4df096701a093b8e21a70dfa8dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had39a9f27d88be9d85716d95e9e20c3258ff878928b282f28e1f3aadfac82dc27b645daef4a0719bca61727352f91b6b6797a83658165f1a015213f635ebd5e2d62027dcb909bf97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd37b2221191639db80e1d050a335ac8d6bd9983604e757df911566436c4a6291af3fb44b72024f9ec6081d501063069648e997cb4c60a535e54ac3cd157ca6a668ae9b8aceb0b2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebaa31898075c457d739d1b1f6bc1438edfd114b27eda6f3d9e75f9972b108717aeece4553b143896d39775e83df51fe0630fe9a0bbc068820ef3ae6b8de00b889e039cd78de1ca0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16f221895030361c7a11a6d4e9274d30b85935a5adcb0016c462eb53ff87826a56e2dc2a6a9c8eac30fe842b77a99f52957c5410b9fddd370a34348882b326d0490774849d7c0d3c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h159846ef62605bcb5c24d58a3d49c015283da57bb7f17602c7f07718d6f98dbf9411b0022671a0a68c8bafb6e56a22611f583d4c0724a5ef0a2c034e0da6d30272a3c0192a7471e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d643a962e47b4e87c0b97c662f436c9bfd41cfae4f58e78265aab1ff3c4c35cf66af9f5d725a4aaeb57f2c4c546c327067ca73d07b1a5384b6ba62a898e1aff56f01bdd686c254f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd629867e0f1aad050444cb83d7e25fb27b535169f4aa238264295f8700676fea12972cc5fdeae0dde4509771b5baafcac65d8eb225d8ad8380aa230376d99124efb758162dde6bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76abb17a5ee617a7dee2e76245bceab63b510965a6488e3f7d02b33f57fb027dbfee9827ffb243eed03d3e00b2f78c51534d2cd2cc4763df3b7981ef7cd40ac3febb718520d3d06d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc23a8e7c37e04fa48cb00da101be5c84300c83e9a90d5a93ab38f6391b9387300eaa2284e35e4a476a21f61161119ddef9dd2dc159cb6c1cac89801c686f0de27293ca6cb97a99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91945654b7a7b0869d66e7f9998b080827769ebdedacd5637738bdb76b5b90be57089964929b7cb7365321091f1f79173544d8acc47ca9f04325a716c225a70c8332477bb0305626;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67e1b4e4d4e2521c6841d70e6e2a2dd83b9755f6c0293b4890edffe62fedcde24924c57c93e79606a958bc01df64a3effaa4ef07ce0a0bf891c8e8995ed8fe4cc66b0f293a0b678a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c34420ffb829a9c0b25369fe53fd1a873a545da34fb5cd3916a06775bdaa220e65f6faf646ce9ce9c7960ac48a371c42fdcca4ab22688f565f566b160a2e14d7892e5c936e43a8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e7c783613d9a158e9846a10bae1c0543e69ea7dcfc22e7974a5794d3b02395839cb052a1b3cbeef3c1a570420fa25c426c49b9b22ed1adb582932e36eec89312edf45620f72d35b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h552fa9c0275cb801b091328f7253b5752e168012bf388f4409e4874b7f21a877991ea1b3a421d960cffb12240a8d126bca6dc872eb077261167d4917ad0de981a3fc7693061dd4d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6c23e6a671f56fbc58adaa9000b815fe57697eefca81be6b4c675ff106a619f82868aa09313397eab0cc21ecf6d96ed6c08e6e4b4eabb28558bd1464e7aa99370f696ea9915be3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h654780551eaf2184ee5dbe460e6ba5035a3caa2b69f16d1c7b3af0aab57c4c0f53c8b6b41de5acf64f7f8234222bd039602883af5e59a2f69b6741937098589dfb38d3f6691323ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0a3edd4b2957e21d033e9650a6e234ca6fd87d52fe2771357d4a9790ae3611f23fd16fd4b5107a28f25c564dffc66b43a0781953119d9c32ab1d759c2fda34007a1bc81c78db24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6c3723da4f93d5c11abb144de3d8e32846b76610b88fac3bb28b7b45fa499bb5ac1a50ce1d4e1d0431f66744d3a5c04867aa1d29a244bab19ad9e1fffac48489c935557bf34e2e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67dfec9723fc7d7a707653723d30483379040115941ab66f997bed49d5368e6581e45318aeab56c197109d2e89caa3705c6ab97a049c7551514bf7247898291b7192816c2b7f62d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7777ab9ce9a344c5b912ade94e1683a7f0c4c261ae9346d7257b4e0cc86f245c601b103efa49155049e25f7190ad9e85e3cf6db1d619a1242b0eeefc9c56d05ccd858730a366453e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90d9e2babfbfcf79e486497df783f5f089dff8b4bda261c67c80554f8ab2b14adcaf943f47ed01c27b3d028ca1ffec24fc86f69469eca42b78d4fae075ecab28014e9c3e6be3386f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20a4edc6c07d0b39badcf020749981d9096dc08d10f15f19af05a49f669815096b3e052a86793bc1af64553722c9f82254eb53adb54fa9fc26c3c15e90abc3c439f2c696b64e346c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13be3ad6ec78339720122c33a1367bf8034ac995a87bd5f0104f2abcc9f56700edece858d559140486f98c45566408bfafd72be18809f57f1fc1cfa260fc31f532d0b8ec822b47b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebe449ed693457896dc516b45f8a1931d5eda977dfe4ad3077c4dfc4fe15ad92eb4db44f39d85a1b458dcf5229f51408cc69edd88b0e17a46080238ca0728652f36c639e634e77f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcde562744de8ef7854a317d6c5df0da8089444517b0061ec9bf2124a9210f3204ea1667a6623c09badc68c1bbf00a168b276b47160324ee746c5f3dd89a6ba9c9d7677f64294b6d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h105fd8f63fc9ecf5d2892a974d34857ae6055e2a04da42c56099c69a1f216891618b1b1362bbf241ec0fc0ae7814ce7efc9c2ddec882928a835dcc68f5f921eb71171d3438bd2e6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fd587f0fdfb5e1754c66ba45b7960c3f6739f7c3504240d6aae7822361a1b521876dcc32d69d1609bed1855b13ca99afbb5035d3d19e2b2b7eff84fae587d4b4839261e287f8c66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34e28e7301e8b12171ee6c98527afc39513cb96fa1ed1d68916dd9b2b7444bee1ee2a588f6618760cb9bfbb5496dc924b4bc072069a62fb252b3d0f5988ecbcafbbb41394e211aba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18705b0d36a37fca8cb856b63adc7695c1e1acdc6916191c7c3d4d5e1f297458fb83d771595587be3d2b190383322857e128172f5c28c43d177ea4caa71e46db086d21ed755b188b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87f47fc9f6b451f209f0fd2932c17bb8b5c2857726e58e85abc4e5029f6b01cf21489d8663ed6e79eb26b023985ceb7a4ae42efc57958fa8ba4c5069371353fa0a91c6eb0bfbbded;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdf728bf797c10907bb5dad0c55989c76d7408c540985a457c3a6b5a3206d10b4ea3c16d9b7944f807d416fb079fd2a9db834540c0f2c6d62c6e0907b6f63712a647c4369c72bb1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe6adf6474d8a3ee81d328a2013fb60b1bf05fabcf33137195517d57a4fb181602e0aeffcc518b4077bae3f46571f2b0ee4cd05aa41012cdc2626e3cf1b969c30e3cdd4c96799d2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82978b1fa9f7a939957ab2b5a9970e1b9778ef095dd88cbacecd4f25371447c7bf3044e3c8a809f2a76a7dd5de521a66cd90ce3c5f4393fc0404962bea6931509bca22e997b92e8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6c6b944b0ab2b06df2b954124157736ed7b9aa6d4ae1578a7eef91fc817a86e34d8b512bb6579f8a9d704ec732461847a697a3f7c6d287060f90f0d218546b2d3f2ac06fcc8951b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69d44362f35e36fd8fbbfb7d1143da53ba792d5913c9ca8dcae50f3cb78e909b4b101fd3f86d56523697953d32757f2d05798774907d3e389342828685be11e1be2eed0a3c784751;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2389678078236090dd0c28ca3331c6417f2c41add3738068dff2c2da73eeb4d827d72a8af11f876c3da0596646da63e35bc17644b0146cc62b1dc077b4d8cf358938aac39d8f31ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92a1a51fa677d596f3371150461c183445614c849dd1456f204a8db0bb63f7f4bb45468cc548933264e53fa5b3102fdf589785da5212e9b0a3741238ff182346afd66fd9f1618777;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1cdc2edd6061e01a99dfd16f78a8b57da3c4c5805f11266664e7edeaed26aa1ae3b0ba5d299e8b43b7a700f04c3f304446d56df2c61dce4b53e6544307dd8ee56bdf3d34497b7aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34569c33c6ce58f1c610de63bb020b04bd5b63a4303e4e4990ed3ed62ae372b507944ded922375228a6d56f199a49bcc730f9ce351b353b13ce66a39ae871e6217d0bffafcec2aa9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d3bba49586146336e9c3a164a6192870c251c57bcd992e462bf12e6c02255caf41e20aa86ef947f14285f6ed18752e36359749f1d3eaa55d593d88e616f47041b9d5c5e5234b7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27a848eb463624e4c5d0049cffa9c9f56a59fe34f908c79d4ded3c46fc8c7bb844a540ebfc86c4d346069d3897b212ece86e376299531a9bee8ef9b021d23f3d3ceab3562ddfa7a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf536b886f8b0c819a72106e322cadc542c015b15f5da656c84b93bef39ed6bd6fdf01bfda9645e6b595e941bc4261e3a28a1fa2f896eb7f87ed637fb3654ce96a37b2f7acfc1bbfa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h460efab173eba531387b8f28e75436fdd6165924acae1ad5cedf2bcc471d7b645f241f0232442ab748fbdfeaa1ce620432c231ad288efac5cee9a810b3fc973993da27e36bb67baa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h855fe299fe4af783d15b2576f78505c8254a10fbd499017b9decb7814588f4071821ffead82ffc2e253cdd3b4624f8a41b9f240baaeb230e07df5c1ebd9d2051e41edf5e79720229;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87766cfd0900ae8ba9be9b7602638a5d29319f6e771d3be43a5366da4dca19295fb3a807ebe179f386c2fe2f355b84608b176e78b209f8317a8a7f0776cb80946b11add1ce6e96e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he08bfad8b612764f0fd3491f08d89707b3ca2fb9d4aa15cd1e48da903afa70372eb99db75cd39794b613a1742e3e8a1afb7957ab1936eeb02a80941f628fbd47daef7487f0d9870e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b10c33ca45f1be8d5888f6dc48d1bfcf7d119013cdc5bf21202c1297ef7e3a34f7f5cd2963bdcd6d064691a3753f4f20a19e039740ac688dcd8c314b8b5e742566d2663b5a7088;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b0e3290c8d26f4ef38860814ed8bf60edbfe89bc8d6ee849865c6050f95aa9a73919ffc0192e41ca668ba6ef3fb8b78b962bb4c3c16b6dbf2b01aaee01fdcb38ced03c452de0325;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc7936f22ec7715d9aaebeb928eb9be6126be22f0d18f297f5f6f8b99d7d9975b3d5496a401701569d20eb3c22dc93f21ac0cf13b06a06a91ec892d10c86e8a37ce3d3f6b831ee29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6a1c8f2517b1a17f30073fcbd2c9ffaab87e333af557e017f2d82fe4a159556fba7220ad4853dad789e17cf50e0cf718b6f72f70fe7c048f78c4fd1f7a3fae5e44aa1db015e0a69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f71b64840f18e3deb8d9b87d57282ba0f7a1e83f524111f4fdcd022ab5c9ba4812d8da001bbc1438761eb2ef92959d03cd9b590faacd24fe54966038f15f67c2236cd1c056936cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9b54161118bbecbc079db7bb7482aba2578724f5e0196761ab82b0033923861d6508debf92d202f0d1705319620900ab93b7ab80876d0d5d5dbc39aecf085d208bffb0e72bf8d66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83045927e8a746f4a7d9afe746aa376c726806a9c95728130bd1e90a1103ba77fc0d7aec41e1b24df593cc7872147ebb389dd8e07709a4ef80aa546b9c4db045f06bc90784e73b06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19aece0c72a5fb6175fd94244121f9ce1768747e5eec943e2075342957f9a5b81f4c604466b5bbb703696cfb380bdfd89c93563074653c7ebd3564b0c1b4e9ef8935bbf21ea0f348;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78a9d1393fdaa575ef751431f046dab39ca89f64ff4db68a2b0412fd36320cf5003be840a54c0ccd9b856da0fabaa5f4564dbdfb2d4c250b6df5f9e0cce6513ed3c962d3caa5bb46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdb8362222b95e6b37a9f26c7a467afb06e9e9ee0c3ccda13be4c77dc171b45102d847002283101ebc1593433a2bd4cee189faefc174ac190ee364b79c28d03ba9f3d5cb87e44a80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32aeb5bc1deeb498850412458c1dd4e69f07573530b145df75599c704e365a1fa4286c7f9a6cc69fdc8b305aae3665071b2804a5a8260a5b73f1ad88c1b8e891648d98c5de50c02c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e342114cfd291b4ca78d7df9441c441653005be99b5bf7593b35f7ae2ad3e197d45b645baf0d759c5fb6c5173d68f72fc3c5426aa39c963c9c2fbe1c60a40d0c917f41471c71939;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f5c7b9a81d18bad055f3ffece7488de7532a45ef695479982b43beeb10a8d9851f38418a1a208d8977ebb6f9ddac356154a918e115dcdb4bf2eba5fef2f37caf3510ba1c5484b7a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82a45329cd663b7e2a3fc674c1a30897a0e87bea6acf5c6bcf4dd2753ca8657b56edf52838a57846095c43b0fa984910b40cd68be4cc65779814d87add256d40b419ee2966543fb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1aaa17ffe29ae32de061ebe9852b2a2c976075744c589319d5191040cfc723a7e68e5cb780dd8a0d51bb4a543f461cdd8accbb15c5bd6ed5ce477a267a44e85c4d8bf24e55f5614;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3df5f19823da2d32115b532ee84c0faa190cbcbdbce56dd0b7a6e19028018054c6a396bffd0515b6831dd39343b560524c7036118432e95752f01fcd2a777885af209379afce1de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc83b4505a4f3d3c886beda06258256a7dffe3ba13154680295f8c98380334e6772dad67f1b4f2f9801bb791040560d4980ef1ce19ef2d039421304b88ea0c6ae60c144028982d495;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd29cadc4300ad67a629181a23e497bfbf28488b9b54a9e10fb42bea74e6cb9b50a945e0a61dcbd095c4de68dacd5dea7b29292325f8cc347176466dbcc53b3cd7475e497cf5690f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43d5151d14472b8f31b53a3e0fbc164010f7a9f2bd96d673b7820d1d8e9f4206804e0c94efe115f777642622e3cd6764169d2a037fc5cbcf0815017e2954bea25c7550a1fbbc3efb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h559c968f45f2638cbff6afc0f11da39cdfafcd3744baf907a8f71e9bf73d06acf2a7104b798bb64d4e8a932af7bf2ad534ded8db74b104f584a1110e02f418b992b39256f21ad77b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadcd62851c3a77703cbcdf4acf4feebfe026a708f07b5c48037684807843d93a06a7ba4480b64741150e211853ad1e062f577f9a35da59c85a4ecd830cb656fd286be6f9848a6561;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd38358d5ac474caf6c8fb66e566c01b89c1f128f4f268fc17392574f45291e1575d757ced1d246a06d3423b48c728852ed21f6cd57ba199e8259fa7b95e3b73a0acec34a1b4db706;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec896f54f1f9ec801843617b1fe31d1baade36b8eb0f0803f54289db2c5778c340465e5d6ca62f460e0735811dde55db36bc561845fa51d8943035a6d85aa04246c1c98950ef7c8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he35200d49280f4a0cf5a900928de00a93c01f3a8835c6d5d93028d7afda707b9ec2b20ff9c77e8c4302a6881a35aa7ca9f798c881ff0bf8918af2771d4d5cc1d810d88a1ca114502;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h966b8d459115d07ec7dea8e3eeb0759042615691cd9224890b016595f6e6e2b8ccd4b3be831342943c87f1a506edd90610cc15ff912baa31d93bf89a762c379b9a81725162e40027;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42df1fa8641cf6d555d67059ab66e83253c6033e32abe8568b8b9c2cd0a229cd8514bcf14bb12cf0a470f270cf1226f2264816e0b3689832b6f8c2f61139953b6a6af2e7e081f58b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda4208660840a8acacd1522c416657a41ebee5bd58abf2bfed690b5905fd20878cd7feb1eb35b8b675de35f8885aecd4b14d0a0146492813b98a0defa828da8ca64c1e25e9b409ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64d31a4eb605f0eb8062e61a45c111d963d1c838c838afada60a8c569e956b0641b7aefbda841dba83a669e75dc1d054d3196211404ea2b5704ceaa428f2b5cf5d62fe62323d6887;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18e70b43f2a859b43fb3e5ba83ea5ce9fd5b8bd20ff34533745a9254a46b319218577497d1f782ca85e931c69c701a2020ad11c1a25284594fb8518677577f4614e77290bd0e22f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf1575136169f30c7fe7f9ea8c49e6ae10ef81f53fd6067833438cd1c85543df0830b1b9b5a0fc3f1c231e0ddf487b4c3b20507be75c20450c32e2f2ee0d61a680ca177745ba6132;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cfaa122710d81fde9d5d3888facdfaf23aeac111a6d19a1d2dd989e82cd86475e3e13b0e5deafbd38d267052543f8e82701af0eb9357140e7a51d1619aa184648b13c256ba8c5ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h830e3fc44cf416d8564421603a3b06953573dfb70894836c6884f9ab83b3d8cf1475b5a7420b91b46a3f9dfac260cb86a6e6fcf2315bfb9057b636a6aa3da66d3b1cb75718e5957b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc2f2603d9a4c5b27f084c66890e06efeb2837357ce23f700b1ccfd306f82f9ed2fe83ee355ada48e4b48e951e656cc733f1cf1249b1259cdb12c3c0cb7505f5a2941b97a157f88f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7182b97014df37aa39441e83566d4d55e2026fbbb210dcc1cc1a82a59c5f82d5e12a158dd28986d1695c35877d25761760c32028e487a8ed0a2bd1f54236fcaf37817703bb0f0b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bf0cda29a01ab1e83587fd1a156d1940a1bf8db1892b16eeb21ddcb53bdf22c732dd74f9914749110e0221da9519bca970df564c62d04d2989ad5bdf3dd204b9f8766c05e6acc76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44d464396bb303b39f9ccb5aca8f2d77bf02e81baf7290fdafa46899ac91dda9e7ef62299d90fe987b5923cee0ee87702b7666ffa00618d8608612c53fd9e7fa0377fa35ef60bcfd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2eb2cf139f074fa3006c16ba6f0272f853d7fc21ebef419e0ab9657abcc1b81117f6c5d88da68b370bce79eadf0aeff3f7b2ca48fe520845b3beb02eef58835834ee1787ac2e2a9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec0f83846c21b82947abeed792ed77708ef8a80bdfe4001cd48ab691eb2842b26115b201651b7932fde64b94d32561caa3e609c8877be8b193141a9f7998a07458e63ca25417abc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60cea4c84277cc5a44fb93a82034f24c39b9184477716825687d05e9889e2b7c5458f76afe7d6e8bfd693759b1914a6ddfa459415e6e4bfda2aa1e910235b747cf1e01fffb48c26c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1ac7284dd155fe8971f7fd163e14daa635fb59d1618d60f2d122a4bd3045fc38f96d7842e6c772185c7a731718c581203c824eed84be6f50b94ef0827347c30450485fd0a791be9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4d261d75efaace27274dddff30ba197b2e5a24a05f18b578a0144feae3a4c29d81d5740f8ee6baf8b762fc7bb026b467e5d40df6745cabf488a96f9fa3656b411fe3f3e80c2340f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b8e9f5ed8df3c2584bb68d820943f670e7590dc9fbd2b5bd96010f710eac5610f9bd4480adb2941a7af108120fc7d25697548dedea2ee89ea70182f61643f350329fee361d06e95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc99b0051bb9011dc17c9cc6ef8fd023d197a8870860e0923f165586740cbcaba1368729826b796f0e481272f186b336f2c7743f33d5130b1b8e2744c8b0e6ec3b76911db4878c191;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bf96e553406d16bbf66cb7c529574058a58e76856b8ed9c0fce48006a0c6fd594cf6c52c8b44586cee75665eaf256b936c24bce0ceef7767aa14e20b821434f43bc98bdaace6253;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fa3fdee63bf4067b7823ede6ac99165765f0ff5595e1d825b21cfbd1203dee6cf5581b099127d1b75fa0326f0eefda39cbd8a879a68a4b051992dd12f05867505a6f3fe155e17ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99d4de9da9dfc077f4b7e3f16756d6b9618523ef44fa869e058a556d935af989c962a5b8bbc66ed9acfca4c7a9059001766a834c2e08d22ee3711d61fcd333dbff784aecd8bc622;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54e6dc4f8d61bdfc58a369ef320a2178b7a88f0a15f70520686e311e4f83991881af3ee02b5e09bc4488d559e10552fd7bf3000640b91c86a94fef33eee454fc5441320dcf0a7bfe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f783b940a04220385836113878b634c5168fb4e231d3b09a922dc21ef2550113d80285d2e3084b58b8df61a6fdfcf61288ef0d0218f1931e72e2a1dc3ad939dcd16b7e1c5549ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77173bbaddc996d29fd19fe2557b38738dead4ab873a3361a8a1a7496e03f400e81d3f5def2b63212cb323251db14bad57fe37dc6ddcd03d4caecc3b40cc05f2c14f816cee42a568;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he48a265d91850caef66cecdbae19b1590ee0a85e9b449452f7e15169b77a103c01faa1a02b50553293861610806fce6c6f3bec9adf5e7b6380681969a99a12619e8c586f3b52b31b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e7daa4b1987e4fe5d3e8c9c0f7b05ce698df6c7b55f3bce7c3359394191c8e8ce060eb8373bbe8813a0f97a3afa763da76b5588aa0c10df29214cd893f33ad6ce8c01e4a0f4fa5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadd3f4b56f2964ab5ee7537750ae8124f8e0b733f86bedcdca3954336536e8a6b9f7b35b7255cb113d174b6b381dcc227b332e2e28aeeef95182afdb8bc83445743afca6e3727dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5deb37f198384a4b58151b934ba98ee1e6da21ccae452e42d427f3ec16fad08b57db0da8e6014ec7f7e36ad29bb77376b8e23ce0e935547e461eb4ae90918490f0dd26eaf148091;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8242c87fbbe5e8740d6c47e248803dcbc9dca59fb26b104f6cda8754acfd7a97ae71a37d4c9fed42478fcb61afeddd47fce5aa73c3ceab37660f3a5c12a1505cc55c4277c3a0aa2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he66ab6ef48fb812040e2d560ee11ab120ba25d1e01df49bc2188630316fe47d71bfe78f1084f88f5667d5861bfdff58d569eb26f404e582823a81e8d88861a703fab3d529b305690;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81cfea173f2a7709c4fa63a399ddcf33fd9797baf08b29e98b199a0827cbb52df5c4d2d05e9aca0699f5e8830af9052acd7c47fc03ac6d47a9a6cab9d23388300892229f0a2b3ce1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h689e22a30130d0de4f53e9421c09ceb2de79005bf770196bd6a463286d754d6ebf52b0f45876c760731809abf0831d4f7eda7c0e4f839dbfb07a69d9969b14bb26ab4daf8b5590b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4746eb68a997ddb30147e78cfe30986e8d3d7ea2c9230d5eed38955d48db72595ab643ac0d4efb64dd2f05638574a79fa41b347b8b7a9ecebc00222c6e7dbfe879ec6d1b3ad261bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h843bff9d8e6872c643c4644c6e62dcb2df2996bb87b78cc4e031bd393f70c058d45b73fc1b68a3c35e3d8e4400925345486b7b69a45c5ff0bce63bd727964dbdbf35f262ea418e43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h607790c30e224450306ac6f450eb4154d7b2e9708b88a5de4c6e332391dc295d4199940b3922183b933503c08cb8b74d186769299c745c5f5e04260b226875f77e257115f8a51452;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1b68b1c394279ea7dbaa0c1901aa4bdd3123449ca76755fde91d2412b0f0734222eb493300e31c425ef5a4398dfa3c4d1562ce9925b587e8d04de14222b8f9ef5d2ea875e3c7b5c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52304c02199349f48339b1dda59217926390a065577f0a6848ed33c2ffb9b8709296748afe58592bdcc55538543267f52f04bca42bea827ca52bbec284081c23fd880466c666ba31;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he35f11a11ad691d8b97ee82451734b10eb39cbb256ab50250d80c0bb4552418ea65a0f9eb8e6ac35df9faf9a821334ba8d0560273b97a62b9a5247d53ee43b9f406c324352118b8a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha492d1cdcec9855db53970d1cf840fb349c69ce900f90b1d4a3ea91f97e4d02e9da284c8f979742f278bad7b5faeb63e16830b8d455e16e1127aaedc2bc3282b3e1858ccca44594c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff44a1bf91476f4503f1f5f085e55b23a83fb472252e33a54592e75f9ec5f986fd8df84eb9005bd72f0b20b0bc463d49399734b57e5887b9526b736635c3694964f57ffcdcb551f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85edcfc6ff047365574d6fe15d3f18ac3330cc33bb5b0d0ba730f6f0feed2fb37836be514919fc08d60bb1ab6ae3bcfb60a4874dce8734e01f5c9f4883c69bbda27736ac30bcb7d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b9f53e2127308ebe61232058568eb76dd9556c0607988a3fda83c834cfae19fd464d7e3a2e23ecd8048c685b32d5200dc673fadb2951359d1c263df9df6b5ca0245ab508a5dbef3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27816fe998614dd48948d53b4d761568a4159fa4ac69a36ff85f7bb4e267e939f5e2648d67eb32c7037d2cbc3c6e678753227850e6f4d277366b6e1ac7b8bfe4b81683037e8b0a8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2eb423b878c85c830a0bae43f393030912a0a929146401ddd0f69f464df13901f2af001d1edb0818648891149b6a2a050f256729f97292942b7dfab23715a3f104740ad63b94357;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b872a232fdbfe61462069159edf1645bf9afbcdbe1cf61ed5db1ee9b326ffc95f444e64bcb2d3c187504e3e6a7edfde1a774606d9b985e0de95836060493442b7ab7b3b48b2abcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8df00a8649819ea8227512dd895ec584d06a5f71e334c3c9eb044b4acced16070cee8d7c2a14562a4f0288f0a48ba6daec955d56c038301841f465863957ce9101b523dc8b04f2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0c2bd054d6f3b7348b5a7279e7b6ab1ff30368e212b927fc34e89990442bc8c0862ff550a507373564c4a391fc4ed98cc74f0a94d551440feacf9e80fcf9a52372b045716384743;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h217b4f6928563d406548a3ba5d7d9dc8ccf842cdaf2017af3291a67f56d377f1e747456a3c7f34cd754108e0dabddaf7076d1c8dce88dbbf4368eea1cdf37144d0398345c560622b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he794199f870d40cfa85888b48b77663352b1726d44733f7bca1c18c6fcb19c0ad181bd4c6d353c6ade52aa1d4dfb8ea9c3e7e8e3848d6fcaac4abfee45504a6df5109df92a2c3073;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed2a2db70a1d1c13db09bfc7b3fd94e17a80ca8512a31b4a817b51ddd975616e0ab66284af8a32f639f769c16c6a1292f178f451a4c3792dcffafbc55b8d4211fb76d052100f7a6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1e59e1269e97766ad570b308bf593446ccac573529d99ca0b4e38af4819011bdd18b63da0518584997c97427e289c1d6e5ae050ac144224d0ea5acb888467594301ca3daedda0f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1657f8061b1340d8c877208b28f36b8894c1037fadfe6421d16c86ac346dcba17f5df162356323999776bdf0b1d2e668ceb0b4c3660661368329b77d655e98c224c48ae5f8ee37d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h973975447a404bf9b79ac5f98662c6df9f89bed245cbf3cce32e5e0968de9ebec3d16eecd052dbd2e107a0f28b01a689818ab27c0b80cb609be09bd9e7e23bc102e8b09a88674592;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h169ccd42dbd193b3f9a1fedd77f56dffdc0e9932dad2c5e21541b0890faa8f4f7d8d366801ae724e7e5bed118ce5789c09d7c012abbfd509919cebf575d344b7a95693f5fc59e57c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25df03f9122b6cc081e71702feaae0fea404602879d6bb7c190c51240f2a0b70e8e41056ded97c8191f81aacae4cc51c6ee652f0dd610415e6efe61645e7a0b9497cbedddda1275f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf82bd60bae030d1b28c68a2ab125ecf824a3b8d8b1b555d755959914e48af64db57e5ba882b55a4217e868a8929dab867f71c40ab17fc14ac154e5a5e7d84cb26f9fb0b6d12834f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f2d01971442692bfabed0514f976732012eec3b0f267cf6a28b09f9cd30ae83ba89628f735faf471e10c7cc77db1a5c9d0cba1e79a7c07e9ec8cee5c4de737cbd4516d77b42fc04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99dabcf14a39505f0275a1879c8db92ba9a725e1ca079e6aaadd180a6f99323f7a6e6f6f3bc16be7bb24f907b14073213594b7e476ed40d08bad465efecabe4e629fc12a78c4815e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb67518b8828978b80d3834479b031bc5124820ba2d7159e790ccf64bae8dfd06e807c1f6ff5c584fbf40dd01663f9492d2e14c656048a6e8f1b7683ac056be29011c2a8522818bcd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4af2aa8a145848cd50eb3cec402ad36d0fe0cd3e0c7f403f2b2029e7671ba0e23dd6b507a1aa9e775395cb58d8cd2928482c4ad02394e6d65650eb1fbb1eb1a6491f3ce0a598ae8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd53d9c4b9b2c26c6b322b622089aa3f2b0b9877d038ca00967bf0a4f58f942906f98b47711b16089cd567426b155518813427e392c0b12bfb466d3e4697ee3bdac75fc0137cb72f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6063fca856f89aee0cc4e69d130b4be15c0799f8b14c552b9dd220843fa1cfbe46c801ff448902858321af6f7cdeac63e859a7cdbb84cdbefc44a57ce640b20014963dc64f5a7908;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c404266a62ab4f0aee2ef372bd661940eee5acc9af48a639b3e22da2b6d1a8f5aa4c99416289bcdfa4ffec5e31067d434ed0f29b198ee68cff19042c7b27d59a4f4998851cd7a15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he25f58625fa7a47a6f035aa4cb298294d18d85b01bcfdf144e6aa4ebd410f41e8b8dae75227655d249ae82e740b1359db29a371091ec91150dd2991c119f034b1d6ba66546c86566;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4961110a4cbbc68f7c888ae7ba9bd51b6f27b1a89de88b0a303c3c88f77f37350388db90cc3736385a401e5625cfd0cd93aac1739a6f1e121d3876d375edea69e92d43a6553ca82b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66175974298dd5ded1fa15496da29756559e82cc4c0c42b1b4612605c16422c118c876bcea22ba7fbe67ec231a2dd512d4a292283d6ca426c3db32d8571c5234498bb7fd5bd6bc92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha02527c1cd38c4829ec36fdf5d8698578b0af151ca5bd1cfa21f31f4280630d8d487d0bf46a2a995b843a364c9be5ac532a3bacb7380065ca7d542ce373b28a6e6f1478f476e904c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c529c63f7ce09a650e97128702bd54886d5672703a3787fb9b8b0230e26cc322e376dc24fbd72628f8178f0f23a5a62d680dcb8bf26b903116289959aff87817e703195c960b8a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef77bebec16f7a4e67d2cf3a780fb84f1f85722e7d11e597b336e670fdccf805149154a067afa66177215979b5a0962c052b6511cd0bab3a121934f7acd68e27d24647db0acd6fd5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7158c51782b58a9691d9896614058bb165d83d70f29eaa44a064ce38fd0894fcc3d39fd126f084ded826996a58031c382e5fdbd166dea66d27a0bbc255e45d92a2035fdb4cc8694c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e8c9622addc2a5bfc46b8ed681570f72bcb8828ea71d7c1706dc2e0f6a35418d3b88559a2b4c1af01cf3bf0dd11e6e71691095fd9152f1609c4736fb6b4052245ed7d2d70941b27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5b579426790f905305c21b49c71cb402419cf9b6d53848eb495d297b91ec5f3d50d22c50e2074d49efc5c8fe7e1ca60e07ce3942afa06101e1a1f2ed45732805d9e4e4d1f4e416c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha21477fd30eb692aad63995a825bd15c99b6416e48f434a42adb33ef1da72fbb8b60c8bb6175ca5ba1917ddb081740c436fe690777bbec2b508eeef78cb902b70cc8666779bbf5a9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd61e1ff62842375b2c5fa243c2d76bfed7b59c268f94c2a79db285026ab071f2d48c09824f8dddc2b42e6a3b28767253e2467ff4c66263dae994d2aacbe4b8ea8d9f69532e860294;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea164d758916b2abb2ebdea6f6238cc5bb6e2d3f46b0c52cd7502abe6d70a7e3034152b10ce1fc77958a194da566556c856b02c385cd45c79ddece43e82e7caa227f3f07a59d1a31;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h301101f9fdaf5dd94f8a412918115ea0542dab0f0820b4e985179990a847767e6c9f2c6e2004b31c2ba773b32645fa6927a09ff660098ae098e3427d75cb09bb0306965524b7109f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc8e290a54128b015c3cb3bc8521aa1987107208c3a6bcbdfaaf79b7819c2c4ded818cd8201c7457d3d184ca6225037286b8788fa546ff5f47db7911f1741b99a7b1f26c95746d91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h162693affd2fcd1e20bb7d362e9d70873d0717ed58bccb58c2983f2d1f91a41259f2c6e02b98f2b18a2715164cc7ed971cc37ae9427b74fb0cff95036ab70c4212deb299c98d8f7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd553ad65e635ddf2e49f1d9166c18fea1d9a27102da9578cef62b122e215081ef9d6aabf22065f96d3b518a4a4c1e5805e218b7e20c077bcbd975b48be777730f3484cb01e8338ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h692212ead18bb1b52e453ed6eade2c04fda98ce278d86aecee8136c9de540b4ede4a7a268490d406020ec9614bf40bffd9c93d3dd347ef069b258f3869131f7297b14ef415594fd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ae6545bfd4eba9b709081075b061502aaee0529cbec46507497206a9294d2ad94bd0388b6d8a7690720ac36a43489197262673fa2db8c1d3fffa560a7d30ac352d3af0099f8920d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52431a251fe21b62128fb9b4d2636008f4dc9b8b797a61f0cf69a227e983abfb85eb973a8b41bfec3f1a2f2c3c02a1a9d650a637487cb16d566ac8fb2388ac86875380dd17da2f58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5166d064e1b412bba63065724f5b597d88acd5fa491500fb65c1ead3c0453b14b08547e061e113e2e599fdd22f3c7bdcd07d291712655b47a1dbcbfba8fe97a629589ecad83c52f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80ac07ec02ac9773a81b2d63147aac918b413a73a9f0852674aa24d040b170c820ed6b74408405a940ac1391e08817c4d91631232ffdab24ed2c164b4d98269188bccd1a2734a70f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h825e358c17f2db5d9ed8138b411267c1187e2c7d92dc73167f813e5de3c32cdcfa120d0a042304d270be7ebfb3332dc971ccc904f3fdfdb24b37e01c169ddc06fc8e740ea05ea5c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1b2b392e90debfe6e7f131422268aad8b9fdb6691dbb894426f470197f949ff8a529986e8f31b4a907faf5b5e5c2021b6b963029026dec0db06d1d71d0e718d02f2e04fa86defaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4941d79f256ddb01471773c382ea8a721bcb6de533bf2481ac91b7678799520f8c845b21cf6bf60eb390e4f29f6ac913a5801d816165d03d4a293d5cf72a2b3b9604f72659c3d9f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79156c408279afce3856d8a2ab8d2febe8a428ac02fb2648442e7ed8a85413c4d30433d3500f83d5eff01e262878bfefe0d62d70607a7c4f780fe23e6589dbcab405158e36f8ee9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he02874b35476758a413785e004e8563b7c5049a1280305efbaf935e331007b7f386ef258e22189ea2d94ff12b36dbda3ac969e58d9cc6d62646c31a9c97f50c1f9c52379939a7c25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d9b7657190f44fb5d387925289f63899199f516d2083d21e012636d0b6cab036c4f8937aedbda7dd94f0e2cec93f95dcb76ab607c90f799c0481640c68c72529746e22c63c2fa7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ddbcb3c6a3162be1c861ab7b4114e264fb7b8b113f34651f353219cb2597320b7f6109078e88509e5cb50b32de7355b54a7e1c6855da0abb9adbb3acce6f98847a43dd59584297a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha98f3e91a7c0573cc1c00273d17568dbf109d8fa29adf4991c3716dca95a5ce0c20f2c59e32af6d4b4df00651cfbc000118b6ac21370288afc3b4f2f19992add19437424be17bea4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedb6a20a3d74476ae0ab0bd41a60b252ff0aee4b5584b3104046da0bdc719707a96572c994201c84ec31adcf8ead417e7c56ea20d7c9bf1e82cf313196fead29c3b37ae91a8dd5db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h463b95a0801e8c187934ac7c04d54e0709eaf50547e63da1de5a86848d085893a32ca6b67bfe007a69200a455aad6b3c550890bf941ffe1fc49a7f8eb970d7cc3abe9db8005834b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55e9d24c6cf53627149f4acd40dde0c3293e804d889027b4a9671e6fc9fb7b138fe91496c5535af092d90cd6e13d3926410499d69210473649ebe0483cd87a8652bac8016ac2f570;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haec76e3cab7142a0f7270dd6311e1aad268132465f5adfce2fe0336d4b339b2d81a611b5241742bd91b9682e0806e9e63d13881d9f4189dd9bc385c5cd960599fab19bfd0e4518cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ab2592512efe3ac097ee0eb1f52887793918df281a6c3fd0b3a2d3cb47127544c7a1cc6ed5e4eaf7343027cca3d71f4ffac6701dc55fe07cb5ff1151d77740502463773f574f57c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h895ef7b9631d371ebb79c771903da0be668cb9ef84e35de159ce4efc97ea95fe8371146a298d7a3ac1211cb1f41c5ec7add5abfbf8aadbb4fc5c44374f15ca44590d6c0256910444;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40e47191fa0fc8aa175762dc7a2939249544338a3e9261299394cc16d01d17020f16a675bf72d2c34ffe791aa3810d5744a15f17386f26938a97aa320afe1d1f3840a25f42ded8aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3149b814784280e483deeb099661b1dd1beca4a544c638faad40e2b057895372aee13dc9e56ae739120039668add9294aa9a51f2c603d02f50e54acb193d5aff8961366adb1803bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19e6d29a1a258d69945d1ba756ff6fdc33e2be2faceb4b9d8a93088fcd9912574939dfb2697f2e1e4ff01825ce3747d6170ac4cc69e92c603aa5d50f0cd49f74bb9a01657b9fd3ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45b807ce26b7738106b8234d9b7cffcc27531739766e4a92673d26a29bee101d0c406b9664959b968c566e6a0b006ffd3af91ae7d931da7c75eb533c0f25f577547de148c6119131;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3d597c500ecfddf3650885b3328e2ec2dc9bddf3d69cac9f5974d54952b67d715366d41f0c0b661797a6bc0c5810b9bcc9d98d96a0c3825db07f480fb5d6e27932fa5e72a060562;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa90596e81c41eec1de47700caa9ab0db35525da2cd83feb643d5d1d981ab2918db07daa7dcc16995213bf266cf354e5d83e4573f0024d5008d16ac2c6fe9ac24daf55cdaa45a4ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6ca2fd2273eb04a99bf2a7494fb417c9fa2ef6a13e7420188b07ad05e99f59caf16a99b2eb1fa72a81efd40d2618c42d0194c60e2db51835ad68e3360915e57c911c5641cb55f2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d13e08e441548a68c61fda884bcfded37a512ff3e2806405296ba67541e08c9d83294100acb9e8b482e99241375277a9cb0211cc08ab2703a53c25c88ed62f3e1d3bcc4d3b469ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae9dbb581eabebe954c57fb22fc2ab14ed8ab2c24b3e83199534f820e96dd14b6b227022294effc4961d1a756b210deea9a2343dcef30a4ad0d82a066e48ebc6a7a3fe92ddf9f578;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8f030c7993e9a2377539de006ee94a300dcf18ee6a5e2be7e1aa033a2f89d33967bde13ac8f27dffe6c26cebb4ee3bf80931a2c94c28e086bc7e8377b4e49d548186f85ebad481a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e9f9ae3082d71422d7912c08a66f12bff6d92ef257beec99bb4ff8f44389f8ce4be73436e7e59738b6e3d6113598132616aeefda411b13556f1c7f56fa0669881d33a1745fc4f0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a023501932c074a9cd4fdca22c586dde76479f2b18ab94acf9a65f7df2be2ab92304ae9047316789ef9b1d4128629a8b76141260a924c4027ecce989791b0115f556f6a83f8899;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h985e6ca7687f5afe1640a39d3268eefdf6a149f54a2c4ba8ba9eb34cd1c590217888b621be7af8b3047594d97be6a2998dee9fa4b903916472bf4a921de03d748376e5bb45476511;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dd8cd49a275863e9bdd51d261960433c987fceeff3861074cdd099524d35ed986a187d03adf4d6adcd2ad93ee2c79e8667507e2921a1a1c215e127d7b138e76d025668fc1456778;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc09b4d81e5075d2be7e98850493f5067d1a487fa57b58aa82ad926770e2610fc98028c3679eddebd1052dc04fbd68d4ca4e489c455f7520dc0d256b737698743fcfb2eadc8a42755;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4f5652c52ccefb88e7eb439a45e40d6d8038443e1c9a71fc3f99d61a9c5c1f7f5053f5d18ee1389a3d08372a000e38a7caea39858041c78d928702371f446672656de844a21a73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0fef3ee468cd227ee9bbff8048cec3ae45f3c7505beb892a54134e903c54a47e1d82f4b8120961e8b526774f3be28c4fe475eab550040fc9090095ef5b8d2d18d09dcb3c55917f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a506e1ee9726894010460583039663dcf583c290f4b081f3193d4191e7787010ae5c73f4e185d52a1e2728092186537b73b9d491171f87b1d41ef80f2d6def1acffe36c8651275c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8dd7d1e4e3f947967e4a3a3693979b0ada020c59dad4caa357194ba254517ab580f1166151c9df9ce63ca637c1d9bb2b205a14844da6a10fff5a6b50266fe26dacf6e0cfd2221e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8b892728546b1e2307339f07495a2b3014c873065120a6b08b56865f721e98db6b67e6db905311754c3287cb4edfbc663450a3c8db806e4b20a6812bf19574b201b1e500baa6da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22aa52034f6d5b24e1105de17effb95d835356ae24cbe224adf75eed0d65431da42569e4701de234f4150e351a9a9f90400bba3b3bd66ecfc3e76febb240958e7111f8ca1e0cc4e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3a77a1429a5fe58b071c20eed1e688625413e9dc36d672fb3ada5e6158811cccf93b46574c95f7f8cf925f7ddebe7b6ae6d476684e19e6c4f3cd4a762bf0f4e1953e0365e924865;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83101549b91cf146dd2dd6ce9c39fc47ac18dec4edad88fd7fe414ba90ed514e354a10f50634dd8211847843a35d52b416b9d285e32d7009b074549e13fa3165aad897a299abcb38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2937e18415e60fa2bfa6ef4e0e08344b8b7b012a0d5db8094a67ecd2910dd332c158f3c8e1748d3feadb54fb0cb2f90335134747f34eefc220b43934e41cc1f94903e9522334481f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbc18513e13120dcda5aaab01c9d291495b3e7125dd3ddd44b3da67df2ac996ce429d662e04363d9f07889feb6c8c73bf8a0a519112215081bb1197a731e6879ce361db99a39a6d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88f14cc644f8e12a582da437479712527c8819ccd5a867d694718ff96c3648e6330063392d8d69dbf69cd0c13fe31554fb628d6672ddbef1aff051713dbe2a0b8a9a754d7b1adac2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf14e416b50976b8222affd5ca3cf512495576d1145b7476453c22d91fbc79f909d97cff4dc56ee62238daac577a6fcf23ce05ed1afc4d9a1336d12207b3495325badc12e44ce95ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h151200c8450d18820e41fd13ae5876e28b6d15dc0f07857414f2d04c17017712cdb4cdc99f2a805c8078ae5080640ce64d3b26958986485a07f9d9bdb22b183f3e5b1b0fb32d3e21;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habafd3bb2f144e5c3e9d685e2557c8e343cc6ecc2038957f15b964eaba6472a014da528cbefefd09f3b776a9b4c373a92d14b36c46fdb1a9f1928e665f0b780a0589167ecfd58c63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b4aed18c4632cd697c7ea33870523f05d3ca2d1cd988754f296c1804364fd2a3c8a1c8c9b855f964bee22e64f554bb7d6b1264597d1fa6830e62bc3d930d4456c79645615f6da4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34aa6bf63597c41c3351ad467802dc7577c121ceffb11ce868c43339e993424109118e47bd732cd1d47b61b4329319e5cac55b09a5b365d89a7f915c6cd2d5b24d534600ca351b9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he424a56b5df0234a8592992c7c5f3f7691423b2ca7b72697c93c8f7c95ae3c7c83be3a9e1eca5c8dab469e6ddba4b5ecddd167cbe75001597f519c6ea5f8e0331c995321f4ca6166;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbb876c52b78b31e9c1829ccdabe380c18b5b536707237324ac23d05f10b6b23e3e5404e94b1c26bd2dcde1eb4a3be72f2ebae8ff903c8b94e42e2ff2d7f57161414e04b4e9573cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4828c34398056ee8e52c98a4f57bc1ff2f6782c19d4dad3edaa0e45176d06ee474acf4d4c4962e40397d6daac1519c23c5cca96bcc03177846a6bb570e1ec20598718c6a93027c07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44744913f610beee69b9124f74b14466807f84f3647791e13b1c5277cc318b91b33e2831fb9feb6e1800879f51d27003e6dce38b52596c54fbce2a13a6cb2a2bd92eb72deeb6db2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab1507bac9d761b17ff22fd3d1a3896d417e46c709a383c502cff8993582cf41eeaa45265239d358075703233923dad7b33a8d500164d615788d9eaae8ab2c83b4c40d2a91bb47ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f3b78c92e8ddf30c102a21334bc75b2c8dc9f824fd2dc5460bccd0f0e436d9af6fb99268bc74c66ab15f95a9b8e0eb53b269b8801103de5772986d248f5193fa706565e5b310c94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7768db104a679571de4c74c58a8ed1678139bc11e023246570f9e0cd5603d1135eb811565b25da42642fe7f20c6c41394ced13be6cb4dbf4949b5bc6482548d561f97a0d6fc6c55c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3bc8f079c58037d4b196aa6a5ca86a4201f5d22b01190dff1f5a6d17cfcad6ef9d8b63fd4f12489a98e6d0cffa712ba49e5c6302292d556970430e06731b81bebdc30a2afe05a57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h148793cd85f96d4d61c4957255a02da034f230e9ffd3c4adbeec9a1bd3594d4683fb9165322b3d16e43590e2e6936653a64681e2b4e4c04a47345bb3d0ae683d1735b2336e2dad90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dd0b78f24374724a05cf3080825269988cb6db29486a2a46e9a3664c949ee2892565d3870f31cef907c615c907cfc717293735f5a28f6382c02b4fe3ce91cb45d9b5cde2e383bc3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83cf9f93584e0107e393be3ba7687a574bd963660ec922e2a38be51c1ab06f8c21fc87907350ed3242c32c45f76a5d0cfde0e9f24b577769562f1303c7d8ee0c1578e5043a60fc4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6285fe58f9e88ddf3d497840f62173bf1d20b8e030a36619eda248904d694107ba3abec7ee915c90bc38a5d848bf4a371bd502e11d95fc279667bea1a99bdfb9daf70c3a7fbcf24e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ed1a551f177c08c3c0334cdb79679b99d99c9ec518aa04cbca1e14971e805c95eb01d93ca08775e99810bdb0f593319206bc83623f95515d7e4666017df36db34119481d5b8246c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h690b7b03b574de1f50f82d1bb9ecaf626e491b9ffac0010403b574986c6311edbfeda6a10b3404dab8885bc31a2f7013c4d41275f98114489310b25f694fc2883869b720779449c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8487158fff4e258bcf970d86d099bdafcb544502ddf34eeb24b6b8ac94e30605767adbd2de3259a2dfc4860cb0dbee0f38eb31b06047dc764244d3ab85aa2f84f7db5ea5834a582;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc299aa70013103d6e7821d84d6eab1187a9e30cb7a6f098777bbd30280ed609e4c86bd97d8de8b202d32fe21a268c37ac8e315b3775a8f87548811f558f0bbb8d8609db691fcc4e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf14e40e65dd012398f26b7618e1cb22e89e4569037becfa9123061c38a4f82f35bb10014f5bbcf0fea6b96c7cf4b5ee2ef3d6bca177477c29760c35a2ae9838861e926badd67d562;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd145fecb359e43c68a9e01704c2bd6192f9a3c57efc69c9e67639fa22924ff6d447bf3d0d69d9e783683182f4cb85dbcaa3e4a6e5ecec985a2cc9b5daaa4a9a750c23fae7672b06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf577a8fcd23b4ce34ee666a9247ac4f629e60919769fa4085723b33c1df4e8153f685f5753e5a2e9a50335fb05fc2b2b824c9dc8a2b332421d3a0c569650842cfb58c2ee36feb68c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d2e1eedc55a998c202a5b6ed2c42fb97025caaf70da6ca8bea6dc880ced3c42b4f078c3fee2ccd0a53592e007a38ab56c60b4eb1d5d6e9f0cec2cfea4f90687f9326f5c9e18e63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75dddee475a5ce9a06d9489e2f162e91a513590c76defae788bf1285826a66c94789a7b9b411864034d825a08ee50596fa4dad6a98b92b4b8fa0ce28109d613f0f1696a90999c7df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e26e214433bb8dffa1233041ed06afae53831b824a845ced84af1981a0a8af572e9b438988ab23ec84af92b6dee0f9b0a5becfd7dea9229f8478af73adb32cf39092cd1bbbd0721;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ffd9d433bf3393eebe1632524188a9e460fad7e1aa67185d27d79a692916770922c1d909e4cbc7979db4e65c86648ffb6585c0dd08def37b26605f4adccdee72c7dd9d6bcf81f00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h395044b1621168064625cdbab1f2efd940868e2ca24590058a733a510d7a7801571f014087e2c603bacf7a1a08def805cf0bf3a354139b936bad3670e4c3cef08d90d697c716b9d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6acbd90b6106e2eb68f1a3d50aae50de07f243eed29413eeaf512bfe462233f40fa76e3085f67b3da54258ac71026a80ee546da1f8ed3cc2216ebf46282801cb90ed50e44f3558ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2560b41bb4e631d2d94f79f2dcc76f5b01a527f601f51e05efd3014ef86f2517302e3a5043a440ae605d0c404aea408934a23a4f07e9ea6ec6655efc252d7205dd73231b641e8ac4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f56f045fb09f247e74f50f4165cb15e3b03764b52748a2e77cebb78d8e9d60e568c7c21622c60f09213ded6054f9be552fd402db682cf6a7d6091913a7e05cc1e3df9adbe97a6e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e5333c28ae65f0f5b6bf4290eaa7e5c885bc6ea7044a3abb47198ac49896cc55e99553f23b7a23bb4f63d0c1bf0e26c588cd91c6fe3fa4a39110ac04c50ed3613239ae71f8ef675;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c83f86e50232b88f3a1e24fc1fa31e1058bc62602e9d3ad65c6afafab0ec7de687071236315e8e79d6a8de02d09bc95370d549eaccd177f482c43854e37f2a706666dd51d780e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa8219fdd7252054490b514f5be0007766ae09c06ad935d2bb206116414de6dcd35f785e0fa870e49eac81727b39f82e92f6f56fe1cfaca08b51ebc89dbb7d59f88239a552cfccca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc9224e0df5ece0364eeea55e56082f83d11fb52ff7a01e82c942137307eabb89d5c6e3779419c2f1f6967e2a08feecbc810314dcc3950e8ad463c8a3dc0e7a297d1982ad9e8719a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a5844e7fa3ab6f41a29fa57b9b04913c80f73041e7075a4362a0f650608b8f67ae286487f3c49ac535b308b10bf391edc63dfe9661824dd9f7d37a65bd04e23db3fb593b6216924;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb18ec9b8d4da82384318349f6e67528022c58bfe720384ebd7e2c1e35e593fbc253ff16010b2cd00db6cb61679f62fe84ae4091836fe89280a6d74decfa91190cda4c539fdaa189e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1776eafb55a3d722549982af625f28916bf45dff12b245088044b336281bd85fa0038d17aa27b70f5a334a9c733ce8061a407f805c5400bbf37d3c4c900a0c508e670aa48efb591c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4392f5b100f99ba1d5e160f3022d2e4284f4631b2706413673c8c4e9c63eb421ab23de7a3a15aad5572b351f9c3b879ffd3df997afaa42eef2d0fbe27c95f82cd783e417f249c83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3faa84adfb687647be7dc380ace16e02aab26440dbaaa1f05dd01fd30177b57927d4802f9abf1495257135a45aee1bf3d78bb3474e66c89ff4feeaaaf12ac2569050863d50d496d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0083dd95bf77a775387e556b97387e5205fe12dda0c17cb8817c6420f81846f8ac42f9fa49c9088d141c719b603e3193b1ab8c27b19e33044c48b304a8945ae740936b9cdef2c2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30334bfc7ee56630f02e809e551618f6c1305f086b21ab00c855677a7b14fe8988b04f80e63bf4cf9ed34d459643e4127b5849bd81d301ffeae35899486d2f37264b890703579d69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h648c71002258e3d5448cccb737b398a8e3fd6791bb52c7c452c341626386ae3cb3da506d49f38d3868770bd88ee1d0b005790aae1ec3bd8557a1f5d424db808b82a42b440930795;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8839b8e012d13dc48d916c671806d36bfa4c7fc5dd30a2515aa1920d2b088ea154a96f5ca94c26848a3b6ab3376c84b6cf23296718b7ddbe1f37c4ca59a0df5e1174a14e7528ae38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc7556da426915dc21a91d10b27f8728c015ae919561970ea11b8c9077d1005761050fd8b9e42f9567cfbfd684343ad8cce9e7458f24df58fd621d7ddcfd808c76de61a2610a062;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ad6cbc241094ce69f3fe92966c41477907ac484c70d1b3a27788a2906b433a281660382ddd82b026e39209ff53962efec6e0f8a7df60843af711a756afa40e9751f57e880065921;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37efa83f012117a653b2f922290744a0f4bdd505fe1066d78c296314c6f4577ad48ae20b0796970a43e23f09052843f5297586d39a48eb898f8c60fbb1fa19643940b4df928f0e69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc246bd2db1b3725b7df1ed2e61e9f739d89ed3ccdf583ae44ffdbc0e4894aade4e026aee8e282b228895358ef9ee1984460121b1a605391d8ecb81930e89c6a14a5ca618594c65c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a09f7547f4a011c95cd8889a9dc3daa59cc2309bf34d4187cd464bb6dde547ac0662d1907987addfe8f6805ec801031c0c907de9637f2c327ea367e69dd77359e9f994ef517609e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c2d5c38ad5b5914de9309b2906a60ae72f5888a4c740a6f12bf432767249aa9e26a86eed5b32730bf71953697bbad5cfabad1bff4fac434030521a2398ba61371d151c48d9deffc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h208a1396808a4bbf0343b98fd6bee0ec76abb19793af04e52f465f170f205224091d6663b133ab2464ac55677f38a51e9acd1fbd8a49b49809f4d939d37ee49b60ddb681e12a2465;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h817dabcaef5b16ac77f660e8d62b126c442b2d85740207f2ac4fbe0e516a01a3a2cb6c5a7de7b0e472c34465c0ef01558085cf94c847d742577a6bd8b80e23511c5fa91ab0d60d07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb03c0c110d18d7a98eb2345cdc8893a775c4244f7f993c3e44a507f9fe4f3d4d3e51f32419b874d21b5127a0f6c664e0e3c984b3316c167823e0cd613ea3213a332ebc5991b33c71;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bf5ae75f2e834c2e2e3c5f4e88321febfe258a4e33b0d851492c18c70902f2053ece87630f871d85ad8fb5e2d6df468cd22859f3a3834ef57acf298b8df3aa56938e0a22cd2fd76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb44ccd1a37b42e4d1f9c9341c616f60cf6eb27b4d472e7cde2fe1a5c96c1392aef586015ee1a5bc4d260ae2076ef0ef9741516e5483626619f9e0c39579611de50e0c0a69509fb41;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e45a133081ba72ce18b6e100f5af8e956fdf1f157b6a64f3c92d98279463ee2398a3cd74dd4f77296501ea19dc50323fca4a386e920d04ad0dce7e219246ddc91da44e5e95724b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h922d2d381d0536547d8f36d1181190a7da21cb9bed4a60eba5e7258402b998e8e4345fd126057947624458a239199b6229ae24ddc03fa719afa895cc800e1f590934b655f4657b49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64338fa9a1b8a774e22c0d09e9e07e92f1449df0511464db39b6db1d8e7b97c109d5ac126b6f6c6413a047402bc589e75d84d1017b18db37b476d242aba4ff9020f17cd55c3fa483;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f56e88aa3f1e7acb3bfe361fdb91de208dcc2ae1c32f005ef48640664a884af8ed8a42e2740ff400db95dcde0b9a31ae7b5279dd5924e5d4ed442d9c5b6e088db09dd7cbc5fd5c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3814fd83e754a08850ce4ee32e52fbd9c8889c8875fd50a4dac66d857264680cc6348386a21b56c2ac8441e392af4cbe1d64797ecd53659fbf3e69e5b2cfe429abdee7ba98945eba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22e0bdbc1dd09b5fb39dab57244d7c7f5711c8326d2ef223ab0666bdab8372254b11408bbca7eb80d10099b9477c760f5405c092aa30c956570bc7702982715f744146aa1a914cd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21da2d279e2c0913f7f0e9e703dc5cd4376c78f5aeb6fd92535c6471a795ad8a52316b02cbe43237624e83532c1bbfc53488303db02cf4dae2b55fb6aad2b4ecbf818749e17c69ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b91380e5bf188527d3928626237036fe03642c7ffe2067bd545ac219d24c4101468cc99747bfdeea4fb06847b19b1e7a68e01cf6f63e38a4cf276089d3e4dd7c2076d90d2de51d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h883f09d7266ffb63ba0858e2f5bf14397640c1bbc7b5885722854e2ef4225426f16a7d83648120231e1c5529c9d3d1d5b3c42e64b2d8adfe555b9ae2e94a90926a6f15ed54f8f2d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd198d9a8c4d24da44d3962d6ec0b74f12e577fb60413750203fe62e172a312454d1c1fda668ba9cd78e3fce00b9aa3cf1be57c34b631f4fc66993822ad758e56a5741c6928f4226;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4435080c947fd46df7d61f3634aad09eb41e4de41ac4a8f02e5c404e9f4b38ac6a2613537f7e7d35fd5e91df66d200a2b9cd4eb26b630e5c290af16bfe71608fb3c36ce6c03a9b2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82041c29f435c43f54f78852de065e0f3ad9c99555642387ab971ae6a9ff24c96435de77dfae4bdfbc4e0a00a5df2f9ce2b85951b8b85aabafc1686660dafafc3666a38cdb2d0879;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h677a80064ddc19fe2be2dcab658d72ebd21b38259a42d8fe3665f7705a843bfa8064845074b980bd68ac5b8cfb38d6d1e3d7856c28b4003fe23cb9f9556e967d25faaad3b9b0e964;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d5779386e4fa4ab9040c3053ab24e24c417c204b1d17881f1fcfd5dc45e49081753d33db2d499de3b0a32b3906b6b3133d98a2910bc80fb93f056c43ce72f66c498b52d37da04e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1a5bb43d727552f1440f9df33b7680b7ab1723bee65c1f96e99a651b4bb76fda5fa6aa3c7f4e5580a48b59866f2d1b4a6410f683a7e1e328ed95a6bcc535ec7d96083a48f1dd952;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0711ea24a4428110e93b56760c3c27305c4629f2b3aa0d4e1ecc33a76ec63a2ceac0cbbb7f257d2362339ef1917bd517997961031a18ebf94e059957bd9a794ea8f6bc18c889309;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c671ce0fb1802ce1ebcaef0e341607760033efaabc90540134e4c79ffd10d24bdf2e3fbad4ae164e81a503109a7d949a28096db0d1286c631ec871887fc1167378f11bdc5322ef4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e90c648000b299e67b9fd39627a773ca18eead240c1f8ca91e3d735b677a296351467f80389493e14974e1942bceafab1e610ee93cd21978eaf323bb94b9deefde0ca4e0402aa77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he65a9abf433793a61df15736a289839a02a17214742836f4f21567a4edea07a54174fffedd85a5ab7eefdf824cc6454f67227ee2c89dbf912a61b81dbdae978eb12c6c692585fe0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5ea960e7c73f665d0be205ca24ce4fa16f74cba757a4272b38e0febd63a9191de6f9567fe0ad6d5de3f944b516e935ee4365fd00801af5df8784f64f638f3066579af249187ad76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f1af832d260b60725bd96d06c7d7ca19061e156c08f66453845e4bd75e5ab2da69efaa414716456957af1f400ebccb1770b09a969d6cd5b7454f561440c811c35d7822fa528508;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd98e9eca1d8b0244348d397280ba9991750417370bf74202a34661fd0926b96059a77731e57b53523eb1a93e10c6b4721c7180d21a9eb6bd33e34f94715032eca99b56fbd04a04fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcab97991e268f8bb1d91c2e70544a0b38544a99de9480ad4bc523b020f25b0813a50330d1a4bd12f44c2ede572486dd3731e43ad672c248a47c9690d0f7a2dda54ae54cd7d9ba1ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63de1c9b02a0260264cd4f438621b11cfdd5072654ba6e659aa42d95825d2048e483de623e760ba5255a9e26cf9c1652f7acacae88020cc275655246885e50186de9e3248a1153d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd11160fcd385b285beac0ffc3d6458abf68fabcf000695673b845bc2ddee492e3f16ae6ec04805681fc123b1ccf73161cdf1a5f2fe4b6bfd6f0b41b56776d55648a28cb97f4cd3a9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbf2dd21eebf918671a9a16a4ed21e5099cdd3b4353a99c24ea255c7c1860733f3bb5e4678a68a017ae5b859b8a345bea73466abb4e0f513e1bb1ee177f6df45f3bd7c8155056ec9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b78e014692d8201f919ad6b81b4231da1a25f012ba595ebdaba6fba9a5bdb7bd0b09573bf8155983caab617cd6d25801b29b45d071c607aea4ee80a94183168cf0aae29bdbf1fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaf60fcf8582558260aa3eb098f8fe2b04ed3f547f03bfc0a1b21b64689101a6a1b86af21ebc63ea4bff916598d0a7947693c8b940fc0b58c1685d8d061756d9aa462ca769b111ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4992a28a867fc0b6bdffd69dedd99c7fe95f6d8be00372652f10197f7547c2969ab77bdec0f422d969dfa9109f081b169dfe6f1a86186a00a756949341a4e27a95d2196c503174b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfedcc8c93af4aa345b7da1fb343690ef4dfa5b416bb6cc7bffc90b8c90f940ec34e5c8f6b2b602d89fec4681ea69752c0300149e20254e21dc16e4eb8a66e9d289421c281664851c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6471e8af27f16ba1afafe820094055db9d767f9d7d5bbd4f895a96f0b755d741b9889c6bf72d5e516fe0d52e63933e53da75145eedcb997cd70224bb46451261e06755356f09751;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95d902e238cf941042b7711168315928ee6a6a14d5c61dfaec75cafa3360c1d229b34b11bc11f6e8e73b50de8ad7a25401c894b458e04c4b6918bf31d405366165b361f94c62072e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f0c2fd0ddc3b4657a188f71b2c1d992c07ecc02e900768c70e7e9289ec2de2f504d1698334d82c6efb9ba49543119271325cbc6095aae954165d349b718712a9a8ec930d6ebc39b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h791c9f9e6946ef23d2449665b90682135ab10e1f76d9639bf3d750b5cb470192a78f4be0cbdedc24b3b769caf8668958c16862a98f6119d60c20365e9d7a742a7d172e595af3e300;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h467d9f164c1abb14f19cd8a0bb690121cdac0c63509394ce70b757175bcd4a6f8e91f8f3054145369ce9c1c550b553381070ef0c28a8b376486ac2793cc4d004c3779a7d232c2336;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e77906aaab7631283ee3cae558a2d218a427390560077556370d77b01176df72429744a56b8b20222283abd00cbafc80d0f23047eef7cfdc227e5a2b2a3257b5403ed208b47f0b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he21a704b4305501e31d448c0c7a9f40d46ae1e8f6394682b0558ac0129200a38cdb92263d21b3ba12e4661441a4be7b3684f26b4965fcc9087cb962af38468cccce878eacf090d05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5c9e07e981f29025e742f89ba4103d3b37a780cd6d095f4224fc7b39e355c72e03b981ca7027509d74964d8b76d36c7a3f5454b6c235e20d9ab51ce5a69fb87441909ed2bcb7c9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d9ea546e2b758a115be6516816360682264d933196ce0dc7cc71b9d6601d333957163af9a3f16fdeb9e78e1f62fdbdb81013a404cf86064c4b7dbfdaeefff1b190b3310f000260c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5c04a764652692fc807cd28c6fcc31b9bd1ec60aeea2aba956602e1fd601db424513ce8a9add29ad9e5b5b91a021c9cd83b9abd5e948be9f18ecfcc76f0b8c8f05ebe91d509f7a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5352ad03e4c8543674ce37b8e299fd027a0c6277888ee1f0df75bd38bfe3d4e3ac3b6b0f93c667793f0f54e658b796f894de5207cf7c5b0eb924e6d993f1220245982ee18470b84a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hada1f224906a8e1dd773a82b91b50315582759a55a5e1db74da23601f2f5f469183706b556e895680296d5f4cae83fc02863a12652324c0b2bdb63e4c4e506fcf002c495d8598f18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d4a8678368412660537eac0ebd3e724299e0ba3b5e1787fc90fff0068ae6743431c091d8f472be66c364dec39a8b7535cdf8058b28715acd113b281f039a0b8a698935078f9723;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e8a07f23f9e1303209bcb03b7a3a5296e20640a43ccd7521998c42113a521dd2ef64acbbaed4f7b01c3dcacaf299df053ba18b06886000344bcf3171999696eeedd4931ebe92f2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb322e533c9f21521a8eaf422f0554771b754c89c16106783888db1ae5daf1ab73d7f55bd445a9975095a16e6c745e26f883c3c2f0c84dddda9c883be0c4c62c9d7dc237d89860356;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39f1bd6d4c5acfeaddf5cb1c45e3cebf5988cb158813ade3605a0cf8a8a8cb5a1219c91a0ead0c65830e9c0ae9926893ccda57ebdfa776a729a848cb701175bb9b951b4fd869baf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8612735f778bafe909123501d6601677ed65c9ec3d1b6648e8070d2a5c7e97eb7f75398b4df9c0e5cabf6ce52c7c221e5ff2b3ee36f4df2db3df0a0a3bfbef3f5a8f5d0913cb990;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf99df849fb86e49124ce377fac3eed861e32944a33b8db964cfc49278076b6b078f7080773bd8025920ca1cc82e64bcb7975c15ec528aa065124ecbdb3686ea27c06e0ffd46589cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e8215507325e5588903916e54c862b6a14aeac25da28e6fba9c46e914d69b5d915dd30ef376cb594edecc1112439e6a15e36432da4d47f049fc5cd9725fa90e2edce52392b81358;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc664ef73ca4b9b040f9383141b44d49f1fb87a9dd452bbfe1c81f4034ee73acd650a0c18bf3497610391f18fcdbada48fde054b9ae3b5827d75fe2885a49ed543ee3a4263b8ff91c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c658dafc4e03e16fc1bed2bc1d5de8cc297bf03f4c0c493d49061323a9dcca83afae790496b9172c0c29210ab88febf7af9a503a27d7c4eebadd39cb6ad5fc3a66532147e86a7d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1670178991b0ee2518076a1f8dcf0893ccdc54298f412703414c5295ce72f65a199de81099757a25a85e4e19ebc01160aa1fe42492a8292818282390816c8e3ebc23edea17a4fba0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae454ba3cf252fe6cde589adaa922068f200e872ef5d257e6d975bd1c01f1e9914934e7d5942f7a55ad90208dc8f98720128b94408874310eca890755244d2420879878006ddb7a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ae4f3fc32932a9bc8bb09f71f15a680a9170ca371cd3a1ac0f01d17c771d0f77d3d1239b5c3e7e4faf154548e90bad3ffb4681075ab2c3a44bcaa4974a17d0c4dacc680275db623;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c7eb618c7b64129f8ea98c28743761d109e85c0d445b25982f2ba3ac184ea590c4b4727f2d6cfbbaebdf191aca0171484aaa6fb705d0134ebc3a5e83e87dde40786b738d508e12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e2b5368df09c794e5bb37572d90dc63ea0e9602b124b7f8e76fae3bca64f2928dbe14f260dd98044ea90496d16bf047754b20fdda44b63dda587873bbe63128494be7867f625ed2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70599d7b0771aaf9bfbbf9685e3d5eb8205035f7e9a82220eb11397811f5549bd15e3340f4955000133ec10030ab6e6d2123a090089ed4d5d0018d5bebd72f393b2f2e36399baf64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf40979474b5214d44e1fa3b12d2ff451127e72d3b6d406bad59cf5d7c807efd07b766ef9ffdf2f801958a9ef96bfc0fd6176c124f9bc8797a443998d12770d1d9cf595b3618141cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbc5d8749a76ecfc5a9a629474dab04f5028fc8d7f5279c45d621ab8bc5e997f72a4a0dfe84325e40dedddf9200d3e2edc8100a738ad7ec08bd28c9a95b5b55d689490de0a449eb5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69238d2ddc0260693e2df4862df3b5f3c67421d6817b81be5780e82636ab95b11a1b774b245d76e654c467f0ed1d9b3f8d4b4d26d66aca393ecde175ef4318ab92511631409ee44d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heacfe3ea4e08086f9edd1fa4bdc71e4090d586f5f914f382885bd6d5a50ba76362ab38c6a3d84153977c3955fd0365f5499f42bb39be24f538313feeb374b7d836c432c116d2069f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8275647025bc364b4d8393948cdd5366cc8dbb7d577bb2382dbe2237e6c957d55fe991cd683a0d5d071c6abbaf72cc2ccaf1d7a40060c3883a03d8a846971ac7ee7a1747b160c1e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd55a8192ab105e68ef766f46cf1f70a53a5fa81f9750549b542c4eb93ada63a2db2ac448740c705e4d1e75f0932e526c3c67999c876d5e3c310ee4f6bbc03208b46830a0ee73c576;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6d5e26cabd408f6990578530fd06ea93930d3738aa4e3374db4cd5bfda517d4878306e297278f9c2ea809dff695233ea5db0095f116390b7ee1f7217f160a5ee2e10d8636b0d7df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76f094b2c9640b39d718c95231d2a321849942352d79c9a07b3851863a46a60b6eb6671c650ca7a8f1bf68363aa9237040219529a095be80017c9791e5488a67c15e28a5a95350bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b750c707c50b33366095ada2c411bf25faf9bdda02cd0995a649ec08c80d7888c320232b4574f13a369d6dcf5448de3211c19aeeb97237ca5b65fd670ed1143c4e87c94d999fd1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbdcd6edf14f46a08bf530dc6d5a334a694c42d3905ce909fb3c5365c0001f194337026377d4440354b9d36fc1cece913968768fcf9eb06196a002721931df826e2771cf6839cb1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dbbae7945553542f23cf8eaa4285070f7a04e49b66d8f9548e89349ba408843a0c387a406b57eb71ec804636c02eb85747ef46461b6189f09f0de68e199964f01d72ea83842195f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h339fc004aec6b41a6e518d9a7c8b0133b01645b257d59836958302f3cacc781610f9e1cf6fe531d88ae132bf394c975d134b4ad1afce961bc51f974bf49c269328503c912246d08b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e7da93dac704e652b48cb44a82a284adf6b3c74d97f1c724a74fe2c5bc34e1c3cd8638f56db27a9467caa41e6b0f59481fb64ad28550c0ea96cfeb0509577626191cc61c3896b49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b2909cff99e6b6bdf5e8bc816970f81f4cf2b90068d0b2b8cf2fe4822618e8b8f04cd6ae8bf8f729b26a1b56424dca3e3d3736544604beb87d38476f17ffe3b234f5b8a364297d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b156bca51abd1e7f1f49e63e703d5c10c4ed5c3bb2d4044f2c7f70fd3e389ef474813e4951792498502912dea11cf8f37a980705b930243bc3604cf60b268af80e504b204929f3c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h858b6fbbd646a46559bb044fb4d17d53f2d36a7d54114f7b4ec63eb88d92c5793bb1052b549c95172302f3d7516b85bdfbf16a15c72e95d90d3d014a5b1dc6551167cc94cd285e18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51c19c515c477fff204e35f279b6114fd0e435cd7c4d55999b2a127fb2cb7a4c1b5bb4b15d7012102b4e77aa7ac65222e092e64642d195535b66f025ab6a4eb74e34445b37c0a725;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70b41871c225d4c533e24a5a704c784011d18b0c4aaee93347fc8568faac406da7982fffef69760fbd29fbe9a8d8bf9a6da87d1d117fca970995181fad709057f1b848441bf98896;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1a5b4aacc8ccc60795e60ae4b824eee1a3c7f251d00e84a71e80d7f09b1fb7877ae6fabf4dc7036e76e1c99974add18d1f044d4b15381ef28034b81b1b5465d71aeade5fcbf3ebb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82ba0d32f946c9214b04bc5256170d62aaca4e19306308ac9cb7e56bc0c8c20b5f132a20b790328950d70f7a72fd24c7d6cf028e2bbbf7f012d2d5fc5b2ffd96be79965375d3ea70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe0cd6e604d8e61303413196a1c62633bf2eed012cf728bd12e6b0862802c2d25b6bd41625dafceeac52a74475baf2a24910126e18d39746fcc44d5be6231e85189ed4f83ab01c29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5af3f79cf11bdad25ea43af3997ab0f6637fb3e454e22f055948c4a3f17dddcdcc51238bd9c8b28dae4357488862aeda67e5be6208bab2efe27d874602ef1fceb10942c57a7ce63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd204d0772f987ea6dca815a52a36dfeb9fb80b6c8c0815e881db9261ec9ca76f5a810074eae4146e8dd3a36800b649a678cfa3d7ddab88b8d8aa948839342075c3af6a520a194aa7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14863a465532cb4dfa7ba7494adeb9f581ddefd472b544246ea9314bc0753d1fa28f50db20922157fd6fbffccc174505c89e74b34c1c6eb52c725ce70c96f82197585f761767230e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7d1d46f287c1b21b9ab61e7adcd02c1bb3a7ba11352ac977fb7bc2e73198e4031143594879f59b7d3cb2e41c0b3cf37ead0421f3569201dabef70a6029bc117940631163a3160e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0584e33d62f40c4fc0c4609cdd7ddc7ada2c8fe16e1e81be9a9e39ccd7b7703683e6266d0d761f3f5d1ad3517991c7be0599f88ec9de033643c5cd7e53a71075d32d0f691e8085;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he20659b7fd959791f23d40a0f601ea1cd413f1de9482af451a54253f5a5a27926cd7fcb85069fcf135d93fbf7f0ee0c336e0946c3e5bbd2de78a9731965e441b092b3f38c6eee2b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7c889da7c216f7a036144e8902f50feccb6a07131af229030b3f06ae3b8de31a3a9343390c40e5330078da725fdcf6bbd955787783988017ecf008b8d59a851b9682aa2ae7e0357;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13c4fc05a48c34a6336180c84a847e96e087ff750629d04d4380332d4f5d7485fb26f900da962ae891f4e8babd1631821929389d60d6a0fa58c036597af6f877686da7a1694e63da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he33d192af8c56850873ab17193520b0f4bcc8e3a0d83a745b872d8135df664c743654b0336f3d0808d54399cfa2359e63e50d348a4e3150b6922794402bf88480ec9193eae16609c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ccbea83c1d5bdcfbb00e83bb31fef178af521b682a3d8d895a7a6f7fe98d366979f9592d3400d4e306827776d857e18f8a3c5462a69a0111ef10035023022c8ec7fc4b1387f21e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba746ecfa7a840d47bd9caed1d9655a3346e64d91e9f310f6f9e4e46725abbb74b46c20294f81d86a6d7fe0cf6d257a6c2c81fe4efa9d60a3daa0ec4eebb36d2b779dc65b4570f9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7a752033e262b876927d5e975ad57fc2ae80d7117d700a6d1dc144513e5ae37610823795baef9a3dcd3abdb00743ae33c066f487276c8400d8c46ae4cd53a090c3ca9b7ae867f94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84357981ec898e952cbc2f4f3ed95d9359907596bd8545e697e345925e1c3c404990ebdba550925e383d74493bdd8d0c8e2546e3572b255c847f4b1bd9d6dca1a9773021446d6f1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h586ce06d4476f3e8c04cc5c93ba3349d5960023a4403374e90d17a9da68c92d23d8fb884a22e92ce7929a44f5aa1807d975046fc036c9c3eba2990260a2102b35cb15261eec20d5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6111ef050a141660bd8d19cc129879c75285a19398d519040809a91b5bd53c1e7c4a956a9ac8f091cccd4499b9b37396c9a09c66bab85d115846c36f72946140bfafde3dabe9c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd3c60ae1156800eeffd2e7836ce2ae59168f61337d9cb7471cabd3d6796a4a0292485bcabaf9847d80af5b5352d0b499ab404a3776cb398eb47fb82496c16b543bd55bba8e626df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he17e86582d43c01ede976a66dc6ea8c43f7c456247bc74940288da79845e6f14833f072f4e1a0efc0556f74416f9f95c6f705fd11764b1e68988775c4a7a18efa997e77a7cd2fe79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccf41c5d94e760c2eb3ba204ef5f515c16e95118d29e17f353ccad9147e9eaede5155fd35be40a9df40e4cc4a84616d0c0ff161402383350560e1433ae02e21f531d6c6f5a97be8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had7ecc489dee085dabb1ce97a1f35ddccbccd5418fa2945805ff8705cd6f260da1aae173ad84375cbbfaac234bf2ddc2e02994b82812f4baa3b30b66219ce4b32ba0fb954a8d4c6b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43944f90e5d669bd38172839bfe552b5637dc8fa4d3c7e24a6e23c6cf9362d4c07439ddf0ee3ce3f45b602eedd2820c84b964338cb1b502499ade2f112b2f02d28be51a81137059c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ca60fafee558f37d31ba7126fb9ab5e7d1664033b1c1b53540d44cb615ebf63ad20d8405eb91939a3b06600660c36f431d96e10cb281f1af0e77ab8eb2f7cc15ab25966af198cf0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h338a17968370822bad5a8c18fe2b7d6be5d4edf330ac6295c975fb8ed73f321a97ce013b353111af3a1085dd8ef7a01f7c03c56195e33fc3414bdd186958468bfde37272d617421;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fa0780d433bebe3c41e18e3c17a054102155f68582410d682f2780eea8f8d6fffefd8829abaff0984855ff87fa4e2ede545eb0c04e2f8f2d6903b7717b557d859a83d7a5c716835;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78c6ae4dd43f718a1c9fb79764ed9c915b9b167c1ce1d5b12df8dfed19274a3de7c521ac7f8ebeb9262ad4006b6667d5adf072ecc6493908b552ca2abe45f5a43f6ee79936915e33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5860d8eac7f3812f1bdda14872a907b1e6e9e13c4c0dd7f796673502d1cba0009b225be103d1d7ca15f79838274c459e7a7dbfbf2b3151866a33a8cb4ab188514710eccec06d7a99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff01ad5f90e94b6a20f35388082d5fa34d05b7806d5418f02964aa5f3ff0b1c5e4bf2132eedf49c1cdd49ca8d3c8e7d23f226d48f93bc4bc53f193e72e9065600472306d6f7cacba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72a87a959e00dffbffa3399d3ceb21ee96a91e17fb29104eec70c1cd8fd8a3efba0f4258493e7e1360798f280687fa7c5225939c04adebf81589d96f59d3d3b7db5825920a554fd9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89b6aab4ecdadc70575f9e225960db577129364a3fb262094a18cb1194eb3838c0dfa8bccaa5031082342b570b16795f9a9a85efc2c3620431368562108cb96a9cd9553c495a626c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1a23f2feff75a25ea5aa44c57c6fedb8ec30733a1e4c9f43582dafcad006153aea03a36826d6ab00e504da51fdd7b7bb7073112570148c09b817c938e10aeef4a430b7869121829;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa9dbf3eee1df77ff2405ef765322771faf854f9c526d2509e3c654d5a3f016c6d24b44e61a0151c78bcfa0ea1a9f55d6a620675e9e9595475ae77f7bceebb4599fd68a29254aafc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95a1e6b616bdd7b59f68e790b71069864c14774f8c8f8fef626904de924d3daa0f6dde87ccad4d6beff1f836a3bfceb5ed8eef8f512da8ce99295c05c5e5e78e6e6e83852db06dde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h932191280160b7f679a27ca84c1ea1e74701118adcbdac0bfa5171c8f194bd076abfa9bfc9d57a56c0f848e4c8b8ba73a53983b6443b2d3944d6f2d18334b350f3506551b821c59b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he167f795b43d2faec04a154bb171e5ff7a1c865a5adfa1f13f4583a4695acf92bf7317891088ea5627eab25c7bea80898b1a80bb5bd086991b912ba16e2b69275a84ad48db4badc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfed0c23288714aa85860dfe5a6269e655cd9ff192a5f6b681e8177ad1cf96682dca331bfe36537c9ace6622ed663a3999812a89c1b81283a51569b0ffd17bb794083d08ded89ffa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ba8575c0fa380e887706998378270423c4adf44e42a97005e78e3af447beb3e9f65293b2d55f54281669ef2bf31c1be5fa3e257bd4c3db1dba4f87917437a755e649a291b211e9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8ae8a9ee64a7c97e811865df18586dd5eb309fa72a26ee2fe742c025253fa4482fd846d25c318995f4b6a22216011a778c8a3bc9a1e0cd0b1afa45e31d4a6687874b7112431c0e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4071c322615963a99398ccf1c36236e0a74c4a3d0345763962701641890718b0eac4b3d00955d0a60417e163928f0ea8a0ce0a594b5545f9d5f8fe65425f3638427bf1a837d39f38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h244bd5ea1c283db96465c0a6a22b16d048424019be2815d336a4bad14a30dc188cef255b48b72de02a297e3e8c14eaad43ccf665bc5bd8a43fca3210982776596ea73787b4a8e7eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79fffbc5eb0b21b03ec59117f486a94a6ebc80f6d65fb52e8a590bce87a4423a5fc503676ca76d092f449a4f467616b2902780f4bdb82a108aebfbd63be29db5a35527d68576c60c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h790c389ffd4d0bc0aef9f82b130c36e2cc0a760a38bb437626ceffe13da7050cf7ce171f3ae81265552623c22de23c2710a3625580f1581baa1b365f4947322d467346ddda03c392;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55322bb3bef08997210fa6967729378222eb8e368a35ee61cd04ed4c80117fa1e20f00d610209ecee7529b5f0964881f62f2dbee31275b1aeee99154128aacfd32450cda5fee2b32;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea6532bab066908e418a85d7cf494de767b6363d21dbd47cb025d778bcc1336f6ad0a391b4a31668df8a879ad267a2bbe6a2e5088a70c1ff363fba48ed19002a8da345a9130ce656;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h951de25003e3308c9ee76021f003fd1ece549432d0ee5ff34c7a6a2712f381fd15fade43293d0661f6a85804dfca4635fae55360f905b9e139ebb3379a0e042b284dc95de0ac167b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ffc72fc2666c109bb666d3083a58020e1155680c3f5358e201c14128c842bb7194ac7dae333600b0c050c3238186dc67bdfb1d9ce7556bb3d696626af927bb8d02ba8c52f758b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f02d8668c4d33e680fa717be232ee6e132941a89a4f1026ade6d4086c26792dd9621f31f5493ee2b816a1f67ab6d14e52a44e27b03acbadace9bee6b8ce6dd30a4ee636539af65a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf92b1f442789e04d39f4e600c91730f79a8e04702b9813b1700bfbe74196d752c788dfe914bc447383cbfeeb63584038a5290a70afcca77421f4dd642981cb323a520021dfaa8ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha08a7c3ecf7162cff011f111046715756e0ff0fb8dae2594639d2e7b529041011f3def0a903001e0f33e433ed92a5f907013c52980a0d98ddd998ccdb6af6556b207f9662e8bdfe6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f6e84de23627cf3f7744c9925d1d635520ef970d10b679c19e3203ac44436237424a9e768fcc5dada8a56314f6f45c2b7f3309677dbd6ba06df400f0bc6dcf3b2013e202759d6b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe68c6bbcd232cc9cbe252e5a5ba6c0444c2cdcdef9dafb62ed3dd43fb33b865e5a168b1717ce3e1383557604741714533e93fbefa2d5ef3219c8d5d72196a120dbe66017bf61c8d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6176a5f5c1a643d5c1f5d79dc133d6ecad5067df37ab724192a84880838add118ed9dfd2ad52494c6332718f6e5e486092659ab1956792e48579338f00f1cf3d105336607ee9fa9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3ba0262599a742459465d07fff1271f938a98aca039a6fe01cab5eae3ee65fda74761c0cbecd201d7e9bcdfeb985c8d63741c05e77377a3a8a786469c26801ba17eb5ac444dfff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3bfe2198a2b079954c52ed00a5ed68f3c30da30c8b2d3a8236f5669e630d8daa3ccdde1f2d38824b1c6230987fe1fd2c80553e484787d9a3f3caaa70ed5317b33bb56a7a54ac389;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf536e69feb4f5da7229c1c38e16ee9d90a334145686c3af5702a1154dc25beb4d66d4f05b4899207a62e1d060f6af9af826307913041aeaedf11d3ce619bbbb26a833132d4edb8cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb46584592061c105e9b9b79eef19358cb6dcb7e55b723a9eca2bc684fb0905f3ecd830d32cec4531623c3c76bab0f67d1c6a6436815ee5dc6a4d4ddcae40503c27ac21588f3c71c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd35e9afc19e051fe350fc2e84d6347077387720f408ca93ebd2e701a224bfaa8344d2a8259c3789bd7477d69ad90b34c10dc13bf6aa9268147e9a2ff5ab29b881e1cbc69f2f8017f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2db8248b4a55652f91e3b964678f29ec8bc3284b10dd57230f660a29cd50fee9099fc6f30376693035c8c4c1bb61f0005bd9e2e9ff5050763dd16d805b826cf2d56111e2d8f664bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc87930326c563a2607e332830f263b09872012333659225534c8c945b66ac72f3a5bf3b3990dc93d8d73845a1869b6b8735e6df1f167d8fb00b6b039810ed036996739c401f0ad4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cf54a70716917142ef4693832755640a38f2e974e3b2b9216f33231732b41f9cac95949187ca3f78128d1293d820836fcf26c2311205fa2b0bf0a5d47c8a15b84816294f5431ce2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h719f7bb2ec03f2e58e40333f37fd1c84cc1734585a6c2806bd5b5187b2d2d6ea14bf384f1107b37d29efe105268ef3fb395543eabb9e63b10203b2b5266206f714fe6ab72b19cfb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ce206e4e9da462daba7180aca398d348260fb85a8b7001e02360ab5088c973d94abf2e013ea28f1ca912904441c7597838335b2a2041fca3b7ae61b3dfa99117939f4c36b6980e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecb30a8d6a187bc6073a51b41b6c53e8df08e34d0fe1fd03ab575a6dcf677d99a8bbd091dc6beb8ea232aca35926fe57f4b035d5b32119e32824c70b5e99e6c77e4950c99217e200;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac63d2f36e0b5119c57f3c404111903a45f36160c3fc5fd1bf2d6226f43545f337ebd9795a5ff42521a166cf8b1940d0c7bedad9a6f6c3bd8eeef68f1aa1ef31320fb0c86bde5ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc487fcaae59aa96af6f7d16ead0149f1d62dcc9acbe2e720eeefcd609316ed435484bb4df9e85f8a420a6ba798a386d9196ff5c519045ee606e4d67ae94de97b36d7c3df07545a86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2e4d2cdb28437ec69ab3f3c62e36137fa7b28ce0a14081ea7401fbe71d82e9de1be059a6ac99151f53e7f3329caa60d5b50e35bd056a4795ebef5d2a89ebd2ecfe5dc11268ed531;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a2a5b7bef31dc6ef81f8dfdc8c44eb1925e5e586c1adacf317e453c5753263237be80b59e39f147532a09669db36a5b56d8d6395e73650c5c60ddf1b64205b0a178e0e7c2aa3e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf49aed64063c6505ab8ae1f86c714c0c7dddcd3f2b386c57fc6a6dba929610ed46d6f37816b6ee8325547263ad9d1fa4683f19ffff7d6ccd4a0678897208d1c1fe66769aafac63d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf505031e4279b735229740f611a377fae33de288833f5698fba2cdd443e833a823033c8f31102a80ee1b2f81480cd64cada0383b1aee72349dbe7f0904ce70b3dd8479f4b6024183;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26a8cc2c9724d07dd17b86c33de9df885310c4d2a141af19d5236623a3071eecd580655ab94bff067ddd0ce3a72315d038349d7fc8ba158876a52bfce081de03ce13699a810cd9ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb909644b7f34bd3e262cee6e75d47932f51413bc5868ba3bc89985b99261090e15eaec665f1696b47ab6a573161bf9cf4fcc145df7917068b2472627c5bb400571d08c28ba747a0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had3836a2e1c51f7486e286818ca45c57147ff8780aa705e60081ca90d69410422eea2617f329c8b68c2c86f79b4c9d745e3cbfdb7097f7a4d8e30320c2086bc81fd8eab3c37bccfa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81af19e04071decb481fc51f70d47942bd01e7bcb30910c3067f02dd22fe6324066e698ac531448fae63a723537f331e78b45f4cf9862e9afb022fdc7a1d24cb3699c68dbaa00b67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97e50011bd14ced99ddcde3acc3dc6343f5c740f3e88cd4008c9d8652f98f57cbfbf17cde0c3bfabd3a5d37f63803f12166de8ec28184f4a16b2460d7a695c6a55ec3597a3aa1a5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68e1fed58ce136b81394793bcf8379dec22e28ffda94672340900bec28f62ce47d33cb82a8ca3059183c57cc429e887135bd3aa78dafe007afadd3d51465c1db4c99183253546dda;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46fa059169794af4ab13a61e9c92730cd246edc523bca1000703f780586b5163fb5db31eac0af21939fadcfad374a9d364463703cf763c5015754b616db3b69ff33a71887511271a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h472b8e0c2bf684af484ab4516933a337d0b1dfbb90eefaa3c7fcdfc0d8dbef8879f0d8cffd5218d5b312e981a9f9c5282a5cad5b22eaee588617ecad2fd08593a57e23f656e2b6af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heea842435acde26740aeba1b43be79285651242a40dd3f6202b433c41191725561242c2015dabc53dac612677c92eaceeec67bbe125a8adda5ad04f94d31607ed29c58f5b183b665;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4468db8c1c1600cde992da410e813c12792ddfca70b2dcefb653d316555e2f3ba6f1a36a5f9e92d6bc077dba1eff30bc90a210b87ea38e5c1733912a4169aaec30329362ef438270;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf09a9334e3ab5e8a9d9778d738d989dff884614e5b82aea0d96179efd80a39f38fc430967b9a12bf22630a956300c8a387987ddd6b1030d16140bbb070f1fd7f4fbcbd6fe189b792;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedaceb1d77cbdb1613a2ad6dc41f94710e66be99b5adfbf727d690d3c1d3372d5e80de1e8adefe811f17cb648f8f52700c3e1bae7c78207adcf35be4f62e6f7c2e85da05404b7ab0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h465f9610080d2bfd314d275a60daca895eb39abc967c2be9c9a774a21047854b9d08ad730d1aca982e9658a437767f97b686eb59aa2f5688bb2343411743e53dc1ba633442248b24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb529a2eeaf25c20e86d42df4f12a49399459a3d74f74aebae0a23fc079d11df108787213ca026c9227e05b377d1499026418b8f60c8caa821aa9ab606fb631bd6d074fb9ba2f359a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcfba1f34d892c25759b5a892ab2fff005788d9395c009e041bf3243e52fa6c704bd0b084a00151aa4a351ffcdad8bac4e15280be544e7417d6131a5f2bab30b8cd36e0e4a074145;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6417acb1ee938e0b85214e5763bd94ad549ce039f4d0633069a5aa6e531d5eea900949de4929ab1b0cbcc210c795fd1ced38b2319336f5ca228344bbd6ec8634bd5e7fa4940a1b5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h508d01f6b9d3fca00e227436707b28f5470c3cc54a6703aa100f2caa83c36747b5fffe6d67095107fdfe07b84d4c813e8bc78c3c75b6b67da6537d0be1b01d22b4ea6459a4a56967;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee52ceebada99fdfb87be03fb0c76d04852dd5f11fe877ebe8e482d19dda8ebe9d5c48e1c3f2e7c634829edb469c048bd9f0a8ca89b1c4781fb353aad9f6de8a9865c179225de161;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd716b2955706127ceb72d0fc7a15409d8a990294a4b0d99503a2fcc6587d8cda94e8fc16111966e191d7664c43cffa50a9cd6a6eb49edc37f4f42a36435cb26b71b124ccb1663a3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4151ce9c6886fa244dd420cc68eb8283c49582481fe744cd2900a746d640f2904d9da79e3016593790e4cc78a91f42a582d7c6a2531cb8dc1193c2330eb48999babbb82cc8274e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d3c64dc57b2d8bc8807a3ac590c7d165291006371475676974746ed491e7b23ef7e3059deba4841185db6b1d78385069b7cc9fb1bbe3d98e3678c360ba500f007ba2b25ed436088;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e693c27839838272c57ed8ac6677ce6606d1eda281b290860cb47ce5f5fff027946d88d20c4c247e4f76f164459ccb74d5822480396d44c7079ce4ebc1ab1ffd457a643ee70d575;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fc4fdd82ddd09e8f6db65412e757510aa81d5f60e38a49d6d3d08bf3e8b1737e442f59a7c32eebf91f47cd192bfe34210a7abd5316614261206243e6e38ede36ec1d1a159d0bae5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h120bd9bc7e97416605ac10116bc306a911e4eb9c74f2f264b0d650dd7a1952c2582079927a0ef00c0accd4a9f9843e4949d20fea220ca805da00e07b51e2d44ff0f69f4658f18c30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba524d1a87afdc2ff213ff3aed1d1e632d5bbe6196384f971c76fecfbee36a43c89207a51789892fead89289f25a41b35a1bf736f8b73b948d907ca3a4791d3e2c7803dd8915c051;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h669da3eeaa70cc0e262c3612beb0ea24e81f06968a108c53f0fd76203b2060a7575a28e59f648cba972e140c9cea50f85ec83d81dceae47cecba34b92e8abaa8528fe8ca76623f04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha49969c5a67a0a52faa3eed549d9655d21c19497c94da8e5ac28b93f41bafda6847f5a955fa9c1b9bfdd37cfb8e2b2a88db4afca3125d51145667e3d72bd5a6fdf3fe256527542ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c07c51460f0264bd12b812ed025977271c00dcdcc1384dcaddfe169796653e0f5e71a9ed9f3628c4f27e2fb3c3fb2d517caad44a53b1051b048930616ea273b67a8b81d14d859b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ca9467a478bc3e314d4404923531693614ac7a2120164938d1d8613769634a70d3f0ac226d4cb23a9ce5645bd4edbdc7650c755373189c9ba9555d19755065cd1736197d85cb755;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3742f851bac477322d63fde07cf9d766e2a5c55d29a714077f949ade86f6122deb8ded4efefae7fb083336f5350a6c143dbac8fd5a0354dbf22ff223ff8d0d2e3d99b634d2d0e405;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cc54b5ee425c07591f92b240dda2964b9f6034020022195c62006d3fc297385fa8668d776856cd27e173dde1be6946f698434817303a97147805ff3cfcd8353af8ec2b0f532b6da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3aab07b7d815aa7790c5dae3df8180ec1611d759731325a2a6bcdee1fb8bdfbc52c7fce0495ccd512c5a972b5a6c97c6c04df994d900345840bd61cadd7591c2c9fd45d36a48b2ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h644a8bdea8bc242a58473aa8360da2f4992f874622567a111a79661f88cc9fa84905a8afbf3eb34437f743b838d1b8ca3eef3ff8615f26f49c1c82bd096475d76ecca13469a3a4f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd26ae49751cb2b97286b1f011b6905c6709c75bff53419759e7a8859f574e22aa3a3ba574239b9d97e23a84ce0c580c8edb73d8d4146d5f9f880e521f4c95f6e43fbd1a9fbcccaf8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb19cb33ceb01448b4f7637f722e78b6ae88512c1899900db7351293f00c278e782cdb93be35e305617395178b82d29f1f6cef0a4c898bacd0baf780e24151318bdefed05e6fdd33b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h576019637d3c3ce6de7db9acf393905b7030dde1612e1bd1c062d31d0c5ff1bf01ccab3b5fd8fa220dee88b066455ef5fad2b27bf47887b44d2d9aed060a0a809735c062bb99bfec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca5818d3508dcaa3d20642ceeb0b3e993b4f19b7f97666435e147a600a2f195e169731adf7148cb19d395083e086b985d6208b03080595e87abdc35ed7b62b0ace5f3fa256f78eac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8ce08fea87a57283c26699d16e2fdfd132a00812cb1e73346307f7fddb9604b6fbb62d3031b61e1b954ad1264d84e86e2fff4f64020f744beb401608d652a6f5e389fc055b4a954;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h837aa230866110f5563050fb0e171f0180387515d70eff1f1688a5a15ea160194b08c5ee7e7910722b24526dd094ae8574353e919eb5ba33f47c797d42076a286e4895a042869989;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14746a94d78d7285db67a1b05258329ce5e64ff59c4a4cc5a01d36daa36ffdcbcd9756e69c075ae02b66ad2458020b38f5292ec2db45318d0db91d72c924bb639be132023f3bc119;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c035af118cdd00a8e2b32f54fd217083d0c42732b9feb18221670b670415543d0d2e66ea374b6841be2e5078e1ff0e4a31aad891cf058895f749adfdebedcdff3b48b3add4b05c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85ea56bcc59bf54a234b090f563d7dc89d423b742ac0aefb86d78100f119de1c26041ac74200ca5886172cb190b3ac127d24a61d342eb5d237af57399e1ceea2476d9c7f446fd475;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1956944bd5704a333645f6e34f00ebd48de52c3a3ae4c4674daf11ecd948ec3c01ab09031dd40d86ba5caddbb03ab63259256d829d8cc9f8ec044e019cc97bf67638a34c10bd5e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dcff921f394518581933faf2494e77ae8b3ece21d80a5c959325f22a079f0293ff3e89ae20a950b2961e53b22213ab0f319b91c4260a57cc2d21933ddb5d96278aac811560a62ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcabc33ea6ab7276961e1ff735b4e26736585108a2c1c618204a2c00854f0604b10db1797e4441d12bfacd5a0c278162bd3a9391df5066a02437d24183158bc84291efe4dbad70c44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc5fa232f63c6fa3c5d1cb5d03b84c0187edf0468bed84243741b8ebc6ddca08a97ce9a9d90e3f2d85609d3c2bcafc67bccfd4c543c3ae001b8978f5332f06d6c5fbbaf469ad757b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h770925bab513d24758846ae7ede3bea448afd178f1d90d781e6696676dae02e20140504933082b8b2249258e68eef6363893873c34bb972d115808f84113329965725912e228cc37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32a34d11f29b8aa81da6cb3c2544170153970b991ae071683bddc87b5090eb24841560347b6d9be2fccec6c09de4b68bdf4a6f62aad21a715461e2cb9851a05addfba1fe23508a41;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6c212d0e2c34f1f8cd5c752b1bb639e0b999d85639f1d9bbbdb76a994d410bc266d1e3f091cfa6ca026729be6ac919d7336116e4917700c11e22e5cd4816f9f1af5f8e6528ba1e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h606bfadf088dce6988d95305e2166a814f4468365a9b7010862bdf3bc9a3743b152ddc620a989a72584e3ff5c085fa180ed262e01558c126c437b4cfd1fdb5d057632cf55d2e1336;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74a97646014bab08622a58ef5ba00b92f3c3f3172ba4d6e79f00e1f949dd747f6261a19ae09682ce42e2f440273b1be58c60af46a07af8508f5fa5a9abce751c24ccf25e12f43169;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95d1a391019b7f308fed62be3cd4880b70902619233b58b1ebc36ee5df33f83a83f96c3f6a27b92ca8d41ef4630333dff1b41f7cf7d5e6a11833446a21d9134a00fae74ba7e77d6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf75c6087d9aada2d9a01f38a4855e76a3c4e830fee2d2204d6b912d85d43c86996f13e4fb83eff97937e83a620b402d3275dff85ac77208a8dd913cfdfacca184932d12a601cdfcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18c0595ca765c5858417fb6ae5832387a38610f4a55b6a10ee3b969982849150aa2664277c3554918ed2de2fffb22fd7f0f74087123f3dab1806b2e8060f6deea2aa52e3948e16da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a10a0408fa26a97b2f799eaf107728b637d229272e6daa8aa7fddab59fe6251daae2aaf7654a0630bc8c163e60c8f0a0ea947450773488c084ccae874690a591c31f33158a4a1c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf890c8b7966f430cb274d4295c8414aa84a55cbe96214895f7c35fb6eab158d8674a37a108c8c9fcf4a09b386bdcf5596b091367f07980bcb747724d4fc6d1d24fcbec5a0821e572;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf24db07ea94beb055377d08fac2e573151d16ffd63e6acf5d9b931e7be045186639331ebd782afc81d2be6ccec1ca70d8b8d0b499281401e5d4b64e5e9bd1cae93ff42d8ebf00a2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d2a1609968041591ebda9dd6c1869d595eabde5f27bd0e60cbec550cd96f311e806e8242e52cfff91ed22a002644d902dfe729770e51d80a8c4781bd7aa5816d4c36ca24fd4cf08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d506d3eb5f2850631d10387be20ea3350bac57e614045467bdd60c32823d7492e2f087e16b9f7e9af2a11b7937ffe43fd55ebff4259f04850d650cfddddf2c37d9406f0bfd27ffa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde18408b1e7ec09d27bc983bafc390a1111621c5d9d3b7a0cb98e7a40ad83acb65f145692af7b3bfbf26f87a54da4711cbbe0ad79ef475109ef93839342f1f1c20c6b5137a5b245c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59419c46123436e499c4a594531a85f924a1c3e9b3f5c323f0dce9b68dc79762ed65df75c125f36ce1ad92d718b70d69eef1acfe137ee015ceed3a46ee5b37c0389d89a64561d4f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77ace5107b54e67c2e84d53f87af5720d7d221e9283a90eeaa71df3a327216fa4c71caba357931942992f9a669b2b4f498f3924abaf341cad57923fb75e6722f4cbf155f8ebbf6a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83474ecbeb029a9859765058eaf32dce6a653760333a9a077ab32fe0a743bc6b6cf7de0a49b8824cefdfd7fd37201b80850e9426dd427f4fd562a76d4f9782528ac60b1f3289fb44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5346f9e61f23d8b933ca6edc457bb45dd9bcfead424aebf16c62e893db91b4a6939d497e2e8ce71332f1d2aa56aabaf2bf9d80a0d180d0563c1e7d880544259d43f13fe14d3af4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37f3219dd86ef05db0da2725192f348850a807e6028a8a6bfb5529a0dfca665281679e15cabf85cbee0368f27d6947dc72d06648b0d2f348c03e271d3abd0e170095ce4a2b0ed802;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39519c450e04a056369ffae9e7b8e3843cd8b9355521b0e5622b45a0cc7961a8f65ce099b160c56b5885ac5ecb7c03578c2bde812063de67160ae1214385c8da63c437d3a3a8df05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf99a09b57ad6b3d34f9b75a6b3464dc6061dc34c4e8466a0f58cb1931a9d34df8a350d8d7faf4c59d56d2f0aa9668b30f97aceee87c42031f36be1896db46d3034b7a2283143ad2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0153401944990a9f87f2fe9a942fccb1b13193e16f6cfdf04431381e987df73b9ef1f7a435bad88de16a617f313ac0c048047de20c402c850480b5acb77e6091c0b1b679b1a15cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0f85038ad2aae10023031979c3df440afe669fe4b06a0795d138e6ee7d7bf57806ff58053c5dd88e85e9f4ad235414a328c16a7410513893469968b942935300be7c68b5561d137;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b355d1ab7b75d9aec5794c3679e11f7fcba59e2ed3f19444458d9cad86a060ac562228b506d952a690f2ece5ac2ed982cf39058607b643687a10f92066fcaca04c0b66db960d4c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf15f28c17bbe6f0b1511b9850f451b0adba33adef1141fb2910a3eea430a0dccbd9ceac1d99e9ae5b70b1f8558f02c54d63ff161c1a38a17375a199c5dc6cc20cb8b7d975adf893a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca1f346a46c25f8a4f57a6c0ac1cd1c9b33da418a82ef56bdc26b4dddffd3d9909fb60e7f79d7828b625d66530f50f77d09640bedb000bcf6acbc705e6648ddc5cec5f3ad28e3218;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6171bc7ab2f559f36f0db90c01e41da7b4a932a495515a7b9b8b7ce1fcd10a5929d2249bec9ae4d8374ae82ea32992e59c5d529f9a9e39474c58848237f827f457a00398b12668d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18caee6bb483a7e34d8c924a821ce7d73f8be0e3197393b33d017eb484b95406dba8006f6b6b8c46c574fe3fdc0fcfdcf2c089ec9678a17f92204acd676634265cee7fe359cb9221;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he099070bfe751baa4e17951b60bae5dd533ccd2f129e243f7a010500d0dbfdf15fd0c2b8cf28427d32373e99d8403df9add50d9d8a12fce80911d7d4cb16ddc266266ddc4bdeb638;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd84bb2b94f3bbc39d1a98e049f8fde3317fc45b9db7dbd1e07c5e805e6dea7d137f144255df96c4061fb6b51feb9c0d169d7026c9666c1a7c7f1ca99790ca569dabe2954a6b25d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7de66cd84cedbe6e62965300f1e70216c21b7ce07b32029f6ac0b000331d8e3336da43b75781b0b566aa909cd133a238cd1a843723cc7a5b571799c025b50192e1103650216e76f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f94af87f78456386033181f5d0f50e6ee86737e6dd3023d8b275f85a1c125250f15d16499dca51832dfa00a6a9021f1556fb3879d510e096a37b975fe8c5135f1a0d4c2bd3ab2c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bfc78d19b730305c9989212e1b8b350d10498cd9632ceac8469c0211874471e85c9034d5d719e24eba557b83874e00e6a579fae559f6be79ce5dabc66b1e73c9c9073c22ef66a2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb10af20bf496aa16bfef5cf671182f4960a5502ef7849015c0935a73bd269f6ceaa7dc20905784296659fb72b2c50a16f5ac6698cd8c6e27828422e5235eae0bab1dd7325e8089ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0079efcbfebb5a4479fb7c4c6d16efe548c22156403ccd8a59c666d8a84694e47919ac06cea2b831ed643c18887a935f327e7a5f1d6ece0e25ea1319c24d75a5a5b995b5c35ff4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ba907df7e6fdcba5b203a6e93a8ca06a0946e472bd0ab2cfe69b7b71182999b676655195ea1d8bf3b4f121549e2b197162865f04c8c7140a5cb579636288dd57dadf3e0ddd0ab67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ecbae6e91d0c5cb016d17ebe426ab5fed3cf7795a7b1ad433b1afeccce8850714f6abe60d493ef7c3db4e95d72ea24475d046cff0a55025197a941ad9238a2204de3d017fd811c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8beab7c0243f5738eedb46e062f2a5542db6f375d896fbfa1dfb4fb7f9a2c753ba273db78251ca773d9365491d2a7a97dfee23d337e1b94aca6bb6f53fa3954ad9c5727184e7cd9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haac251c96cf0edf310e9166931575d28f5992088f77936553c19e33470c5dbb952beea874e94bcb5a1c6f35f7de005cc8fffe06a062d2c787d19cf1bf6b9b37b4b36b7edace4daaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h793fc9cac79ac45f954f69970785a85095ece872928012a4166122778b0ec98e599480e27c16ef66d0a39f77d4a1ae5c2bac136f9477d0918091df5b44aae6fda8e5a62fa7982f1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7f91ca067d2fab35dc2ee9ce798e586c7dc83fd549d19549eec5d817464a5250189d80f5ef7e72b496699a984001d27160b77845efe3bdad1070551fa31e6c5f5202835dc24c1ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323ac232a14b8ce8c2afa5adeed286767174d09c9e5504d76b66ae3fc7dae8d4d0958fcdbcf9b8473d2cc66580724c0068f1863a8bbc1689b436a03ee14c122cc48603e61450ffeb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8cb493c43906e4d0a8695ed3a08e6887696f00adddb977984962ed8d802106160f8754bb33dbf7ee420a1c78c3ee717dbad0dbde2f3a180f047bd6ed8a5454e0d2ae864bbdedecb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h785384b43be55b9d96109fe3ba4952a6266a7ea736a80eeaf7b8faa9c70a79785b86474cefffeb7245bff236817a9f139524229e0f637b2fc74be7ff721d2d11e4840ae361bba580;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50326e55812a0c211fae8f1faac34335761574b489ed9580b9794db2cf5d21b6c44372b069063c8c702587ab1b7f4c67ea4345eb7e42308c8f65fe80183b40a0e38a8f0e3e7224e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4fd78f12be0d2f69f5d6fe8698fc8fb923ee4fb72e2c20001cf8d6e3e33e1597537c4a56b9445fa6f811e2d8fc5812e4afcd11f1669a1ab26a5fad05bfa3e7772bff68097b4237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea5a6703ab1b1b181f48cd567321b553f5bb81c9e197c8ee89c752a46b961208b7d033e237f8cea3c3a244b4ca9ffd2d4e1a80345481e96fc500fec52064f6ac29726692a212429b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6eaa5008e51184f5651b1779f7281b8fbf35314689a0429a3547726c07e5d73c19f9b394fa28660c0f5e9b4fe5f879c4c28bd27cf99b5dafbd1c3f8a2c8efb4de5fbe218873ac95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8a9b3b5259e8a073730698252938393b502d5ba879feecb91da137c588fa0f4c4706a7f87010256b0161c548dfbda7900990f644c8092ba72e04992941310bcd8a6924542d27eab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc24869ae06a5b0aa66226b2ea82bb0f3e0d4b67a092a23ec7984b0d1d6f5617e8d56111aed1e00b8acc202a27db121f7ff4029f695a25cb4660a34409ae5afdf79eb32472754a769;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca45d6b978e58193cea9d0f0be6ac8aebf216f8f3bd180b7dde6dba9f48d6596d63143f4422ddf650061530e09b462ef80099e1e90c552d765c4f348e9a1d17104b92e33ecb18987;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dea3f923e9523a8a1e0c99898d6811e90492f72b77d5dab4b82719a98501735d6eb6e2d7992d4361de265b45cc0aacfeac3a59b2a9f418fb9db371a5ace41a96d78c91dfb319d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c117554cafc71b4d8d5a49dbe0675ce6c8597e3d34aa37a095cd9cf2d48100bbec4ccf488a5999e1e0a9bdb5bcd9a79b5b4777dc2c4a1daeaa30d1457b6d2af142a5dd16533ad97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27da15d23cd99d1c216e2ecbcf200bb3d5fc404f3d2be0797820eb2ccc289f44f584fd48f894731ddbed175702cac96645896d76da5a750acfdb299ce96c79b0e12028138bf35d93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9c1bca1091770299e8bcfbff6e614a9be3257a6eb45cb9d5bf47aae7f4db091c3046ac59a6880fbcec237d7874ad8881817b3ab36ae5593990abe931b8ac57d8e672421349bfce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f208165c2277b994c2ce99c770a10ed921f24abb67d7bf46bc14ef49a94d7ba492d4f791d9bb2b7a7f352aa25c1134d589ca80c19ecb475a3d308187533a3d486bf235d1048ae85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8b00cff7055aa50b78cf6d8bd1999dfb32551c8fbe85065f8a0b32670b566798347d1d6cfd821748dd617358a0440e1b6213fb1592ec9c394003c85b8007fb0e2b0e28cd3f4edb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h600918c430c59534ea3dedc582824f3aad8aa0427a5593a5d57674eeb98fe05ace07e8827dcaf4a2d570d74c8b8bd58eb957ade9074d0408f75acd7556c9efbbd8d2c88270430d76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc91ffa2d48ef3a122170c377390fef723613f6b7ff035d27bb8d9c331a41477c8edf4e6e0dec67dea72fdedc8e1fb45624daecc487e7a543835d07e4d0559f86fcf0842e49775e07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h647434d862d80b4b5d96e6e938750d0f86bdbead8610423170e1566ef78d176b7f247f5c9ea75f4be1025538b5753255e557a2afeb6747624e6aca1da4ed6de6c8122d3a0236791c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a9317b280f0aa59adc73af3d70621052de516db2864af717e31f0427e1e1e9bcf38ca2fcc7e0ee5c9a9914aa1bf2c413473de7c976ccd1e860a282070387a8c7e102419faafd55e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e8a44d060353d1267d055152dd37a4fbf39e39eb753a2da667d25f7dcefba7618d025f1dd1649cb9fe437ecd03635beb4dd53e63e8d45dd02ec034a2b04657e8a3a0572f2d38178;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed1d1eef9ac7bf105ce7ecc6946b7cc1acaec13f44f619a3e91cb90e44defcdbc713949074b1ffcf2b89ece07c9005601f8cbb6fc24e6dbf5cc5067e91e90f73cede9fa1b9582d12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5c72b111502512ed9772829d3a8ff43c028557cd709627e247cedc6dd9cbf256d2a27ae0e4c6fa58b093f0f11bd569caf0b409b0645982a97a4bb7cc8c358bb6c1ae927339ef67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h686fe4f5084ff0ac869cadb36b5c3bcb31906ac1caf80ab45045d371128015e0851dd282f736987af652f026f7048ee8eb662a6f6e4db15629a09748655ebefe987d6897fe94f2b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65a09386d32a2b29a47c939245ce0b46f80605dd16ed972bf09492b220553ab421c886b646ecb167b27849022afa26053e6e78cf3a35ac332445f5eb62d3a01d4350e8b533510366;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b80afe9eeecaa43739e4bce0e13c0773241c8d1dee22e4bd84b67a7949cba58b3a47dd748508de825d7c07f52e09dd954a08b4f46739e3de28e3b4cb757c7d2d553fd124beb0328;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefc4a6c60da0e36204c500cf840e0735202831b4a186701eea4a0c1df9ac56b48b9f4f0a09f6300611400481d0167a12c5a274d4dfeb1d62094bc46a5c985433b722183b94e41b5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf269ff1afc6a329c0f0e73c022f384d39ebc93e676b2598463acf0eab1af4b55b8163a0a21a4cddab84b458e52a59da5bd17da2ba04ca7295da37cb29ba2a0019fe18b7c845ed956;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb276e622af3c3c8597eac47b481a792defbd67d018bcc0e4531d2fe227b7b6d132316f8bb8029e1422cee9ff4e25f7317bda0354d3e24459aed88ff55355d2c7404d23c9bf576a5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b8301cf9d5f5e0c61c1f91bb91db5d100b2a066e9b625bc0960813c89d173ee625aa932240af3b273f8f0ac7aecedee9a07e06a4670994f9d38332c4c33a4a38b0e7c890ea76881;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cb19af65b41d87c9b235351da9ad2020d932c274c17d8ca1f13d854199d83f8495cc1b7a587c12f2d8a039c948f0cc5fc558e3760c9ec9c3e00ba9d4fe526c0a0dabcfb6d3fc72f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4132e54ef7016b6502a2a2911d5e279810f785a7d692f8d184af674a4716d2848cee6d7191c99232e0a7a2cb09e32b8b43d39b468b58278325c63dc3d30c120e10024280f666892;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21b448e8119728ed67fe08594bad28a0f188f23b9f2785de75295a120561e6a5c6f59ebdc29d83d5ba225a60a4b53c3314305334c4cc821c07ff70235617b394e2537ff8c8588a8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2118256820de108f866f16b9768fb0ee55bae9f714b8a395ddb8ce9c176424e3f6ef91eb015a23ad93bd8a580f90d5914410c79d4941eb7e3c29ed6ace90bd93dea0580be8423355;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c0bd14cdca34ae0886677303e5bd8e69a15297f1f390e5b189d699b247904f48bce3158907a1eb49273b613b257328bb2f49a71f7fe93adbaae106e25601fc283cf6ee01c392758;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7fa7d7112b6008b57b4037d2b8058ba67756e23a674f036a67460164217f2d6d880afe0d52392905261061ff076cfe485973277b8a831961fc914db29fdc195cf28e88280a0fa57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a73dc20863ba366bc082baa9c3fb1b4af04f7f5a6640824176bd684dc81a404547a1ecc0d6fce65d3257ed293047dd70a4bc4cd91be6675b8f0191a3088d7c46bd1c96f4143bc07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e8c8588a086124cfe248b8a40e6092a1083fec668479c69b9040dcfd1b605d6158ab3e551d9186b7edc719eb20061f0ea9ee2b8010306566c3d7631aa1e140d07fb503ebd7fdeb0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had548cfb1a3c15810da5aa0af716e39796e5a7900a061c2dafbc7d2f2ea53da8e4b6ece250d1f2b7c9279fee6d48b85b890dc02d9b53d8213868700a53cef20bb44ead75347d62a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb75c483e177b5ad051a84606a2e5494efd5020f5d31b4e3666341c57dffa29b68f06aefe137fccec0e904e939e747603eefe7a616a6b8333236335ce1f89b9667f60e00100caea68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc45ccaf404cf706cf14e9d9dd810c8e3ceb401155ac6c7821606384c1716fa4e5177756e1eecb06741c547b9481735a05fc9d5495a8799be158cd23778e8b79c8abaf9d9594acd63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h183b225ef924c7eacf831cba000f911cfa4855e9e4bec8c5347bb7769a3bd30a82b0f4f568d9f0cc21d8d230ca14831309d0dd7304c8c7705a6d0d13e0ee15f6eb1bd12b9554a7ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h625f911aedefeacd94f71f0b9c31bb48091d0a4ed9eb24363d256b8aaaa5b1c76e161d10b18fb3fc0872b1fe68fc698b3f6dc1df79ee47c0c4d652949a84b0badde52690a743bc0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6930c45208362cffef6cf8e0772b4b403a870ab1af96c03514f8497b33b26d0c1b7e3cf343d5fa069800335e7e101425242177b642f782868f26c3da1c41d97ade259f71c4c04b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26363c377196d327421fab71859bf7fa014c0f1fe815259fc7e2de8dc34743945bc5d9f0b284c48c7dec3074de8834d5bce6d87d19992da1566e18a756042184c8e2da847e68fa78;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h761fac3c39292155893a5ccf2a212f6c81b4abe7148f0d179eccea864e6d8af5e349842501b8219443fa9243e23bb51a10e1dffcc4c7951dcc7890cac1e2205bd5673279124abcbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f9f18345120e50895fdb8431a121c0fc8141a458d45d1fde411dad7667e51c486c666efebb2fedcd6821cedca196bc7b3abb51c5b2ad1596348274682a45c726e2567e6299aee05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13ba0a75b5c8da22921a9ff3ade0d27fe52d550e3830737b764f9beab9291c399d5bc23aeaa507d3d6da41262dc5c0435b65b971aacc89fc3cc7f20e30e68b7f16f49a7c2d5e2a9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h579259417d6c601c3c2785e1518fa4c75505e2b529e254773d01c7804b9c7e65bf71656fd499b9bc459453b4fbb1ec73b817e11237b8e62e8bb99c280346d9cb239ebbeeefa43d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5729b31fc20e6e03cd5e743c5bd14609cd5a04111ad8726ec3791f6e8725a734d9af00071e9b9eb1cfc5b8c2e5d3fdfa0a9e5adc128d79c1e8beb7064c3ea452bf0506dd00dcc1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a59ff318a0a8433b7bd210f71b9e63c276597ce5cee88d0f78af607fa00fc0309306ee8f08e787e316df7a76b1c0943aafde59a456cfaedbde37240520f6ed4f70b548258f0c024;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ca955a2452416ab3b55fc1a862bcdefe32b4ad91aeb1397ca6ba8a393fce8772f1cd00cd8f4be49b5897f0679f661d2f7487fb4e4eea66745642a4bda8d59e859577bfb759b5c26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fcc34c477da9956de895d3b02acf2eb282c751f13c177ae7bbff5122c1b603945bcbf13e6bf843b5149c5ef84ecb1320819a052bfd61602ffd537ab9e9db43932f1c79cd7f8ee6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91bb917f2804521a3f917d1f7a5384aebc686a4ad277bfd942eac09cac54baaeec9d9babb8462bbc3400c19b9fd5c08bedfa675e3479aa370b0241b6cb8f8e829671fa12f8656da9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5526fb42448c5358de9b0713170dabec371ee383da382f336257ebd3ede6dca34c530849bdb329ede28499dc0886f33d623acfd03d1909957148eb7e05711761f5f2020192882d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha337d68ddeebbd0caf64ddc1caa6651a9326f508924fa874d5d44c3960a38f7e69adbc7babf2ed8f93a1e57cd08c7830790f16eb4733aeee14eebf272ebb1789c7cc0f8f439328ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde311a69cd1e7bb486a0329fb860091e5c8510bf0012fddf1968687e040096b961e2b8c52faec2ea442b24c83f14e8903b3aaca49b8cf6392e1adc294b4b643e13347cecd197aef1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c1bf1e557f4839593d55769ae81ad37a302d1b207395fe06b40f0e0d4b8688ae8d640eeaa9c79bbc22bd1987fe8cd0c04aadaa51608ecfb5a32081d862ea6db964d9c3785546976;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef8289077d063572ed3f51d524e7bbeeac28d912e131c8768c61e7ced0e61d088396fac94630f6866e9c0c650c058e7bc707f5187e2b40c7231ef1dff294cb88f0e6ee84da5dc0a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb55b3a3afbe8790120bb3a9722d3a2d89eb41d63d29d7846f06dada4d963f1dfa702a044ba37c2d979d94d2a20e5b066124ac6ffb3c4102df00c28a4af7569082a908ec802d0d5b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h967daaf6232b01729854c21ff4f9a28b36c211a2163fa187a9efb75bda879e81c9a93fe5c295451570d9dcafeb0bb8d27d36731635474dc5a9eef1f1adca8006529373cfe4fa4058;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf50949a5d1f445a20ba8f6d8796b07fd38024250619603cdec46825b47a50275890f2f736f22e1f3cf87474f99ecb0d366fe03f7918c92418e208bc796a49ff87ae7ed68856d180;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b14f00e733c910fc3b4f899e85f7fbc0fa927cb95d0e0f1e08b25b3186b0a3a104e66c4fc66f73546c5a5fe73bf0afb71d8f410215dbdbeb9fb1fc612e57a2e81bce728e2d380ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbbb2b2aa58767fe3f66e29911380277e94228dad7c93ecff489894532f6d836a53051ad5e89312afd4ab2dd9a7e52bacf0b228fc99550de4ee763975eb0aaf78fc2ed0bd01883fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h320fa9eceb2f2fcefd7c3005af242d1517ebb4b8923316a4a754f969436ed2800898b475e41000a5355e7b6fe6bfecf6aa8e82f47d53d01bdea4924a27bb4b5dbf80753a264bacfb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60e9eba1ba2293c3104545319845143eee4f841dc4a99aef4c2e5fa797f996a0243f775e29468ebf5cd500134f40f2fcd1827381db5059799ab248cd5c7d12f8799960548821dcd0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha37c978171e4931ddbd2b59c69e3e3bfdd1e06a34852f51d22fdbcbe4f34c9f1953129b1a76ce854ab67d56aa211a35fa8da2c0030fb33bf56a382b68d06a64a241e699eb8537945;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7edb4c45b68f84f3994a85efdf952b93f47cc2df08094ddf01f5dfb74ff9708a892860f11d2df4ad5a3bdcd681a83aa1b625c7b16c32348f2e3e895ae6c28abf32a80094e1c8aa5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8ad1fde62d7c8ce371b10c245154b8dec50cf97bdc70469cc8b4f32c1368e9bc38b8b8a3c5d7077ef36147286af59f3b95659eb9f5f55657ab0264b8ab89fe84e25726d9fa342c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefb8f58aa9bebafb67d1f24f488b45ffda54428f65b6812ed5847007b02ca796436d50611002ef6233ce357311770dc60ea5dd3067d162a37cc11172815ebb0845d36ea1032c055a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2391f0b8ee58942686efa44cef440898c963a765153ad0909d44e8d1d848139e47670d44f61d7ab00999fb7f701fd37e902e5a50dc4acb39b8763167c8f434189c54e6d8c09d0f2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6503d0705f1efa5adf35fad95d8125620e73d9f76b26bc79c6f596ec9ac066e0ab26ebd9876df99665a9528bf71cfbe03c13aff3f4c93aaa808c0b7b4a5fbfe19a4f0e69fd392ca1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he67332af75e8b156fcb79b4985eb74f91abdb1921e02bf9fc097a37252219e9082639c274ba5cecc9573c5df0b5b540148110df68ada24373653338b40fb27dca37574ad07670fa7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe823f60e1790b364cf063f4dca473196e76ff6ef58bd4933f10acd07da46e79e474c5964bc82375353549b1fb5252f4a72a8fb8ce0891445abbebd622299ba1629c077e7195f480;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0ad03e34cde328d90530f6f3d801e454b23ca05f857001e4eb0b36fa07d87e048ad345594e66d40e14d918f242d91b375e6c20b761f198f1d96a04fcff480dabecb3eb8e9f531bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5987aaffc397975aa1aa04f771f006a0c7592cc92c9809b780a5df5531e1865b653307ad93dc47dcfbb816f35081c74a02854e7b61f54003095c77544650496e51bc4597c3749825;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb97c250f35d198264af789eb8eb426a0d69e076de23a5291952619a622a3349a446d21050033397291423cd20a6b946cdfc96cfd7185cd360e64328244e76efe9c1b5902d31a16c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32a12cd5197e9b309c4be5480ad293a020696fb34a0fd330525302a1e1645e0a47b8d82b980da2025652070daf7db76ed0549830f4634f96858e2a33496a32ec29750e2017c8ce84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22def44183a92cbab6d6bad98065ed1016e9e54115487f587a1f56530ef86b53e7dcbb2c4738f8d886a24ebdc0b621e6de31be87fbfbbebca1a0c4866d192ac27567e973991cfe76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafcac15ef17cefb39959606374bec2f8457cf5bb9357f74ed09de5a161d447f0c83a295576322d58fa0f00007bdb4fe82f238e6fd0f949ae6cc81108b66c84a4224cd3d4bcb3954a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h214200b90515d6494eb09b02cd5a73d589fabb39d8580ff5d5d5b95216893bf33a66bf3ed9ab606e9f1e585af01340abe7baa5d9ccf3c6e1d1832ea779f7d62ea9987c7964d7aacc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccf5837d42b7ce7f2c1795fd5a24b504d702c623d9e508660cf07e0dbe42734dc8eb7b243d47e4e6df841cb0c05eadba37b6c47bce833595d352089477aeac96dae2e64ea73e3a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he51ef0fb5235947dc2df0398fe60b1f59c5fd8dfe1460db02f8f743fdbc737f7f9c63d2ffcb69c26c1907753ffd2d5ed26b06d3999c6612e256eb0465bcf8236da931b6588cc3c80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he861b8dc0682dbee03816c33364da8f0b29948442dc828e6af687a66b79d31bcb063fb5365aa969fd67313e992eb594a682673c3b330e3cfc951887f7e30212a93e81deb39611c8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b912451000e9b04740820a2bf657d053b0b638b2d7d17f077974a2301558c6d86c0768c6ba57b1ce78f0fcb574454350afa1f2005bb2196d031f201f86ae3de429614d24b801272;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f263be301cde451e74e7d5dcd13c8a4779e5ec1f0c635fee87b969fd32a6a09668b1da664aaed4d0d748ec97a8f2b9931486d53550982258de2a03bceef1febd595dd4e3d733e12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfde2fa613171d2fcc1d93c72848d77a722ddf3bd32a56b64d3f853693bb38561c43863f5f416ff3de2eaede8341aae1755b7aac215b809c2c4945b14f23a6af3f9977af17c673e83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86c170b1db83f33cd05c188434895fc32b83404c8b23a53d3486f83f92ff05bbf128b6a073efbe98d1ed983f552cdf811c3335d478ca764b679e5f23c0526eb741c003f1dc47be8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf86ae50969439f8273be35d513567cb70919fa97498307577c7c910940478ade79ed73f27601695a3d9bb28da4af7b393c0ce897718feb81ead87f150a976211a87fc78ae4646aac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf3d19a89cd3415c8338a79d1d86ec11e54cbaa182d17875d753528123337ef3d04ebeb4ccce3b37ae697b389bef1bc5684f67337de87a896be3ac281243b5198127a27df3df493d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22a9f1d0f6afb2ae1eaea589bf9526dcc6ec076a77b2499ab38fcbd846f9f9f7dd47dcedc1de4ad01a2d711043f4d42f543028a0fbbe6789a1816d6b39911058d8266c0e9bfd70a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7aa21985e4c55f1a8fd6067f4388364a62a89c7d5dd4ea28c0350313c20f89b706fc262eb20bcf014eabe5410cb40d7a28c19099bd0339711eb7b9b608bc9989b4ad119ebffe4aea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4333e8e7a4cc16dbcfd796cea426cace58d3c2214f924d4f96aad848273812d52e94a2f605edc563edd96eb3fce36bb9d3a1ff2544b34e9a62ba8e8345df837f305de81dcc6708b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ea52d2c4c9546d32905b7e8cb8a9422d76a65fa9451736957673575d8c74909726cc7bcd88af85eb9abb2f24ad4ba6236e10f0ea216e7ed37f507a40ec0ac545fac048dd8f87f49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h394077b3158a78482e8fbe7ddcd822b3eea012e69d7e5da80b144d99315f70b32a652f94928f2617bde56529d10fdd9fdfc8cfe112db45e16ce14e76ce34db4024e82233ca00f18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h830c5e81ea5c1408e1a73f9d0072a22f1ca22955c6ba4fe3d707384391479deec192453455b946ccee97fab56d43c6ae6a51261760632ad1235c44931ffe878db6c8fb508e76fa35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d7ae7fdec5f4fcb929ccbe0eb929c9ea0e7c4c64e54b947d708f987b3b4f0acd08fa9911cc1541928b999897e7f00b2ad164b8ddf37316285b03b80afa3cd59510a73c58e58800;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf870ce953aff8bba9dae170a223897808c3f585ca4f5abe59ae603d8239b52fd1b1b585e40daac49b990f09b17606ae6a500bd7afe649620698b10806a70b8f99ae774e8684f0b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf480731df9f55b6e5ef1effb303ae0d0f0d0a895f7cda9338dbcef56f48ebe9ce326261bcf4e02ac3b854f1c64d5f841121ebea9696e58d48ae8a0f811607abb21ccfcc5a43c123;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecd79afe4fe9b9e5e59d2e5e174c4ae38f31e35a55657ed6a019438e1ca808667535a920ac944230296deee5aae6faf7b0e6b939423276b96a7185283669468f97c2c29558b735e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3c969aecb06e9d5213163986bc3749d32d9e7bfa896650b48f1698342af8eafccbca3b87d93709d4560516602b77e8c7bd5e1c387d9cf695c09b8f6d1456500c7b303fc5bd2e2a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h368b27156d41fed8892e9cedc3d94c08b34f8db4d2ba496461d47a2e60be0ed03ee116714495e2e16865c73fd41c4f42a903cd6e63ed9e869b7da89be6f9127e952fd40ab723e014;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d54b03e8744178f22569acc2c9041407938087bd7048f8ce936a8846c26cca23ab055ad4ea8bad6c7e36bf92293c04c27193a03d79df1860940bb50c8c33b222830aa0f19d9a5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b3deab339eead2c0760ac05af887d84c311327e237c268330008a2da28f122ac70ff3a14a70b368cc4c12a462adda585c0f5100a73ad8954002ec82738d8a5028f1e8251281cc5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba9999868198044622aa001f1529f44185051d4513e2cef8ddd17733fee9925b8aac7cd27db8e4c8e68d82b3ad800ea0f8a75fb1bfe2c92e0689d0ba4b366220e8be129981491d44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8c183dba9236909773208a47de941f0cf94e2178ef35360038d3d88ce92a606efb6f2423dee414bb5c49e8732570878d27ac87e4c005d37635c15fd5004891ec52fa50e2131484d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19965c4204d0a747c286f6bba4835dd2c93cca01012bd9869c180acf92bdca4707b32146ea02b01839bfa7b6fa5abe6fc9bfe1c4cbe4840315dca29c76eb0d7ace648e24ec1bbf58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92c461ee10fa3e6674832bbc35d6a2ced31b14674bf6b9b9bf2953c367c1f203b296ceebb6f89f0d4d543e6cb7ceb4f81fd718b5bdfb56fd67a9db69383436f6f0c503367c87a4d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha880b5796089e8f8e44743cd4f4b8903c43f06ba04f7a268c5a50f7e6c16cf77b704ce677bcc9144a19f62f52b98245c35dea628e566710069a67658fc58f0f9f9fcb96485013afc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7374799ac0f56999b2653d4d2a5fb571466d63e7242086d14b49a06333b52afcbf4503713ba72a2d4e191508aa248569a8495cf165cfa5803e37f8f929db25548986fd6491c9f265;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h810c51435e5d80bc07390fb8b1cca91e7bf1ca093713241a9a71d2263b7c3133a2288790cb2b14502e2f969490ebb18e8a90917dafa6dca2af50f9794df6fbb57a923cec7b367b55;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he08389dddde5d16321059a9d532b5b1944a109770edc41cfc0a8fa171a5faee33c2d46247689585620d0f3d5f0e5bb46a48c88e70b67237a4e61fc9b96bd102b1d15848a9898c09f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88b5ec8aeea35a50faccf0006f9a6b4febf44d820afd7b19849ff73a16b414c28535156cd299cfc7a332354d1492bf4ba4486d0be2526fbcde62492077a0019da52bf8a6cf4f22c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h972f0464a373bd4b32dbece9fd80905342867468e5b53e675749d38b733981acc02e4e937151a278f1e39841cba0d376b200578885cc418034954b4b6f20827c42bb24fdc12ab998;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8506c74f661d84208ebcbfc7ab3684f6522e1a79240f942049c18f9e6fcc06471551e8b65015e63d23a927a13c1c037a558d5e88fb8d825eb89bdce8f016fe4d48835583f8073a45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b4c258a69778839deb79047bbe8040bfceb3711fa00dc076764c0042bd3603ab6121093f1adb6063927293e8ed6ebb3cc80c25daea621f5f2acb6662d93222908ee34fc50e4f281;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20e6e556812b014c9eda6f59847b3d474231858d29c685ce939f6bd4c2bcd9213e646905a642be6ee5a8edb1d17a299b1f3fe5a40ca94b3c78b55a08e7ee59dfbe46b2a812352907;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c25a36b392ee52932e5e8575bacf4f0dd8e2fe8146ce9a3ccda2c05d5185c55f390120a7e0808b5d496024adbd0ac72f8b36f2234a1236948a9b4a9451482c60b687f4e2edd0f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f947af6e5dedb2437fe1c518b7eb7332bb09e9ffa2c26f4ed33c79ff0f993d46933897ce16df3dbc492592507f14a49cf7979ed4bb775051a80a4ed36fd6193f98e4b2bb6de05a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha85833216e8f2e5bd912626faf0b8689cc848a40702f0e3082651e4dea0fae52d9c516f4ba59768117041e4f6359b111d28eefd91d17e26b8d5165c9eecb06d645fb39b645d26158;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1a767cbfda54b6eef107a47716cdb02752e6aa4a4e464794f3ccf0a9389be29f47f70a6016061705beda1433c612098eb502b403fc83861ab2d29677fefd08dbd9ce47152f6a4e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40f7bc9add53da46a9830ef544ee0baf7cc76d654bf8487fbd7e3fe8796345ab4a50597e8b0d1dec0de41bc88a601eafbeddb600356c9a6f51e512ad5a03f32a7cedaeec909a5a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde22b52860995716f36112a16f8305b39ec83ff36865c2ab3a15f15abd29f140abad2d1aadd72e0cc69e217cb6b5c653544977091324e84b11c53b4bee9f0c324a3f79cf364131bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1727526d8cff6ba74c7a0607aced9e36d0e0daa2b72a9e4d8da57804d6581fb340bfb048ab688b0140dfe5cc7a71b77ce1158094d95fc463a8e8ab04088f6a7d93ea2c9a902277cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf51c2e38d3ee1a5fa81564067167c3ee7a203a143ccb9d7d6c7d23ab73164db652b633c33db2d51e2d74f34353711eaaf3dc3d9c28649e7bf54e60a4b69496b8e0f011c2c25c1402;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa5b6b23f617fdb3d0d3c9bd8b0e34384320931d723d56b47dae33c59e9c090b8738a4239fd51d1869e0d8895f081148dce38332ce6e9464eed9eb409074f7b79e0b4f7569abaea5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9b4d15d71ed291beac0476c5e41f6441d1ab780033c09c315f0e663073ef10372d223b32502543141912b1278fca1b59becc436b92db9cfae64d9685f1655454dfe291e972085d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e215a9c376cca5e3afd05a4023edcff48f2ade52c70dfa6d2a0361a2bebedc98afb9a061d09ab94171cb2321bf702fabf84c625a9ae597b4f208f1447cdb585cbabf030e6302cb6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7ae75c083841e94bdeed562a7b5dbfa138274f7edd5529462bfa020c523ca232999a6368348e0191ec3a41c1f56bf6463f3f6689413ca2c222ce448b119fe54ce60cd69370af387;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6ad860319a712561f39288624852b251b936afe1f0bb31a2faa7d825e1b77b273ab14ebd62d56e9cde045cfacbe9dac55c0a7dc85964fa2f81a326e5cea56025502d5d33ceffeab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdecb7d70b3a5d487266cb41da9aa20246437d69ac790112ccfe814f7329f0dc2eb17f869b7fcf171e62200d0b44aee99dd99a449a5bcc96c7833c062a4646b7ab676db9fde57f053;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70c857df252bff5adf3f72639fe9325a2c4731e6c3f6253ed9f338e4e6b649102fef674f19f93ddd45cefc61114ae56c8a556d7c0515cbb3c4ffa9d13718953a9260816c74876ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57ea6a53b8519834c67707ee0001dabf9484c285c1c0cc29136a19cad36202ea3e84f7af63bc90d8ddfe0eb04d3ef5b3200de225279f9f52727e34912c8dd73dab43de62a9b2ad00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6b4c0e7b1300a889a588503cc4d5e7c53462f3b37466c14d0a20093f3ccb0c9be89a0e787fe14e7de03a1a84b843cd0fde396bca718fd7400ade9022f7aa68dfaf66081646a57b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48eeeda6decc5fac22ddf480311c71df5bf4b84fcf137607b82791b32e551516292074f86e14e763142582fce9a4ff2721360a1170a200ed64dd1dc98ffaeda93a730ef84afeddfe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3e9cb628b62b6179dc71dead7204e630a7d2f9d56c8d4df880be31d8c22751afa06c43b95edd817ac764508081b4b0e886e18dfad9e5564b2356b01c41e07aa5966eb4da86e2f3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a30e3eb9637f9f8463da49494498e1b28a95a6ed29032740a2d092f6a9508f070aa037830d3a1ac0f1d7c07ccf98cba09b295fa5b15b0926554318dc41046e005066fff1243a3d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47ea26b2c69c0883ba08f55b5f0da3632e73b23008eb3da9f6d947fd9b6d059bb9e4c482e36ef82cf2ac3285b90a15cdfd32f67de6b2a59fb282d614e2ed767f23a6987dcbfcfaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8391ffbd837f30981382d6462e12547a33e1b7ac8fc7c3db92d30b44ad7fafe62e662f2d5c45dac926d0ea03c104215de0c80311494e0d4706afca511f2536678a6027844b811a70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1391f3ef51d273a3ac18120c0fb97898a9c76b922d79c6f9b0577315c2808126675ac7341f66465c761d21620e07a82833fdb9bcd2a2b2dcd7105c011a381759d5b0b774926648e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7836958657226434b55336d3433957f6661230ccdba05ef2afe9853a5ce8b9b60c1350ff04a287778a0df21a3ed70b4c4e40fdc82859326ab8a02ec02ea87b07fd5f56ac1d5c9e1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1baec1542be1bf912d4728fbbbdcce05d735fae60ac2e7c63ec0473760ec8ea9c8eb2215f15bd3a2645b12fd2d81c4941c16940b5fe2a52509b165ec3d7d3684014aac72de9cbd43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a7017ce4e60bb3f0e8399cbd6523b61399a6385c8b34077cb6f3b79d648375cd6db9b90358048fe3cf351ea2c665b43453a025cf382b3221ba278cafa06eb133cd0b03936433e24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5fe5e7a79d3c8855ab66f4959139de5fb64e44491a6e270d280720c066f629fd0908031bd922d39917bbd2110a6eb0c478912ddf3dea2c3325b0b1ac6caee8541a05eb02ea37144;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddd704e8bd1f5d96d8d20430e3bc53898cc9f263c374e99b8062236a7fb8105c18c719fb66c6f71db1576290692fc67b54e52ca02d9c08a50496e7c43b3c3c55cc66655c6ea520b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcea41f97c0a9585bb417af3099308f2636e43650d717504d0b3711b62883f71c4d0321cd45039eb4e40731ad72331843fc59a004a6ad8f68472876d24e13fe1282a60d2c64d653e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdf493928d630c38790dae8298489484331d6bea9917708ad93c68e14fb82ba3b2e2bcab84368c64bf69ddd5f4a5e0c83f99054cae0194959f3d90aa80c41d4790231a6a3105d22b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85d26316531a83eebd6a503f5f9d7a2a6afdd7acb7310584c6c13f76a30010517592cbb319cb596b6811c07155b4a1c8fba4f2aa08a5c3ead8cc0d6532014fda5cc4114a6955eafa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6287ce7dc0be9a151e7a80b8626f42af3986bc0a7ac9456d9c3c1eba58bf1e7096cf30daa6501933116c085d5cb838317c66e45c6504babddf0667346262d88da847f2c79e541b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h334c6338a424b293588a2ce632d7d526afa83804025c722a1b04a5007ec908429c5aee07964476aa85cedbde53f6c75df83bcf1f74a954c7880a190ebbb489947c2b14de78cc4dd0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he62aa3343106ce7a3bba36e939f5fc98524c9e5dc23e50b0c7437ce4cc0bcb1266839c1993dd5d936b17d9c8ff7996292e0cac22484a9c581b85142b6247323f6d63c791412ac1ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b433b46f718bf37aaa42a58b448e3d14d07d6430982631429f8fb48a1fc4307906cd3cdecbb34183e05e860b28b1c7d0a0377af0830617da115da7785b00d3ef22e2827d261cce0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2443a46c1dcaea21ab89e87d7727184b4bcf513a6107214b0c9e8434f1b93d8f142b33ca2861fba46f45f8e9eaa90454e04fabf276c1403c60b31acb74ac691a53e03f0d259f359c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf692f726dcc2bad7c6059814bd4ee8e1aa478d796e544d4b8c108559df1fa0e3b238451a1e38acd503510361e25e76ba76132e61cf119c41e9d629b30b9f7b51aad799d504e7945;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf16d95ae95ee127d700b169fa17662f90c14ab6eb62f8647c09b1abdcddf1193e976363aad0c577e97a320fd765123ee254869f916b14d6a709206d2ecbdc5079bf8206991d12dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf69542cd89b10b77d3a503a54de68889fdda3f16364d4a7d6e8164831c135aa98b4eca6e6c99d78bb6ebce5374a8999dc6c8da854d5664caaf6bf78f6449c08b91b30b9cfafceb4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88f476f5d93b3a3478644409921924f775c163e83cc915251fbbd62f773a60610b51953192feef0df07ff81f1ecabf4b93585ebadd78ce87d41984b8ca76d41a2b44865e55d896b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bef5d958908394c0d547dff11620099d9b31392507c34a85dbdb92245f672145abed8584f80b5e0d1b6398b1b52e0592d4845a08f203acebbceec531302fcf1e3988c727e62f2c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7fd3012e60e5b7d34cf2d85274bf2c8e5b26c83d2c712bdf253a33c8b297ed9d0f6a1f205159d660e5e3ede2a7a0911701c745dee66eebf038e609cdaf90c141e7856ed43dfb49b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71a0f5e17d44ec3d6e978a84021727488b8f43b8c89ec9783af3a86ce5b9576fac200a6955d0060c37839c27dc9237bc7b2ce629313c623ee13e44037738f8bc016f91d8d7d91d1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96ec1589a5e0e08b3aa451af3ecfb49771f4dfb7f8ba0d3ba4d91e7f5a87a2321b7d7b8935953907510ac299892f1afda5ebd00e25662555ec6a44348779c195aa9ab04dbda48461;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8c14981acd1978e49ab984f917961518451342f6e1a1abf57e213f715a0ec74d319f2523c9c73b2232118f6c08d1af7a43e76f0c8ba36715cb418eed8762e0f2eca383fe15ac03d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h559d4eb32626778d86397eca926bd14ab13fbe7824e1a470fe3ab52b9593e33d345bcc53c087e5bf2af34e61fa49b622adae85f010bf6407c946f3ec71ddf773231d09d2429a9b7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd0ead6fa9cfed9013d206fbef184ba7c7b78d747fd73bdd9b4d1480b190026d8b831efe6b7f3372b659ae34046962046c9c349581aeca3aaf34c45b1ed025148c7b9b8c3848062d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d0e04adc9131e7b93f9e00f22652b9cb5c21b0512c3b7ef0a512d6eacdfab704adce820e9b87a33b0be40fb8003d587a55af728109fd79f665cb4f03b86d67c25ba8c960112506a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea476b7305cb3362f4627b3873968d1e842a96ed6f438543426ce76c78978aae208880c8cbc87a458929f467a3045bd999cdd10ea91a8f9dbd6553bd8aa5cf266c3382440c469eaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30f020ca3791fb089c2468560a987b23a47f90f5b39ecc5b00791e2dc87d8836f9f636f2d147a0a14b8a084d4639aef3fa4bad0285f1b54c86dd335a52c0c50c2c8179758bab14e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he45e9ec20eb59b82fb0193d28415160a1213d09516b8ef29c14c2f24cd64ac198cb53280f8f9a23f891f1785025a21b5d833db3b4c85af08781a461cb01152fabb57871f826a928e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb68f981a3662c8f9ffa6e88852c90c4ca6f8347170766a9344771c0daed410437bf00ac0edd92a1e1b138365df76933672c1be7b2057fed7621a38aef5f029e10d7ce65662eb0b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36bac770566d14f18073c57fdca2f71971a1896783cf2a50b4efbdb0c94e8d8d0d7964a9351e0494c6b10fa82dd762e93c8c090f86536abd2f0a3e65d5bd7de95fdbe76259d240c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43c1b066dab23cda7bc3e7f05709b79b03a9bc2369b5dbda8c8c8e33d031919a8ab92da5587e0995cf35feddcee39761acc3cc3d3c4ac4708aebdd92010dacf27e99cbffcf4be031;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea79f2d5e44802f7e789cfa23b2a2b3f150ba5c5e39d4de1fcc7be31a3d06e7341d13a98ea0cfaf93f1be878910e5f88f4b1c5aee598a61be1e1bcf65714ac66415cfd8b1f6c146e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22f469f70bf4326730420b1451b13c950b5d2eea1c33815317cbd1753e8d7c819303f3c184b4e599d751773e59a9ff99f8accad0f9f7ee21baa66e538b214156e4ed8b3129372a43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ecc88e7a4012a9735ec95a3b8fb9bc960048e3d6aca25d09827a12fc38176f13e760f4fc882779f643a60a063dc1be82b19d0410b5c267d67dd9ddf7374a5287cfe4b946a8b418b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b8780aa499fd5690d65174607deaf1af2af127027e0ed62398e2227aa89843d212222a440c54f90d2e8921fe851fbf9f1b02f4b294eb8f1f355bf09c061fd8dc00179b4c5c0697d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hded7e80c0398d9fabc06586dc1903c574d218c63c952b799d630779f7bec629d19e665e6ffad024f6fb76ee993a215398627e2554fbc25698f7e6e9140b12834685a24d9f9e256b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7715194a1a8b66fa13b7669910a6096de9cb7291abe1375471119c12b14fb08f9c555ea76e125ad44144399c31f783ec8347fa2aa8f2eedaaab7f35c2e2ac666fb9e4ef85f50247b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb3dfab967919459629971a425439f731f7eac3412abfa822f2b41aa49c0079086b41817441b61c7299023d20e48a1960ec13a05e602e7bc771d79e279c2e04ee0e82545487df0e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b78935223fc68227465cbd22fed3b688fd174f2a47fd0d858c2a355b3d59743d170b525af3e28297080b32cd8d9c7c8a5026ed38b96992ab7924fe70965691a52027946a11512ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h310c9f18e0b9ccc151630051e078e059790737c1662eb348829919ea97f65c6423ae4e80fc724542777e0da0e8ddd0987b74fa55dbc47b7194aa4fe85aa78c2348c17ceb19c8ec7a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86fceebd22afe42e0324a1ef815387ee3d14e66c24fb1d3a4da52e7cf6077d943e376dca3f5c715563c837a267d68596b2402e4863266e839aa68958a2ced992bc6bed3e6bddbffb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8d396a63ce492499cc2600aea63b823a238b7a802adb1030fa4d0d9f3da789772f5bcf1d4708c5bf2a25bd06e4a86fb34c21d2c81ff14bb5981b75597a401ab760303036fe1adf5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6323539a18392a85044e2f39cee284f820a6fd62b1cb3ba9f3c08053a345972f390308a1da91207585051be0739a11388a03355c0dcb1e4d8272cff2c69f7e6ddfaf97c824e4a04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c6286d35ea3620ec0abfa10f2621996688057727a63380333d9319d2e025eeff185aff887a91705f4e0d18191963aec8666e0ce1f5b00bb178e6854ff49c765a2129e316be72b8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h168e7a8d59f9461542933e4d586a44b5f5fc14caa5c816e7ab5655975ace3534feec500a58f2e26589f1b673bf5ea327510ef7335e08e16ad5fca7a5975e58f8d466aa5234668cf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4b200e7ddc7f3a00b8e5bb497a95e046ea99ddfb5109004b13054acf964856366566b21ef393c2fb28858de3d218d804664082469a6d2860a486685b0b4734801ae2bbc1233fca9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2067a1545728cf7cc554c7a7278291e50f04a5f1d151a60b8f51a266aab2e3221f825803db32dcc863b35c863ae0ef2493e4b6dd683a3ea1473c5f253a7adf5f84fdc90a1a9d38e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habb6fe0bd30c00ef33398699d3bf8d1b275a4b7e25bdf721470154ad053b04547dd410f07cda8a14755387f96a529cbda3d0825b7a5d6398295a1affb99080e54c9edfba0688babf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc0746f4253da4032d31c1e72549b4b1ec664f403b350233888a7166db6124c3d13d6f5bc0a7f3a49932fffcbf581f2691a5799ca19911b7acce6251a35bff76373067b6171331b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2e37c550e06563b5e8b4684364b6a4a56200455276e4e7d4acd8d719fa0e1a2720af52944567f776ee93e5dfac36b442aa515ac45b7a76760ee517c26da0ccc6b9a5bdfba67dec6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43f1285e869dbb49fd492e8c3f738441dea413649bc8203060f52dc0035c3be91e6bbe07573e2fb857c9ca6cf822d57d5de99d1a881dbba89e16492a9e82782dde35712070479f2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc92dccfb8c6dfcd4e3e3759e49038653496777e897605bd57e55932b6c050f126e7c8ad33185ae54950d1ee5a78bfffa7a91c652139329f41a3a5b921f4a55792ced05a2fe99cff8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd657be2b0e689b80b7a49ef504af952d41241bcc264dbad70f57bbb252041835367b9f6e3cb5b1546594ad69a7d2f523b65cd945f34b150a9220779dd24dadc38ec8ad2ac97948f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb4636e94bab0d858f12d672b8cf117b4a65d012e7a9f53fa8c98a0b4636087ac12913fae27bd8f53f4e35059f62b707027f146b03f1b8141091efaabeb7395058b08edbcfa609fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53c9207427ab1c7f0e5fd1a252ea58ecb867ef0b164ccf677524c5541651b02571d4639356854121809414b46cf8cd86c78b141338841dd61b7ea3918fc7a699f863c7a97e198b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b8cb58e19a8915dd631f4a48ef12dfd6c16a6ec9e309e08382562532e6d55cc9f45e1f8d7aff6454866efc062ed458b98cce86640180d1b77ae5a7bf51d531177a066988622e9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19f2cf1eb5efb674c44bdef87d64a54143e7809f39fef39b4396103ab192da954da87cda7949561ad1ab63bd98d9de64b66184f35da98c43297ef4f2fa5a35484bd3d43ab63a69f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5731da4c9a1c9a9d4f922068e76e24b5c16e4c6c7e62999ee849ee5b7d951b71ac34cbdef53e3cebee55814fe7487af8d0032ca4007ff046b0f134d3b7078c4a3ef00f538bb2bffc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf23ce2febaa7c5d075ff20c86d7b52942e2d0443d8c2368a988c741d6e8f775cee01be8d1ac43fe187cb6cae273a44a20b31d3112a55a3e6ea9c4d419eba5b64c02aa243ea5c0e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h347d9e1129767fbd85bec221f096f858e0b062a51c8c3711cfb1b1b30c723e175ee802c08392138309a8e3250c27be1c746df70c6f9183f74e62be569a6c143e56f915190478188c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd5fe1ef6650e6779d722ab05f9c1f2935077dd749ddb3020806a15fc7a23ad387608d6023a47ae90d843d4cef6e0aad4fd34461b32aa02ae8c03c5a372e3ab10926dea8283bd0f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59ce72464d3c9ea367bc4de7418304c9789f9c248a5e3cfd70c8e6e9216f19736c2749f1d300a3be3d80cc08e56505a047bc3416cee86918b1d3c9ec06fd103c1143a80a7193b20e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8119d3a0a7dd1a48708cb65899a6aa65e3f1402a2ee4565afc877ddaabf10c813c070625a82e5c61679175bb58fcc1e9b86f13a7a45c1a6d42701f3341a7267f6addc1c919d64db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha448af0e9fdbe24a92b204d964ce160f1e3741dc0117a69bb47893057cb56a111238cb12d65baf5e949f88e99d327023332b44d56b146609c4688f832be78dbeb89a4b5249a3fa86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3f2f10e03c6941c41e9ed56781d9b9c8ff1aa4278a5a5903fa117230815447c82fcb447bf6c52edd591a17af812719b593bbb7d34c997deb459c1ad0365ec98e284b821251755f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60ad2ebd32a8579b3d9d07cd3978711c75736835cd0269d537ad3ccb9c0a966f749ef86468889adc335320d14035a65b616bd1a02c57a0140c29f1aec8f0329290d0c2c567ff0cc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bf554b09f094653c11e7f48758cf1733ffb5cfc95e8b79a703352f8c31e7efc6ab2e892215ddafddbc23553264768d30f076bff17cd01423e83ada2210701553482e94d5f7b8260;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7093e38afad635d2d83de465b522bc737a06f6838c3dfffbc9ff2ead5f55d03cee351de230e97aa2de89a3ded6fe03062e7f92e0646b28184f912d52e67e388e62424cd64698eeb7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27c3ee9464fa03666600539a5e5039910ceb041a5139a468d6c4517dd99547da77405c20166cec649d0341d4f7f41441790561bf43f6901708db8358f883085f636528e4c7e765b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbb1762591c8f9c2b025dd955acb3ce78b97988c399ec5dc579ed2439abb3d53be78e06f5bac46301af12f7b482051966b4643d514fad2df09a04ae8f4a91181ca26f46f92ebaf24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf2e35a5b9fdd1ce89a8f5e7961927c8ed265b69313b1f6c524a0a87d6ca7394bd76220cead786fa9db9bb6988686fea5d6cf494b5e83d2726e85126cc8356dc9b3546ba1af057b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9daa41ac2e99bea521d91d02bccb9cc637f07c7a85f5017d12c0334edfbdf8395fa51f382a7b1b8102567830e7994653abdd651788e0ea4f2367fd12afbc4aa2915b543d3ad1f48;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43ac999b8bf1697a128ae1ce6afb7bde0c6a3b124d2ed5d203d9a4668a01d11ca7a9b37d7fa10f42dd4f5f9a503b259c66882f33699cfd9211c7ad108de0336ca92511df15f02ef8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h168ba1598ede1b4b1d202d635ca5072e265549e5e88f2f0aa9bf616c2a2b593e33e12cb535c4393cb11942b56ab62fc4eb4829c5e7d5dc32855adaeba266d1a2ba1db688a47b2175;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17eac29d069058facfff1d1e6040f7fef84fd69d8eeac68cc333bae36d60311248ee0d29a40b4785ac046931da8653d21e10c8e1ec9f5b9ecd453b57fa2cc10ec4a5abe155a16066;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f3ad3be72a38384c0580f7f56e8f4b4cc9bd5c3fb997c8816087db42245a528b93c46e4dbd86da896cd187e9a1aa8f0d3d4b6f7479ebdee0c23d76d9f89bc2b25cdce99a6899729;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he63e9831955d614a46ae2f079a7e72d7732ecf2c19f1fac0c520bad59a82df2ec13e65700ea753c98795731ac64e4778050844e81e78723621e036ab69a8f79e13db8998b17bdf8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd212f848f12472a33cac6efdf299f0928554addc3e9c4e181807ca956c90ef0ddf152df53667818e50e588971353fed4b1c69a98194719256b91ab81f3019750de7a336434200044;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8638bd9e7166dd93faaba7a314648714f5dfa91f6f8bb1f48291722efcb39608134791e0bb6070329a1ef757e0bc7ae67259fd0f985f51067e88e9b8343ea8384d608f76943b70e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf78251a9ee65efe8f924abe937cf7b1a111768dc990a26288cec5030be7c4078325ad67454bbf2da9499acd3852340d8239835f6750e2d0350f2e70be3adcde23cc32def50604c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f523275ed74dd97ade3ad0998e2e917f4f3d17007ac90e0e204d4a2c4aee05a2b0f36551f5d00e45c503d66e2d674a834ff78c285103b7daebc9da7d13a327470907a54dcae5fdd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h802a317a092f7025ec3a1501c68bc370c98ce5f85db3b49f09536a8ec249cda88c98b9cf74153651c2377f6f55c25a9bcd60f9c4fcd917506d63110d12ea1ad46d8cdced68d2bad2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf368c38895411ad1df35d48fd8b1a5864fc22c3adb74a4e2524d44fa3cceeb8f85b31a161c97af59be71af6c10bea26f717ebd9c5486f83de4d52e960097f05d194ca69343ddfd10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ece971699e486c85042af2e8db0b97cdc051a8988119bbfa35951e35487160870b2fade11a3d5e38f3452381da805560cf08e56ad6a203b869122f4a4424dbfdf15e96e91fcaf86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1630996e2e17ebabc684532efcaab8fc55e0b313a1737c80304f670b4fb5d9f8bd29371f69c1b3ef3bc3dca318259f10e455c1e860f61e9b612ff777cb962f74ef9dcef0f71f115f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb93d27df189aa585db8942769197620c5ec135c70dc0991c45f42a17d7703bcda03d374ba2dee8b1a0633895cdae5cbd36dac823fbcc206b08d37a0db613c3b397709b2000170004;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h783737450cf277412fe856e3e40ea44e7105918952e5170ef56727951d40294a8bc1e2703981d69c6068eb54679a5b47af44ccb45d90417e89a50b6dbfb6dc2fdccfdbd3564519e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94b7945ba84b1964725de4b4d4c94dcc34491ee7b191c099711ad7ed8ef729b2cef17871c6c51dcf5d6a67efaa27d8a6354eba2583f752aa6eb28ad720781202b684513a8bb4fe6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h866744f10c892c4301d2bb8ea9a1d529e8ffed6c8421d3b6dbd0f0833d68593f43ff458a5918fd12176fca193ae6af0e6ad83aa14a1113d9528d50bd0bf6a54abdfc3db36b94b5e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1594f7cbfeb8fc41b2cf845a9f9b84536f7b42303ce59129add4b848a71cc055f9840558cae7155ad18e1aeb1a1f88a8c31a955b94f792f9a6cdcd118314ac24863ab04f1ef4e478;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f21e4a4badd4a1e774b5c7795693226f9713ef581b207afdb97001b1ddc58308d8c22fa619cbd32df952d4c203ce02b31fe7b297e2d9ef7fe1b3d2cf5c090389b8fea8dc23bcc1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1a96d0dafd7da10948dbf122e7cc7f6d3e0ca24b9f316efee0c52b0b452508d1cd2c4a974da911589a4ccaed5cfdb1ab2f298bd76e3cc7b70971e0b3c534072089a85a5137d4b10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h955384425dfc2012d0161549d9e2f364e6ca97cd5062b1213524a1733eccdbb4053e3f6d08551b4688d637f403e10d32a763d41828117fa1f67397bb039b8e23eb684bf1a764c5f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf082c9d34b4591c2d5a7da0d4f19616f1253a3f6a6453aa37389b970520e55925e21b95d07f71dbd1411c0a976fd2082a3ced54cc298548df4496dc73140a2e7c1bd8bfafd65faa5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7b67a0c43aaecbd929b31e79467ed29c8db5dd688f81c16956d9d31da70d9440d13171a4da261154efc586e6588269a2903ce7b5d4f0970e9f0b4d3ef9a8bde28b4bfd399ca40f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce7cb987176030772d501c9b1fbaef1dc6e5a96885a67f0205350f19351a7cd536c85f2682cf6e175802cf87c4fe6de5771e73d3906885f8fd1231f6608c6538327bd6ffa3bd22df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha57156762ad04cc8928a219397522ef7c720dffd0740702fca8836bad2bbec8841487e797af94443eb7bb3f94c34599259610fe61618e431fb3db712fd84d666667b4233c00ba7ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc264c8602cf4b302196102fca429757bf38ee791fcac212b5491d77da04d21c65b331355f3b124ddc258026fd527cf90fc7b2c1f9f75927e8b0699a8f878a0be23205317fb9bead7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fa022f55b0781bf03b5f455971a7107ceafb97c0f781c809927565228b2e953531ea7d6b72e8f54e86245b625069f2f8fb06f9759a1d3087c3dd8490420079b544c9ee72cfeace9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7ec2ac44dd2839ad3cfc94795724b46b45437db02dce9fc8c25cd7355342eb357237b0af7c04a89f56e0e893b9d944dd9d4bcaa8faeeb2b3dca13abc84892df4d0ff0b6d9e74259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29ee13cd9b40f592fff42f43e6dc65df3882d6bbc767c7c5242cd7ea85852be80d5ccc414dfecbd035387e8b8a03ae10ca4231a3643c26a759430dc98ff2a4cb5baec6e233dfab1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16eb6991016fade7e0310ac848570b8ccefd5c4011c4a348201aae4c15fb2937654f389a9c331cdce485673e4d85dd70ca8b8dfc78169d5b09f054ced0d05a6d78e63f30c0a95cc2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c66cd47235750da6a9b8c0ecadb4e56f1e0b35cb5feed2c0ea05d31c17388f38709c62461f31e7da667a52301db789e1096464c7ebbfa2d823ebca55c3cea7dca185bb9a49c28d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h872cb9cdf4e9c6c29a31689426c7eeed1eb48adb48931c781ff0f6a008b67e983f41c235f07be80377a5a4ce74b67c1095e6e18fb4748fadccb88dafcd3d0b7f4e28e5341e022a1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7313d7742223e1ac7fb267f7b21b0082cf2db58d809e499ca92daa5bcfe7731911daf60dac5aa646f1fc5fb686e9a89e5611a5edca6aaa0df33082d5ae24a088013ee62e777c435;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78bc712ef553079b880ea8c10050649e0b173bb02a13e0ef7d421b0d3a386a3e85ed2e0d0d20c5f6864ae1d2451e009dd3e806b213163fefa821a8dab4425b7dd659ef9e1288214d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc391511d498b4ef0e9f9e0be34d27bf359c902f19648cdb303f25e04e8f4b8e1b7b7712406938c699e450ada366539f497c471470953630f88fd68b6eb28dea01a8c5b996875627b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8af8bc33e1f1f825372b183697dcbb97c69cd7e1aab5f11c393a42c505df1d9e8b215eafe5cd1a5a717e0e5ae27c889bebc3c17500ac8fbeac20743908260525b2886931f1d9faac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea8ec126681d5ef3c3bb34f7ac5edcc3daec487b0de2b9a96d580d1a69962aaec7802b9c3813008d2011201a0b95145b938f418089d3459853ec1c47da29855bdaeb277ec12ea5e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e7296df60d0f898b6ceec58933472b91e68fc7fa28236cc621e78d2c25c6afd78077711445dc11a8b6961daa6dc59f5c6684a5ed32d172eedd415fa87b2c290332144b0db23d277;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bc0c0bf7c491883cff01e5171f3128e18757e22811336a8259f0874f545528fd7eea7d8f120e3716a5bfffca2b6594245256021bbb8e833cca1e61788037e3cee13ce0f5df93317;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f52e1afa06e181aa62e8beb274904bf2b117fd18952b3d11bd070fa5bcc4d0f1f3e78c4b77456e52dd565b1e9c39dde187ddd9b50d882a620fb6863ded3a597bb48d18f048e9cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34a17efae4fe09578ed59d76bba5755e67873cbdcff896b9ba9a0cdc5f728035c491cb315ce7df956c5520b227c42f9cefa2559bfe3b79a8c1af04c827356c5aaeca6865a4334c8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4ece7ad272485054503a779ba94f519cd39dc8230b45a171f5f5a223c065af0578a95c48e0cbf516ccfc085df6e95ee252785914a3a6a932de36ebb183df64ac36d8b28a877cc0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h612fd6d11fad4718ec14759e7b17f294ca30b35e3f23f03cc70e6273c11ed6a7564bcd1439f5e2c226db82779e7c3a0e2014f6f4b68fc92b338215a1970f9a8c9f78f7a23bd56ed4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb456ef9fb290be8e6758da092b65ad550fb4e1f9e6a5a77be661eb70309ba144f789b191492d4c14aa9969abe8dd6667e46495e0ed778314abaea6bd5fa7c4272f51765594f370b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f7102b5e38db3a2a9f0e66d72c5b29f1cbb2b24ff22ac4bd16ec54d0d07a6fb5f64e074e2ae0410da09b879e97be12c4ad6cf659b5ca2b731399a745b18a9810eb2089d41927c1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1444ba2d785775e1b7bb82e431eb356e5360b112ff75cfc04b449db1c5dc625d1442e5bde96b5c8fabb5686972e184fc8d840910706d8eb13558b7925be4c142e151128d47cff80e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bc18a1eb1181bf366c6f57f4803ed2322ed31246c64cb064930bf6c74570f218e7b8d32ea8a206f67df4e60922423b2b297a1bd92a87525efd5cc65a053e2b08867bc4f8b06f2c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5d7893cff6594d88a5ca58960b94a701d9276f86a74014ef48fa5cdaf2cf26ab18e9bfce9b327f50c7c9bb47e71ee2788d56c09fa907912b898bc8d86c1a22bfd48b3b0dee86dc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef02bdd4815c765ea7366af0ff03d755188abbc723aa5b6ef059b5aa97e1467b2f728a67742cf371f1e1511e58ebf20aa566b6b3b68d5e5690ac27bccec9c1e72c1914c78ee7b259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac8d9f043bbf9410d633cd0382090da98103d5df6ed6ac3245d539edfd658c2264abf1687f8418e8a736740d8fe878156a9949b419766be360607091b908fb587bf9c44ebc37ca26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42d280203121988e04f93977940137818c8982fca38dd99c5ae490e18005dc869c7eba47041ba6cc3939907c9bce8224965a02603214e9ba23cc2f0acd190115ccd2bb74f6776a1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b51dffbed710791b54833a3b7a04e6bc85cf9670de794fe63a0ac4c45b51b3cadced6dd5de3f365fa0e357348157277020dc83e005e3f371f93a4b240d7ca558e546b5c75ab4131;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f3687e33c6f855414f62f5d7fe2ebfc22799bf8f082b349f158a07fa11aa2cf041d02edeca6d6411522570095c84c71537b74b942b7f491417e309c3b83f3f3ad548037cae9c02a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61b208517b9c8ef797226d901aa58694f80a21b69449888ff7b9605d3c5c62a97e78a9f92be6b9e850af5b9d6acf3f87f8ad2ce51dcbd829952acaaff04bd60ad4e58df32cc84e86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3b50e8992c7bf211d23feab71420f8a5a7b9ebe1bd5d5ad78280353065b8ecbbb4e6a5c498dde5210c5ddb8fa72d962873cefb0d20067b665cb94b6476d65d2519e71582c1d2c55;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c1fd6e03dae342886f9a94ce7ac7e11c70ec7c242ddaca1da45830319edb20141229cff27c8d3c16af30d1b8bb95fa6a731002d1b55b481f861542aef99e4ea0dda2b7a75ce4cf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h243d67a31538337e9de6fb60908878250eb33465e2db1769ff6146755e7d49de80c14b99780b9f12141278fd8abaeedfd1b945e752de8f4f7a586f0a2c66615213004fa286048dee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0cc6d34cef3adea5895c920f7ffb5afffa16df7825be923ebb308d2c18b9ffd5abcedf8904a9b74a3b535a8d7fdb70e8ac83fb5f8ed6aab4ada540fdfbb0002f45903234a084e90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44d91f634f96f50b432b33dffd7ea33910325de818b3cd1801a70807f19e16572128130ebbc3c79424ccd4a4fbd867d15717fe37defa7a674e441bf96c61a98aff9d976eb5fa870f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9124821a2cf9adfdd470252ae6f05292c4b25f6ec91ff03ce39933c5546ff88667c4a8cfd0bf62856fcf0802e5d59793566b96ca2209a89330402cb9f7926c08e8e4220759b52448;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ebec695b2152f8ab2a1483de6e8ebd81bf7c1ed3821fa52e07732f27d7fe20b11fdbaecb0a04d09d5c08a38b1042b777365c2bde9717f9dcaa40c1b12c2e05bb02c62f72263defb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h773bb95e695cdf43b61a2a0b5beb197348221b8536ba0325a286067567ea90d37bd7d17af4f3d28e3a8d7f891ca7e78e219d9231ae34e3185aa601fd880c4bc046507fae0bd4a118;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3fa8cb3a70a26aa7c102cee0efec403dd77bd57487d1b40109a41a83be10182791e9d7d734d9f59b2525ddcb24a5cd092b044f8e35cf98032cb264965fd5f427d1e4167e1a0a57b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd474592d5133d74016f98a00413304902fe6bca0ebb42f7a079f296671f37f558e09c0569225e081c40daf4ba8c108f2cbd73f8886bbc13be124c7de5ad299371a1940799aa42e5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h642102fad8bc6074f645d02bc3861d83ba4a64b26ac2747e3481c24869b3341405a08eae8f9e987f97b5cb8287baeaaf8a024fb6be8efdc1ce1c0a3239e4d900999991d54c8a87f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c6b049d392de352d07697555f23e71277f07be069e22c6ada99d0499573a301fba5abe9157b7bff45f3f4573ea5e350bab18a8d376f97c531057d35388a2e44cecb5d137a8a1f90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9217507f1e4971bd7894e6913a0b4db2692cf35ce99be978756baf980656db907e32a24ad254e2078a7dd57da61f635933655c0d82f944f3d50c284eb2ffbb2c580973e4a7089ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52f433dffd45ffea7e025a28a79eb8ef585154d27745718495fda4a56fcf4dcf723078703160383ea34601942e5fe248d1f9ffd127a3431fec62f775f1b70a18dd992ff8b6f55413;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef4f2445c7f3127502677ccc47f1a43d9d63817e2f979d27e123bf4a4daae27c3a291d9b10a9162f34981d0a56ad7d49d9189870617b1e770248219596458496405f305584fe2290;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h345e278c222357a4015fc471923b0d96467e312d6a502ec017fd9d30ecd50c5c23e3c6d87b747098e4194d2aecc67055dbe97082c07929f16e7a89470e0c5e2860d259b00fd2d7e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e9c8ea3b0e3c48246538103c9a65f972e74882d79516cd875e960403c4ccc6a9e30248092a7fc4f5c89dfa712ec1373b3a8a57b56869ddff4fb9e2cee86f9fd53018b8f0bd14eae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc05cea12a2c5098dd121569114a9aa6447665b8d19ba7e3e561ceef5281c583ff2bfcbc9448fd9207afbe4f9ce906f2f07c1f3ddc4763eb41d442cb7561a1a4a2537b46532ff9b19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ac6d448adfa66f6aeee8b57c2851d16a2ab76619f23aaeae724a5375a70823a9821df81c10de368558ad55bbce82a4154db32532ae0a86fd0660e33a15fad9352378b1f12bb3131;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff17a35dac04be97d3d0d87b6de14e832d1750bd3fae52fbc129cb844437bed6a3d122cbadc7c7d29e821455446cc303a0b136ca52a804f06cbcb4c3cb215ea818f2a51dbfaf929f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b85d9a6cf64b4ebc241ac430fddf4aef0545f81ded12afe55124e0beb298449e724ccd63d194e9f6e9153b0d8edcdf10ab3194b65e40a32d747dc0d4dc0836fb7e3f440c4d37d14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a1d5ab8bc751c8d258b66656dfd6dd29eaf91b8f34970517cd686b702fbdae6ba7e26286a9ae2b856de810cf5445f0688ec1c9c1f965b554308a63646408662828d100f62a08bb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c179e0d780eec47481824ce85b37d1f894ef1b42c6a9598f2fc582997f2b76e00b7aadee9ce2d57a5b6372ffb60e45915cc4b4adcb100a67c210ae0b564863d8d931efb326785de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57dfdff0719203333815f1eff22d9a2024a11e87bb83d0ad8897d011a497dffcbd3f94055c9ea1a562f78adf82fb395325765d8549f1d71d7f53b76ec47eaad403bcab9c99f74ce5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h388d3013df351cfa92f5757c4a6015377173dd05067f476cc5c4242aed55d65c19d8f82f55d4f1fc359898f42a3502c9a5602127baf9de1ffabdb4faf8a6ecb9af81ef1daa618e92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha07933f7c9350396df8483d795935ffe31001dc5a751215102845e5985fec828ca8fb8f7a7abaef631a8db0e81b8564bea9b67409fa06ad84c499c3a293779ff333d448d4c608e58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h325cef0c6dc7999d65f65e9a7ef9db03a0c94b84a4527a3dbb33de21f188ffeebc0c14ca38fdbe262f5327b9b488994e8489d7932276c6c39faf37d666afac9f9e2a106fa1d3cf4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4a1209f8261af2e5876051c3084da1ac33108a514ec80cdff5446c24efea97c27b5466eac38afa7fc36636b4c8e621b36d881dee9aaa3cb3644de7e00c94a455c73bff87e190ee9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h476b9728dad7330dafd79f33d23cc3e45d9ad2020b5bce1b1f0c59f200f05e185b73d60dfe595989c7762749459a9908002448cb60f0c5b0ed31fba6dff3c64daee32ce9f7b275e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36c45eb73d6fa799a09035ccf7eecfe800c3dbf792578f02710e8e0a645755c1529af1bf0a3678548079becad3a1b95ac98c182156b70132fd40215c184f06020730dabc8c34ffce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5491807ff566a4e4a1bccf0415fe93c710570b0531c3dd18068e976adc27707543a0ae1c3c5aececf30ca520d1c502aaa3e21710140b8e7b78708eb4d72fbb31f8ad6d0999f977c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24e88a469dd646e1f732527702b2624c99a1b4436b49ee1deb9d4d7b164577c8e3d557a3fab5dad41e926bf7d26f57178746d68d711260dc9cf60333f9523bc4e492b4f14f421bd9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34f22ffa1cac8a389b7102aee6550d6223142ba2f42d747bc8ec0ac39bed6ea0dbadeff81d9f3a5a24cf973996511a4e3eca713f2b2e83905541c3062e3b1482b69d5e85dc7c315;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8307b4b8f1172be454bb996e842b95cd83d9eb1a3049f4b278d3e50d9a0dda9865b88f0e44bb84facbb7c1d1c068ca6c4532dc6c34f7f2f4797b6afbe3cde917b9395639239ba819;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h660b43af9d9d599ce3396b20d8c6df239bc180c8f156a83730f8f928e60c52b7faab4f202e81cb850a2852dc5fd5a3bdcb62b974de78979ae7310d768f25a41759a8fb003ea577b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9b1e338d856c6d6fe51242d525dac4e9ad06da36d97d9c51495923181f799ea2a7e449555cc5a257df331240e19555fb13e3aed1af7e4d0b044bd910aa77529bde06c51b4c210b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefd2f0306459942cc281311e874549b8123f9b521c7349ca72d2805df448eef5f415e24a7745097e8773455f8cb27647efe405767c8f881194a3b5f509c8e2840c35895a602c5a1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dc8ef6aa8dfb18eeefbd9988aac073294b0691c1c83f0f175a544693115373958deabd5a9a8030022d52c5b9f6eb441baeb71ac0e16e9deec2ddb6fb3b70db637e606fb2538658e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd8b551bfb14c6060b2fb7fa9df192293738686c43fb4f3b460b032dcbf1891a91aeb9421132a17e8782d73fc5c67153e88eb68a34b4fdbe95d245b04bb87957a1ec2994593a343c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb59ea52bd7256183a3f2b1831b1e46daca3cfa3e21e3aa050a49dcda246e33b888f32e2b0001260c1096b15334ac16739c189f1fad9112f3f866e6d93dc1072a825238c218f511fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc23a6aa8ef42067224794f2eb1b1bffa1f043c0a8e4010b2c720afd94514dad19497ba2d3dfd8de644d2b45c416879155251b54679f70b7f12490c3372fe8847f0f143534e2ec950;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h322086469237809e6421222936dcbd21061f2761e677b2be4355d788e39efe2a5f1e7f45991e4b0d9f7a51d51b83891934e4ba2f53c2f1cc1fa71de4e29f752c3ed7cd6c28bb7a03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6db62aaa954a3df2cafa8b27dba9fc2b09fb5f868767772224a06fc56c28407325d992fa43d5920d34171efb05e96be3bea05bb8fec66dfbeea142dad0b7d8df3166be770ba3aeb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc138e620049194898f60c70d212f9bc25f6b4657a430d97916454787b9248326b7a7131ac9de866e3a7b739acd30c280f07f3cf1571af4e7f61e7390ab3eec1e1fa6e6732f2324e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf79b447244a638073b55472a356288c85608ab4d0ee1b63f25afa19d5b2dffffecc870ab1832c80cf0021841da512c713ea2b2ac039c9622ddb00607a70ef4b9294b85572cdcc142;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4645e2d165d3761dbf4c012fc217a77c1651f012060e19479900b7da0029c0788a8a4b548e039942218dae6780c0549afb2e4815deadc5bc1483b349991fcdf1a0ceec0e0b106f46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9983a9edc03435fa800484111061cadb8db4b8b26e6d75f3f568cee0d8550c5a2606e587363bc6133775819c24291697479d5706b01df45cdef29004446294201d62ee744441b33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d5e38e3a50e979c1eb8ddf1b4690b81cd7a56682a373ebe927d21462cb7a5229abbda701b04bea17a93933044632505b51ef2c1400bc3f40160bf36d696b81d2e30345bcbeccd69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d207a4fe403985a681ebfedf97f0675aed5fbfde9f2a526bbefb1c3ad6e4d1da7dc9151a5db39bba4cb0155fc7e3d371c42fc07e1bf93fe8a97a1da74eac3b9c0e7788d83f2fde9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc57711abb841450fbb2a10d2e45631cfc73593dafc654241b671f366ee9ebed48b12402e23bf51b4dac0e9acfc9f3b6f0fb914d8bcff138dd8e8ff2ba2c54dc4c98e8057feb1f98b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha36429fb960dde86cf373dca11a1dc9e05a4dd1c03739bd27f795561e975352c372e5e0414ca71a9b271cf5cf346d3d1c9669a25325dc9aa3fb569fd539fb1c61367bfcab10d26ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf25517e4091106246afa66e603c24c92f503d68a3b05cf6431d25d9e47afe0821f0375fe05ffe4938548d1e6497aad670ea9ba83527e2eb09be5b8f7de8845ee3b53950f023b9d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddba200923300fe0b3df0640d4dedf2cb7bf5341c835eed338835982a8b0801fa5d40862c6fd33c3abe8120d84a7dd876f0e090ad563f4c70217bddc5ecc550509c414943d364c13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d909d5d8a96ee0063d7a65ab059f1229562f502cee45ce72573eaacba8fcfa2dfa3b63f5c616af26e259f43b98d7e2b20d2ebe8255de39cad69328de4851761b16a5b2cc87158d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h677738557b8a066bf50e3c25cdabb5b3ca42d8f0d9d14e163d200efe8f74b6769cb4891649c69240bf2b7d6931efac54fc887a820ecff54bd89d0b5c8ab8134d75f142373680bce7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85df28d3eaec0848836ed7b9056125bd0914a8a70b1cccb21a13d1e87e0a20cfe657e568258d02cb60fe628a803e18cf277388a25bff2e57b846a4a7945b82a34c8dd2c535663951;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10239de1e27e957bc241c61addf9f42ca35f449b194fc8e76f4be45f424ff728369d7288858326aa815e7bef95aee453a7a65e2c14cad4b6503e0922a0d526660cf6b0b61550e678;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33f11c299fc55dc89a3356d6be25037f210a1a9a4968ffcbee8228f83b1c89b4f372cd2e1d26f9661fdab4609e1add0dbfa71b48a3c1de6d63fad027b7e797f7aee591add94f075b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bacf5cc66952a298dfe56f48be2b684d98080d821585732b58d4f86b1c8c231b3ce7b4ed14947c77dd8d726c4696cb83cc100e9ecd557e240eacafca6f436f97140cacce67c3668;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dd4e5b97ae25ee84efc83ced2bae7f6e7e93a5cb1a21925e0374c143b2f2f9891fbb8e324e781b60cff16d27b0d2d61bd64d1f57737078bead3baab3c73679771752d49c29882fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3d035583e31458944f8fecd2c1a44da6c6dd6074f948641cd073d0a510f585fa60576fb2007b37a82f98da8bcd1acf5b7e1c4c69087b3f6da7906c131dec5b9f69c02ea12191a73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3975389f4ea1f8f9bdaf9522cd06c1d143677717fe7be98c08bbaadba6180b095b452a55869950c7908464ff088521bbff18b3b1ec180b3dba86801a215de106d0490ad45a08c7ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34912538c6e1e70f8e9cd802f2e13ede099318fc1458e1047d9a28ed576ecc9e07977db0253338298583cf5128683d7193fc844b449ad4aad2c4121c303585122eb0cf349031cda5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h578273a1d7979b3ae023a6db17b05160e83546c69c3ebb4fe0915586c9f004a14dd89877b5abd267bb6aa5b0d35fd7fd7097e4688a5b4d4379e9a7f6517f2b0e82374645872a51ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d015ed053ee1340ef377fb6ac508e3dcc3f23de9c6c26cd0abd24dd0ddf5569b42a5ab3d6da5cbe160b3f0f8883261e1c68af83479b123a7bfb1ca10eae2a09421a7241fb3c1dd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf65dc856ba27666355a07bb44b1b318a1cc32a83c99a5cde3f1b64ece51c2af7e4d84e71f1f9ee8950c0e022ab68306cded770ef29ae5ab5b2ee4b87e446a08a53265d32944e0f02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he794f317f894044234d6a70df472368795634a90304af71edd3b479fcb244bc7fee54e4cac179b86ef52e22aa6bf47c0ffeb6447501673b60120b1932b9f93dc1041a47f6b4aabca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6aa927308c488861d4104caba03cade13d2498fb88ef2d9056a225d748cb9ee38cf4f14a63ddcab29f418cff93eaf67864652bf1ab10bf5db15cc39fe8f018ade104251089441d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb788bbdb483f725f5ec19e60c2f5cd20770306124081a401ce2d374626beeb23d3a2d9ca0f09e9f52159e8d2ebfd060b425d4994d868911610675b80d4390a1f91c5a29824827473;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e409b20005ff26a670201aa6f6aa52e954f93f2fc1a258cec824704304c14c88756ecd0fcab79cb6d27dbc795ec1f2778c7521ea48deaf1de926e3c65fd78da20e40ad89b618bca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he06c11fd204b2490638f4a4c108f7c7ab79d1814693a7216304bafee26a9f67a9bf3e51935ff193f8653688323f022d259b1cd40ab435480d7bc57c012648450f6c0579c7a256fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h840916a9c8a8acd02a5e26e9fd4f18a74edd2b3080e7166484193a6b6ee69d032bf54a64ac1db09790f666380440733c7838912d2e537b54ebbaedca3ba642686477f5a0b5d00836;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h138f23ab3ba363a95fdab5073cd34ec2eb6fb20985f6670498b4868ed6ed7f6becfcbc82423ea4f7e644740d41d0352c55fec8fb97f6be1eab35c6f7baa24394af291d4047c21af2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8d1c80441334d691d2abac2b5478848bfe7676bc59c3c9ebd83c5e5278ad9cb180298cb85d46554eda8ae32e4825cf824f1db21a17a6414c6e632a40bd1be184e2e0b3217d5669b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23566def4556cf6585409a317dca8be4b71cf2a378a688712a385d16ad372d8efdbdd4e52f7055b8542704ede10b89587dbc7c4f95beafadab53074d9b5b2e0b11ff6ca101e9f516;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h542f01d9f9f15f564550221fd85663b8859ee3fed241441fdb9a6fcaa8dbb8d861b66f5e615ba2a798af87299ed0b6ff8ceb32ef36db7c512865fd36db9c6e1a41980a86215fe43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e978a05cf2f69d421eb79fd9b4bdf3dc5ff9342c4172b3a2770c34247babd7e26d27502ee5b7391a07146ad82bc739423e8022b7255ce02055ec50c6509002097e04b76332eaff7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87861f9cbb2d4f4d11ecab128483efabaa0fd67433e3e654abb50376c4b78fbb07d70506cf6780cfe2d6c28a67d0b4f80d11636bfd257ba99cf648998c291f425ce319117cf751c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1a7445a85dc89363e8b51ccb1d6a0ed747d8b8aa54e63d316e27a28f7510676dd5739b331257325b729dba21fad4cd790d9bd62a0d586d0e525017284cc7cd8edafc312b9569578;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29188028888770b70ed1e514d5eb47a5507b68bc026fade0de6d6fc337b38aa6855415a3cf891306b4576a23810632dfc8b27de41554e32788c884f4f8eab428b1958c706f50c4c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6495ec944b051fdf6c3b42982b1437179f0f7f1579285c2ea1bc456645c2f75de8545344b9a81bc716c5a1eda78e5d79fc56d123e774c87e5a5202fdb7d2742d717f4cac8a3a455;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcda21faaaec8e2e47f4b6d64fdf02efc23d3f0210806ff77ab253ebb3c8c77a20beb85ad92a8baf47307959c77f936002646ce6f865b78b6f8e88557c719a11c47e6989c9b19d913;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54e57f73ef526e0df9f1f66a3af27d36af5a237ec1ada8f99f46996e3c668425e928cb8e091026657a8e0607a063a94b71b7efc2d722764e17be1b771170573a16ad879207687796;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea5f0fbe4abf02a8afb260ad2fe97976f6225612ee8d032af23717dd230096683f0fb70ce928137c9e2276c5f196def7ba4f51147ff4c4e275e04d16410777cbc91e5491dd7e7956;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82d87d11b3f78857a6dbba45adb13520a365e20044de47cb6454c5a4ba0af85b6c1d24b98cc2e92bcda1291107bf039cf51f2e70ec25aa66d26de613e4481f1477bdeef94f88f2ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8815e34439d14c3ab8e3a26fcf79a14f0494c3b09bd1addc0ae6f470723fe6071781e0e2df0d1efa7eb77505c0a0d6a80aa8581146567fa38fa17a8acd4e6d615a7fa914466f109e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf612aa9db76a133636082ea48dbb9295ddacb7f97a40d1eaf7a29bbeff5937a58fe4fd458a575ca4a0dd2d5d807cada6483719b2f45dc4e84ad24f9ebccca20e822dbfa308cab6ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf34546cb1e268b2c6f062b9c477422d05f09119c902b6dc6ae89d3e2c301c5cf02e7d553b67cd15e7e57690cb10f94cc3d1fe6654558e07b6de96bca9676f34e72514d9056aef380;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73d9c65c894c2d3cfadd9d8a7303b9fc83e5c9a49c4b8532d6d7871fe78e16f8b3e4151255dbb77c69e332e91b6fd862b8b87160744299f44b3e34fe1548ef9af099487f774a4035;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ff76d03e54d3b9b1d05ae14878b64d5842326728d32e13ecc7b43a76c0643ccd3ae703e63c631f25365d63014c36cfd9b2cc88ed2cd760720cfc66c64e2628b6cb20464509dfcd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95ec32c3ab3be65bf6a65d3cbba2a91ffd0417bf0765cac62812d76eb20eb1c52f42d0998d2e9066f7f2a09956d9e6e932c85db477ca9ac8f28781aa904f3f6c34e3db57dca1e0ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0fcbe15501bd499cbcf65df0fce33e7c51dc5245511bd72cbf34d469c04d69314dbff68e298f597dd27f0f6483c766afe105e0850e6402867f052a3756349b3004f921bfb348a6d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32cfe085e9c76ad4e2bc98f1e18bc4b3cf2d83248cfce5a0d88a47b7b6e2e9bd9978ea246e6cf7868f2e0fb6c433a16ff430907c2a6119610645ea31406a5efeaa18382a5152e4e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4fed2cc3cbeafeeb44a5291199b8059ff093f0206926ad8ccb342d1a9141ea340f58f5a1c58ee242927bd39bc79f55fe5afee419cbe04d40e2c4b414590f197ce0d7b3618d1dd48;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h306c9554c1901f55f1e45a69ea0f2ced962967f45af3a8ee66729af3c81cbe5898a72cfafdba3298db81334224c503d7e81f326d24bd4d59eebd0b42505a3d8a5cf14691481588b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eeff3c291df8e25c4aefe88a46b2bd4dcc283d473b68f82106e4d29a0ec569c2ff9fc22d761896585733494c9f127b18ce442307ff2118b55b8c0426c11ecc7b8a450bde5dcb5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ce9a3a89a2d7c92373e5eed609d4692a1698b8eb14a9b256b2230fa0b634d9d40a5fe657c751afefa344ccd56124305afc0f8c5ae01f15d09f41064afb7668a6135573460388738;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22dd6036008e9df86754a96c656ae444e529fec9f9d11a9388741a68910417ee366d2b8ba88db92ae145fd763b17cdd59e183d091a18084123eff0a05e5b66fe295233447b2f720;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f720a03bf4bdeefa1061211dbfcd16888818336871f3812e02567cd34dab89c727868f2272124f3d3f011685b1162e86bd95fc24b64cc39a5fe1fab159b855bffa93aea105c36e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87f5efed7aed541c3e822613afcb3437ef779c7e22c72e204df90e1e0021d947f8823f82304ae3025e4a93567892165e05bc1078b0012b6dd58c82f6f781bba226073aca553eb350;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfadcb225bf017a48c7b9237cae8d871d20ee9d8ab19f73e1aa9e631aa96a0ca5318c04ec265b1b01a2f4b713b6b3e28d6236a0438e1fad12bf1a5e85cd35cc7b6161fca435a80a68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2f848f8ccc8280bac87565037825541af84cacd282af01fc3a41be56af7202f27b8cc24fa37b794fc6cb431ffb6f7b1b70805dc9bb76543f478af99bcb00f56a055f9f4aaf90635;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53ec2a52ba4e7e4a96ed63a40a2045a893597b55eb6fdd2d024ad4db68ab74626f87e64bdb9e23fd591dd97b1acf7e95813f440ec7ee63e35a38a0ee0246942b540e25bab1fd88ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8e200f7a8633b3ec571b11be09b103af23c2587d4e05ee2847a8f82b45a9376b85d437832368af686d2145f501b6f33ca9a78a9ffaf9b49514f097d19aa9833572560bf522edb86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1340741a06c1f329c638488b2ebe37bc17f28ecbe0e9b1ad0a5719fc0323f52fd5efee410c65dcc557fa9b0acb0e175fca3c1c0707e8d6b2336e467e8437d1413d28b7118bfe811;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e002625310ead4920025dfad3be39f6be990fb2ada3cdde3dca8207c472bee140d0a98fc9657321570ed910c08ba46e9e262307394ab73024baeb9d4d975d1425533fdc29827bc3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36b5852dfa76126578ff3a164d2ae87c5841b42ea3afec13be0e10f4fb0a7947b585fcc189b2db940a5591c3a76dd10b6ca1dd05eb4187383f9d4c53b7399d132a2e7e62905d1b8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5242de2dcff234e30fc2676a738ac1728aa77492c77f575186d22621598fdbe32c779c6260da2b845f6743e5b891dc3ad8d16e025704eb1ed8aeb7c21c2a7cd52656ebf5ee107e47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcada9e9d02336500fe18186c73128c3c1501110095d286a022a6006c7a397ccd59d23eda6826ed414366bdada31f3a0ed70f09e7c3cdfa44d51359d64f441d1173f871ef1cef1760;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f0805b1d3874dddb0fb32be6934a6d0028201b4570dfbcd6ada42adbc5aad03e36ddcb65ed53ab8616818103c5f8d396150b87c91893750b486442c2d39ae8d2be99bf3df9d3946;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4181bf130f271404aa8429590cf8cc04db78caa14c218e9f8c0cf04ce5fb6432e6d56ef4857735d5b868d1d239ec1163e76ba354181c80a02bbfbdbecefc99601ad51db402767978;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h555abad66fb05d132f8800b9613205f50e594c5618a12963240e57d3e56e89fc1baf9174621720eca45a4c1109a1fde9d38f877b182ba99a437a56c7594e87129e08059165b3b64e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d3b8286e913ce9758298a4c31ef515e5ab21601c38ce686929ca5f033c20ce6ceddb5851d396528cf4ab7a0158dd57761af9a0628274a23af41bd466fe37df4d2905b882ead7fb7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had314cec0003632498ecf0701010cc5e0a6ea02a1c2c22e08b2a99c0110a5af9215f59fdce8c66ce183a904742b2f4f682c2017683a3adc43fe66beb10b965bbe6ab8ecbe1ac619a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2759e569fae22b8d67dd55802aaeb8231ff29a09596e7e3b60c40257eb4d4fb26ea6ec89606e925dc3c6ec0d107bb7c517ecf3b06dc84e23522e7b956b0e18283a66900a05da6533;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha26ed70321bef3b8fccaddf018189f23889bacd3c6180868c1359395e90b292f81b61812925d869e2e09cf807ebacfc72e998156b6772721c193d47a4650361786a48dbd96ae7685;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25d48b878822a91a9f92cfff73f1a016b643c62abe952239506612b06e46fa5731879ff82b8a7d751ea9c7b8e9a010206eca11926a2c9a9f057b7e5d392120317bc186aa347ed0ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba224e4022927ebe067a14e0be36583b8284bf176f509d22ef56d959c19a64e43055b617bdea3dbdfe97a21cc1c2d23a3fda55e3230c864b452e1eb178c1161e54bf117d954973ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4649a087ce96c394f20d5ed564c1d523ec4e0c5f27810c1305d98f421b3ce456c0c71665ba60f7d85c081452d6bb11f52e2741397b04e6be6688cdbf1f1ddc85f7901eee7df9fd0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c98b10efcbdeea33c2950fd5844ad2d59b57ad3397f9781ff5921e22a9bbf7e070d46a229d3ebb6d6373d7415195ffa8d6c6e5aacec3cadd7d69557c1df8ee5159042809ed31739;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e5765d6b97efee07e9dcb0a4f772ea304feb184ccff86f3e9173e624dd495f2c03e5565738aae6a9d5d3c3fcbe6991c34cff98a80ed69bbf160b105582f2557fcd27d9750f7ebd7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h127be69c1b44cbe1a63472f5c631ffe730e1eff63a718ea902f643fcf1573f733f632549b6cf6a8145963845b1fe7cf44474fa1ecad08ef13048df38c8b9e2e2033a583213174b89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28cce0f50dbe871fe11d9c83d9a63f0f22fe6bbb2824f5e9445ced68923b66600cc57b3ad70e327e1bb7d67d532e93e96a5a2ae005b2a1f8323a1be650f9bbe78eaf09156759ae14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc90e726475d9943c70b92a645e34720c57a5355ce87e81bc98be4665d7ce238b01e0b43c6a87343867c8e0f5231a8ccf10ba06e5af4c22d12a910a03a4c1ec4b2c0de113db0deeec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bc927cff1b6e1695c1baaec5dc068c6d59c11188c45a5d86a39786d52dd628eb179787b300cc5c12de40e4b25d645a3ccdac232e1ecff06463aec420dc444145eb5c90675594d2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h528df9dc469940c5838d1b55cbca09fac1f31851794e2b8361bf7a8810c00e2979866b1eadbe75a638d3311b0dae5171e8cfab05aab4b08f4eace0e2f5faf8c0ae0c1d8c64114ee5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47a7e082fb85d240cfeb6329ee67b87de38e840283d9e636ba7d52c3a1584e5ee10f8898a5c6433bebe40a393c55bd33e796f0d5821c03e5186980d013190cf8d309d4dd45ab2ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habc9a22e3e5054efd5ad6e48cdd4272f6606f26e9c5b7aad97b6ab60bcf4449710a2446fe0cfa75dcfaf2f3e9c56735f283403205ac382b2fd56cc8263676578bd35e811bb24b7bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c99ea6bcc8527439353d338d5674850de3c6c0f6329501a5921eb7b468a4323c6eb177e0497acbd022647eebf26db8263bb6956728df7af1ed1f0852e754a84c068136d4fc5bc31;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ba4c81f91acc3d22994de00b5870f746f6d35a3f2a3ff777729ce8252dab7d9cb5c4fd3970309a457d73ed75e8e9cf755b078e52c6dd42803e15928fdf30a2215bba33a92e20831;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec2a81094053023ad48fd6600b965732f3a636c523f0c6e0739eadae985d54c66d3604234190231bf023f2b3527b3d5ba98fb4ba8e7789e5a89aa8d4b362c1752238e0caaac66834;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2951eb771ce7216eee3823e109323eba8a6e540622a1ab6333206aab8d1cce6e1d64c7d5f1898a7190c773b67792da3051a4ce48c26cd4dc9245053efc1c2f5832dc3ec68ba8fb3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habb12bbcf30309126c3868f56ee04abf9becd376496cc71495e351498a8065953195090f6cf10b3401af2e079d503dc44ea2604d7bd97e84afc0535394ce534779a822acce17789d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5c8950823e9e145ccba12bb97b3ca6ec5501093c7583a583912cae5e892c65de765ffad0665215a5a588e6f3854607a7b82ec4e45490fcac701037f9fc37bf167de8464bd0bd449;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67bdc6b4566394286b7f7f4fbb3ed03318d18360010f1e3385d9f2313c4eabed3aa762c8aaf18274e42a177177603b44d64e9a0f7688d1782a04ed0644eac88d7f159b1b32223e76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2064f5713adb0d1d596d7d09f78fac6b5d9991df3d4acb566e57b49074a91af5fb0c01f79e24c94586205e2c0ac46bd72262770d2f63f028b5d7e95f25b7507275a8f2c56b267b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15737a4b3f5f122cbbc95a995143ee10624f9176c17bfabd2f0bfbface460d23cdf932388c9c9906ad0f81c61ba75301402617453eda2e7c6f225056cc51932609517e0142c59730;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8046e203d2a815907cbb4a75c8553fef7a10fbbbad1aeabf525b2b6d1c2f1918f2fc7a6c241f5c8946ca71387ad888f2cfcfaa201d5327da9eae85a4d9ae53890cf3bb0824973eaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57d03f6123def4792cbf82193d1e6856f02fb823b6f0f8bbd88cb7cade59268a11069da9b058bc5cdbdc12202d5385a7ff7f007ce78834f7c6bfcd371f01302cc3112e4f0a3c7871;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89c82c6c3319b549e0f7a68eea4a6dba4427ce09ab418e85ab4be55596257c6038140a46e201067707241d361cce9e90c4304ecad7b3fef538a5559cb3f635fc8ca665433fb4ebea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc4c8583b6ac73b5f2a0bf079dabcb8aef0945eacc2b4cf55a582b33819d6cbcece3628a177dc45b9fb391992033dd4bcbeb151926a0b598b7812a794f7e2a7184bcaddc85051cd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ef129ada5de933877ad5e71c00ed963346d7f0d05d0f889f040bd2453c984ab2d21513a8d1dbcb9ec2cd8d0e40c4933b8095b997358804cb99654ddca9391705bd4f2fba3fe376;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2221772e63db177e01aad6b2e1c60ff655a53dcc4b8b9b4df7330cd32824b9b2dc574d69a27929b18d158e4e3b260b12c50e44e8c20da6761ac3ebf296a7a87c46daed411ae11154;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99dba406910c4813ba84352e624ac44cc14aef1b48313fd6b6e97910bd2a0214acba1ca0b41659c49d7bc07c680f564a3bedfcdad37b3260c84613f0425b3cc5a37b17f1b82800f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53039dcb62e607b75b8eb6c7da4b13a084b8f8b0c4ad68b1c1b685d175f991653eab895a91b46fe7332a7118c6d043c0b6025f1942017562efc64735ec92095aae3065f20b2bb9d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d90a136d8d1366372a62e0fb566506dcb6243e701d48ca8b8ca148a766cb0274abb440396ea4a14b9ba3cfc09ee5cfb6b36dd13a1dcc55664f71be9ff2959d97344ecb122f6e430;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h869f7f88ad6793e9be7b5263881ac572f601ea0bc98fb324cbb323042511d410a5b4a0cc1c9b902adeeeb9962c692fda433e524915a0f530827267364b42caf2323c5f6a5fd412d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f145032ca97e72e5b86df4123db95af8ff29fc5d8447f81ac7d927620aa2fb4ca00f6454a60bb577b2f7d6df93ffd726b847f80065d28021770272ff875f61a3e4f003bbd5f00d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba7539cdadca084dcbfb0cdb373189a7b08823ea483156f5170730b5c5d008cd7ff7548d3dd8df2b2128eb97db5178f244755ddcc891b2810cbfa67bba5038b698235a857e912331;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b9cf41ef8b19e773ab693bf01a118974eb2ba30b880643f52b4fd4dedfb4885391c4d34466c5c51969fdc51f260b599bb6caa6eb0d9b6a5da1780dbd5fecbaa78c9189376639408;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8df5efbc8773eba61011a4b4c48405acc4fa32274a14dc6bc4cb4f2bf5c7500f62a190a66030a976f6d2c241e52f4d526f6d585bfaa3288bfae2fd0522f65042b589fde2fe7c45b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829c87093394cd22526e039d256c377788a19798cfca04fb836340f9a57f7cc825a55e1f1ba71c3ad043a40abf97efefdc9d635445d33c3a1637038d6c5b19c7b081fe382582a0f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h674efc3addd74bfc9d1c6e41b2b5f57d408ab2f27b77211173812aeaf682b70a860d70de4c8612b19f5bd098d7a745e58ddd05ea54a86c00386c044e94e69207d405ad089a500b63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27cc4cb74d64edd1d3b9633e40c4a633e58d438f601cb30bdec7aa2402011f2fa9f82e8c6f7755e1d0d6b092f7603eb5da82f68bc21e58e3291a496fa954bba05d02057ffe40e7c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h846a014cc1bcc834ba3a6957d78b4a8125a89085a20214a9be944f6d51512cf760c5238152f791b2e9cf0c4b6f315c358cb6e83e8d2a8c18353554371f689585de64e238e0155edf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d926ef142c2835a428030c2fcd4fd8b52b26d35962229ce2d7866db0561151cfaafa9733e01b2d765675093329e759735545c3dedbf3e7f18d7a45ca5b196a36161ec18d319dad9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70510322ebae9443cb6d97540805afb92db640a8f26cc044400dd6fa8f94938c26c606921edcb8cfa237ce6581fdb86e9a2f478213dac6b409582746ae8da634197440da57604209;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1618864f026f81cd7dd06c65a89e52c3a24247ce913dc6f45d370214224206362e19db6e6e4b6c01e7b2f8414e6b0e14b1587dcc53715487c82bf79357f081e9da51c54308e8dd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4d155804a1b17e6156d59348322cd384ac61d32294a9a0fceb18645561cacc7f8e4fcc8ed94326620552183f505df12fe13efb6a9b0e5a6bf50e0bbdb136abc9c91e20f28064432;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0d03782c600bf4aad20c805c5a580d76812a477c78abc6fb4a21f6a0bb211dfb099f9247b96f87a2363c431901b36c7a65385f78739cbc55ac4108d0297d5e87f825f45334ab032;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0c73aeb1b2e3cc2a9e4a32e801548929e0130f129c4f7b3cd8d310cea1d905172783527b8819b95aee8059ea9e664440ffc4393d2b907998a551c1d7aff7cdc25e72b37838ed0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1d7d44a322b6c449a52c1ccb21f6e1813c6c05c70576a4ed0bf41b25f55a8fac73eef50b19e9d1a397f8ed3488c936566ea6f7901093f0ec6d4ff3332b16c5f4c91b4eec2d5aa6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6dd99b638bed46c464720f881bc48630a6880b94b3bf37df4f64e15f66cb5561019a454f3c6853ccf14ec78282da62b74f7f3c2cdfc45fdca7eb2406b9319076c5be679ad5c502a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b3feab97d83ffdef1644188a685fb8b935c2e0e91767cdf9affa9b67636d999b7ce811a277a218246829478523abe81d7ac1a94ac19e5b8fbf38b8da9c3f4a8e4471d96a9a0829b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25f0537a705b39bd5ae26e173fc1fa667e98393913616fe1dc6a505e8970e07a2a244f43fe85488c4d5058fbcd2b1ec202025e4a75e7bd2e65ffe298a8502870d1bae84f18deed5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47ac53644e82a0907bfcc310379202b3dde36184f9b7be9da65ac36d101f0af765f48e82867a31113d7ff19b4d4c984ffdfff9850e6e93a5efd612ea8c27dac7cd2aa9b2f6a4d71e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c293a05285c0b3d72027297419446821e613d3b655c8e677f656717e8ea05f283aae29eb3fd0b40f633ab3a1091a0a5aba6450316e55d4364029e8fe10d9cf3e235ebd247a2c0ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47e2b5f497b63439243996bc13b335fc32ee1ee8a3b607a76ce6fc7fdc9444c691816a762f270bbf24932c4659771e059af5313e41041707d4d514fb092406af6767f718fc891479;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70dd89b9ef4d48f170f987b495b043b068d7eb1d307ca9782bf409e84d07d82e840611b5381e5a1d8e213508f8b3e864163b054ad9c2c9864d3cc57147fb43f09a9a94ac15fd21ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80753baae76e5a5c40786d38d689b0dcce015690d48622b346f44550d721b94eeb7e1606adfec3dc33be00c683fb10d0692ce4510250fedbdab11ebd8869e9e088b29085bd2fa274;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b63cfae03560f7dec90613cafe6fb31f89bc5b139f0276b31f283574f34894976cb0aaf8651ee03c0e4c6a471e4f00876ae90263b0fbe90a28ab3e39285f5fff2eb81f8c0caf6ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h781e9ab3c7a62c5fc75c2f2e635ae16efa3f9e0d360a42840e3c0d089a1865aaca66c096db5c64d295d82478cb8db124843d2b1fdfa965ca611f8dbfa958822b379af3cee3624499;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a8fd891906f97023c9dc53dc8671bacbef4898f200142639919fb920a57bff18185c425c3686e3ef89081a7ca9e8998f9a07a483d65d13ce798b6437d665c632ecf097f4505d4f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2182c5e9f7b2cdb505715a8f9399bd9a9f3ac7969d9683891f5c4e1a7629667baead10c5a39e2aed600c71293f126dbf452bd04b22ce026c0192aa97eae679851b8b1973bd90bc9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13b81dd048f3e4661baec5379e56cf51684d2f8bb72965300ba8f05a49a35f956f18ee8557b3c28182cea98b6d32960a9be7c849f2329cd53c7a5c737414a046c2192c0f1d2e69e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha48d215fae14dc312f3bc42b1f2002a4eed819470254c16fb3edd63d6e3e5510b537bfd8ae7f9caaef2591c012dbaea131e8e931635229a1c26577e6e33747d33a43084bfec24f00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8c172dca54c3a13518100a09b6707e4f3a6819790207f56e9738f76c2e9fbf526633c7c4bbed898f39531c7886bf17e8298f459e3d68188add41e0a4cb0c229e07fc3e6d4d78ec5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79258f274b1e7e06960827a848c982b9183e90d4751e3c60c2925b0d91e5a1aa8ebdfe2a7dd37507d4017823b5570221ae156f856036f1c13fcd9ba271fb979fbb781b194a79b8b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa4b62619e56e24583096e9167fdf46476fefdbc835850371dafd007dae7179e52745a325cbc55898f0e8c82b0c45b7cadaab2b85eed29067318655933e81e1829027fde44ba5a5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66d70554e5a6480c33b81bbbb515682ceda77b420070d5c3cb7b5e31ec793dc52da2ceecbab61f283114479ca7bd37580c0784de38b897892eb0751f6d9bca0e8a79729fa7753155;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cad9b93685b6f1f10550195072687e19b3a383cac1269a1865c9c8e9978043bb8e62a1d6c8f6e03476837c58512709a5e4dc796a5c4744fce5705d4aca003e50d7fce80d96ab417;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5cde85016e55a4df3f257569f4aaee476000504ecf05345a49a81282efa194198e702156459504c3bcf7d43f6f3e1a2215a41b9018fe375c83065821ed95f82dfb860123d8f082b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36ec3a6156ca3c222cd6b5a70ff70fb60ec40e0f58f4a41f65a277a10ad628d420c0d5f039423721398573fd8fcb930a4b8e46abfb4cedb37705c8abf1fbffc5c753ff34cd792d4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bfcaf707f97bbea4adf942d5340b2bfee7824270edd7567c9291db40eb410bcec5003a8ec30907c25b7f2df5256de13865b74fda3433f814c0f01a114cab62bd175764ee5db6535;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd60e5e256e70e3a230b25b122b21c0341a9bd70b2c70cfded9cfc8b57902d63b8e4457c85772b4519b5f6ff0f9e54a09b5cdf492c48b8819c6103de43420f68a90447382186bdb4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8912647726502362608dab9861d7ef6448987e1607acb57587027c901432d6f72d6949bab5043b269a805c0b15d31888ed0c3ebb2d430540be20379ab708fbf04f29a494a4bf20e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57ce9441316db60e556b0a71eb879fbf119d78164268149a9f82d781c2736e29a1f9dfa6995960ac5ebb532056543875ea6de63df3bd539591ce0111ded0c056c4878557a0e21df1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfecd762a94ccd6c4b0eca1e992301c207642665ec4148602c1ae0e8e8ed40d91d2c9293202306b0bd86d3babafe81244ef6bb1129359976a47c9f9d8b8fa92ea10d541de1940673e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecf798c9ee388576f596a77a9f6c2c99bdff9ff8ffbe693b3281b127cf711182306034a82226c4d3011c6e0478b80279f7c4487f8365d664f7fec3e4107235ea110241a4d42143fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb4e190f7c1e396eab30b4fd3d0cc17617fb46081cf3a549bf726dc881b5d609f235a54ca3128d89cfb30376503f680f03ad294fc65ba7c6dad6ebacc4bf13d2be0ab68b7d735e74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4e36097ed173b1664742e0aeaa54c9bac1b8e9bfa8f0184ee6f2d12eb1a8d22587de34a33c16d6534ac5dbea007b5160b094513aa5734c6b22e9887a712496ef8347c29db1d38e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h915c1a34e8df042938d86dd3b5b08e1c2c81fd6f7230c846d40390d487fe1c07a20369845fcfec0837aa630caea0501091072cc7a87393073015adcbb6ea087e26b3822a829a24c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a8b2ac82beeb196f95e79b36549ae2bbf959d32b40f4aabf01798e8d806cedd260aeede87aa333ce2d7e1c0aaf0397ab9db0fcbe17cb074b9fdf0726911588f48ce18607cfe4fce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h652d55056d812c91c639aba5dd69ad269d53c235c0a4c0b10a0769a86aa4171666d09177eb2160762e9f0a01af332e6c25d4c767155d810a12a2708a01d540ec52c994eff84c7ed2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81c95eec4a7ab10256094ae6eb9b53cb391a264b30bafa486d83e44c438df9d5ae2e62798c7b99972be5569392b9d11622dd7f040088a73e27aad252dc0076c97315ef5868bd0864;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf2aa18b0934d920132727ea12c4f758682879146820a9d981ff78a1238c0830b9a4dec53c90cc5ab3931f1e82ade9fa2c0e4f92ca07b69a4edbefc824802f82eb13402459f265f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd00f42dc3180dfa15b6215c7aa4b7e15d80d07a83ccc1b65260cfc12e2942533b89a9ccefdfd0e5fee61b6c1ef0867878f919a1bbd84c046f811a6ca9d40d88dc14f1190ce221846;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30e14726d1a0473549755ce7b3ba965cb0ea7cf5696c20a8ba11a12393c48bec0428c4d12a30633ca72c40c6fe76ab9a58121eb5c4939cd956c6211fca00f8be2f31adb6f6708f09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c10dfa544d2ff6a77c7ac61657a20f7d07befd8608e4d2ea85ad7e5248d3ab488908d426816daedc0550e877260a3a3443d9f49c581a54fb12d5f1dc6b4d6e428a8de3bc08b8658;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae1cf83ebde28825478ca8849b81b8dbd50a5e9585c74720f83dfac9e0dc4a13c68d3b67b7e9084dcc03741be3543836efed584b901cf8af84679c9ac0750926217641c21b1aea12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3de8242187e87a929ee86bea6096c2d618e493547f2e7021e8880f412ad7c0e07e0b10bee8b1157d0288827be2991ca80d703529bd90ac0c557bbc465d506b490a567184e523374;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfd3055d0b13eac071aaa8314cc1b7e6d1209bf2116f16dac3a4e5279c60a7b8cd58921337dcafba3e2bd75e57fc7ef8c583f65d10a984749dfcbb7e0ba28de70074920f65a8d3d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc438e29015ce451d1d8958c3252dcc2ada63511946782af3bbc2f07f0b4b303d24d43fd325805c8586812c8fb176be6bd2dcdccf03e64db4dd38c8abbf199104f9e1c49cbf47c3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86077417d0902ddd14c7f152b4bdf97107a1ddb60b3b216b19579ba2c0769fc764328306a504b04b8439d5a57c3bc1620624475358cdd64b8507bd25f65d712032278e81b4300ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he20670f4971bcd75ed0f7bce7a7c15d31bfd8af1507331e732203adde0fb8f97d59dda8b965c668b4bad234091bef8cf4fefe5298a9a5a4f4533ece77b3706d2bf51354f2fb6d59d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dd23325a922cf1732379fd1bafe178c1f39f8e97270182abb540e7d5a3c0c0215d265aae4ecf22d5e71a0e32e955a709c244fdde1786cc126c05c433ddf161db872f2ff62bf686f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ef0baf9f2de35e282055f52f9a38437664721fedb13deeca05c18be6bb64ad3536c662284c375575b68b4ff17316f30d0183041511460b82d38f6017e091101b7f1bfd9711fd4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ac31276c9fde076164f0ce65af7ca661981e3601c40ec8b3851266fe78e6d2ef41acd104a948d08e61371335a3f1910c21147dc4c18095a27f8d92f0a72e1ba84f77fff1a17987f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d897bcae81a7651dcd5365a629f3d863d82cefcdfe6fde75524d739203c5bcdb3802b0b8bfaf530efbd2f8f9cad0d1b9e6ede4872f5901930298a1cb336d3f0a52337ed05d23f8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67449349c3e08074c0614f0618d9f1fbfe848963f655e8a219a805f790fc692c53eb337d9cd9213b70ae284f5645f862b8895542e7190a8d7f39eaa4d0ed7a935dde1e9c1711f96;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5e12423e933aa4264404c984a37510f1cb4cd6aaa537bc9a452278c2104b92c0f6d8ddfd0c95a8a0950750019afa77fb4223dfb5a4fbcb9cd2c89992ecf7879f6fbf0a6dc41ad03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81ca82c39f07b2b5c306b311eda36a06ae547bce791f12e2d8c4dc4ef45985432962dccf86ed404b2ce81ceff35306b402620c4d615a74061f897e49ad5a6f8c284b895d5a75b6ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h831a3ac47a1bc0af128f49755d3385958ad198c6b0f079718f9296aa0b5fa0d9a7a7d97395166b94a1f90ed367d1487142e19eca33513b81bbf6e8217fbcf6fa6f7c994da19fc1d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18865825c249ce80568963c3b0c4b4fcbe07c2792f65760d52f816af8a73291ce77f62f89cf34fc139e197e76ef3d0d2c957ee38831aa539cde9028c0d1ca49741f0b17e5e6501;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22ac98e8c23d6b88262d17de5cc248c49f6ec55af96c7e5bb43b79c124df2619f305feccc21c256835cce60ea0541677eac48835cb752619a82f43fede16ccb0f2ce4afc3b719e0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc02d300736200c42ccaa8b5412f84d5e16afdeffc483c0dd81f05f5e28a65dbbae3bae64754fbb0fcad6f0be757d0d5cfe9514f461faac74dbba494fef14985e5bc021075d9173a4;
        #1
        $finish();
    end
endmodule
