module testbench();
    reg [26:0] src0;
    reg [26:0] src1;
    reg [26:0] src2;
    reg [26:0] src3;
    reg [26:0] src4;
    reg [26:0] src5;
    reg [26:0] src6;
    reg [26:0] src7;
    reg [26:0] src8;
    reg [26:0] src9;
    reg [26:0] src10;
    reg [26:0] src11;
    reg [26:0] src12;
    reg [26:0] src13;
    reg [26:0] src14;
    reg [26:0] src15;
    reg [26:0] src16;
    reg [26:0] src17;
    reg [26:0] src18;
    reg [26:0] src19;
    reg [26:0] src20;
    reg [26:0] src21;
    reg [26:0] src22;
    reg [26:0] src23;
    reg [26:0] src24;
    reg [26:0] src25;
    reg [26:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cac584c5bbe1849436dfa1602c019d2167bc605f61a78c3b687a50e9c4bbbdb09906e4a2cbf9f84da914669682095f8e44c3b6c62bf7796792c7139d6276da6fe5f22146268cd6e0e739bf06532e7aebebb8ce76fc49d319f63cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29af66fcad05199d14675a9c77c0020071bf993886caeb433211a63598497fa4b57a7a505db97b1e7910a57d71f357af23b2e6fccfae91e49ee1284e1e3bf0d50b5fc03f1d681d355f2d474c28e83a92f3393401849009eceb54d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4e1a677932c2bf022212b5e27d9b9f2ac790c2fcddc9b58ffeb6a9d81631cb1c50f073ab4ee981b8362bf8e2e8c5d871a2fdfc5f92889134e302b0075ff1bb34941ba2bb37e7fb7f53045ea599c9ca6085c9abf257312c3386a3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc71ab01dc21e43c119e46364e40513eaa1a29f5f5df3d9c8afeec984b98ac878a6304aa5a7b3611e2357c8a4c49da87f3a903afe39614ed5a51f715c96aa9594251801e4ed0b1381398fff8f57fcec5354497846dbd09752e36611;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he639a1e66b5e687d90de0afad65c6cc699600fd71e1ef8a8339b687fdba13972571f1dbfeb871206d9edb963aaedad92a457eb3172f6c59dd8a64e09bf1c7042fc67b3ee1aff36ce9fc2eec2889a9e0c3a77dd7201fa547ffa2064;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fc801c357432d069115fa6f6a496fb368566cd251bb740dca4a8b239b6fef3b23b85501a5fff94ac505f3395a0519fa0fd28628f55096bcb3a6543e10ce4daf949a82a7c830090377ac22da7b6691753f8d5ed04cfffb585b288c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95c11c9b5243de01f48a0132f0f203df43a070555b1a338e219a3c24c927631c862869c77253aeac7b05680878cfd0c4965142f3bee89732f9c2e6cdbed8d323898591694923ac83edcd42584a89652805a092b549330790d0dac6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c211efca8f3ed14aa62856f2efba41ba1d80ce060ee533c051836071372686c1b9ad36d471869ecd7b646247a72223c05a9a1462c750e989bf741ce5ce9b0ee01365bb77d12554237e5341517d1f160a4ccc67bb77cc381ccb5763;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0feecede390ef2308eba6807d2dbac47a7933332356ccc549aaae97203129a3b75e7e13381aaa9f23e31de8c814c3667e707e50902af79bca5b3ad4458c37b1220472b1cc99a7d2bba9e8876661ac7ef5a27e1a5f37ed5b1335c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34a0aeb8a0233af845ec5a994bddab174529e7acb79e4f1f6e69d5b4924ee5eae733381e3ba24b2726e1cb194d6005a1bfee68c27ef42d829c9178b665ebf122927e3c226cef194e8872438122db7ee86cbf8dfb6ef440cdd4bf56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f6747c2b8f967b960a412a877f0ee3490247ba1b7b4ceab6c0a69f65e6608692e16315aaa8b9b78761d2e6cd6cee77749760a59df7c94b803e0d8e6618371894b4d712364d31e2cd77f83942c79a06a88e678ab3de1f19921ff5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d2b39fa456837ad6d582cd84be1a74b0d00f9c59b18caee866bc773c32f1f2676c4f83e919c1f3a0215103498663b2559b629fcb9f80195be1333669eca605ea1c1c2f4b67603be03fd98020b92ba57648cb3a58ea21e8c93d503;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha15e81461aa61fcb76f50f074a89539db31a0f2099c7444048489a8bbe6ab5a05a00eab603fcefff299a5134dcdbebaf43f131aff7442ab7ab597630cdae723c0f068a232f73a676004404c6890b38f34c0aee63308df2b5f5992c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89c92327284a6bcb8aa55df14ea9c3c6c163dbf4abdd69dfeba421520b77869dd0448d4187ee3b85f7af6cbeb503642470e8f388e16acf84dbe5e4471b938a70f05aede1e119c3285824a3c4b24289fe1029f9f73ea8c18e58a955;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha51196021da0dc7034c81f4fac6df3d81d7507a2b137b26967262e818db83217124c4fea89907ae3bd650f2887cdd7f57976e59ffbef1dc7da0ecfeb960b22171cfd01a9794a50563168d2e4347292971f42e85a4809428c4f75e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h651afedb82400b84705cd3657ee8ada8ceb15b52ce70a57e20eb3ae5b2634302a45b554090125f79c11b3fb250fc60bc230aef7bdc6e5d06e2e4aad3f88045da65757fa9ade5271d61ff28fa5c96ee7a331981da592101a5df8e13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1496ac4a5fd2d3420613d0baa7d61f592fc32154a95b4c137eeefd6be273c310d4db6396a240ffce7f50eeeca38c8f9b241ffbdfde9ac859c4f40d100e49dbc2680b730b7b644800b3722aa8c092a07c8a2e32f53fc58409311838e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfafdac060499342e9cb1032906465a23fea9312d45f273a9038cd8be8993c9941e8093a9da5ec8ef935101b23c3c3d317a95f85f843aff353b44a7ecdc70b91bd2629f06a5cf7beeced7084c2a0da0b52b2733025a6bf707b3516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17663621730db4ffa998b7ec8dc2f7e053701163447b29bf44955eb167b8f1d8f5470f6f3c84b39bb6a9217810160a22d02bd92292d63949e0d5f6d9f6b4385ce7ba8b0f09a8a6ed2b0c9e27b4e01fd0cccadd2762af2607e8ef0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df2f862670fd1a3a3e8147646379bd5aacaa911b1c6d1a29373b537ad947527564482c2ee93c00ab0702f409c21135fe0409b1dc2db3b2ac1ae550a09ef248d3e6a52bacf43afe77503caddee8a549dceae206b368a67209f1a655;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc1fd86d704abacf5fbd83714ce9e0155f6508ac119e6974aa5b77d85bbd6822489c404806a3b6f6e2c5a0df4498036ce41fe80dff19a052d8d16c1d230bcf9cbbb3d983defa0380ce2c57db938a22b48fa2ceb75870b472a2baaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ba65b2fab76a435100ae18b9f1d25e34a1cef5d62b743a9b0a935dd67c996c7e9a6023b358295a6d16baf0fcff70eca642c82739ef253e4a493d85e7efc56c965eee34acffa912672540e88862689630619e8d677e3347b6babd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h807d9fb60784620891ea3cae484ee66d5ccc203d0c78cbfb5162f41b393a5f458367c503428ba6eeb7b45e94d6f3b5e11be770a1318d3bc003073844bf88bc392700fc138890689fbdc8c177e9c48cfdc45b944c13d386c4537f43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb118fd84c8bb7a5fa29999e17a7729f68fd8448e72824435ab0d7bc13d3a3e50ae1258bf4f0ed828f48c6d250972d39bfb878e95157d9cc3e404317377b13e6ccae7d48c6f52b37398058f6eecaf2335942dc26ecb97186e00a3a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h778798310fbf6429b44def97671187cc3a1cbf5724e432901bf50e4da8da7e48f3478a41ec7c6daa9db8e77d448ba5b0c080e0b2058be5ac791888fc63b22dcf73776a58b85035168bf63f25ba5818c1e20e31eb51a152a4496b25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3fe598659a5af6d558cb5a37414d20217b84ae88fd80c74fc72d02e7081132e24f460036e2247f3febf0fc745fdd672aefbb9843f90fc2ceacb2f984d4994f1dc00eb309042096118913b102482eca2620f1946bda60fb326d8e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed09b8d729ffa844a9de1c802d5458341144c7a9624c218f882e5d58e192f501b330ff90d0870fc852d35d11a1a31e1ef9ca6afeb4fd36dd17332e95323d5e4b7f8ad0e931fd6c3a7882992b749b3fa97a84e097dc477339f9ee41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18403bd07890b6e26bad29a4a5bb83bd0d719cf6c95f19c6cf716f605582bcb7bd5499f74940eafebc10f2769a52ab6204eddba860defd9e54402297be8193e1c9f8660564d1fc9db3ba4342a673851eafadc2cb4538e61593d4569;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199f6ba8cff5fe5177b5d2da06c23f11dda51b27632ce9922d2ad53730edfc6a2bede6fbf6fed69024bb4506958fb626392c99c0b74a6359fe55818cb388db81c323ce07b3e39d2c49aaf69f44ca2215615bef3febcaa9be3a9f7db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e02fa14b0a59d3bd120fccc67494682159f9e39fa1ff65e4190b0e0dc476b533a28429cf2a2f112330b48b6cad2cf83a8546b68cc6a3409a808b684d4b8192d9ecefb66514cbbfa8906fbd87ae04c13f6018774f603683697f9bfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157a919be8a2ae2e13dd0670389b4dcf6d87f3bc4c6cf6d16a6384ac7dde82004defdac6030a55efc9105d87971194ea59d3c3bf14debd3a530e15b3b6027db6ba1171b244de96c98d22ff80b3e61ae81f8f40bddfb633259529a50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c3c3dc8c44522934e3f8406061c738d15fb5760370b8f34dc73b51a75766bfbd8f7c3ad411a0009f6a43ba3ca813cd6ad48d589505344da7c551934f4b51e4c08e303dab953603db4fda7c01a65d4e23e88f3de3782cd15a58059;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d421458ea35cddf2dccf279c7bccce2686c1f90d905e488a76c8355ea427e47ba0b1415e6a20d07477ee20a04b30131e5d4025582e0a1b766fef2841f28fc16e54e08fae2fa1784d4e10ec23565e92c1abf8e3354286bf9bb09973;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ffe2e01cb0eada35e4f3cbed11603fa0f67b5d18da338b6c346453c174097359b56134a8c05ae1e7e9a08d6360478720399feb85af9118762d1b6f12356320e83deaf35454db4ad1ab61696e5a138af589fafa328398768dcc087;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h954b9cc3aa5a42a288fd2f8dc429b85258bcde649335bf857f807c7122adb470f28d4dc9fc9e02918727732ea5aae8fc42d0e51fac46ccdbabaeb5c061f715efa2c4a32eb29193a192c2379926135fbf57d20d11fef2547a096e28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182476938886cc469a6417581afc54efcdc291fb23f69fbf55d94e39d1686c9be52923aca80abb40449974d23a314ea5692f071070a25256b9cc7d025a85e4460d2e018ccd1f932985d3708bab874430a614ee8eb299d138c17f0af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb26dc802003e280888f9841998b052fd738ae97f8b392e0281e508d9537584e5539508ff325dfb4d31f9c4f4088fea6ba14f24bcdecb0ea77e13fe70fd8e5dc6e0a88f50ab493b940c377ad0a0f27d7797c9ad35491015a8e5ce2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4872f37a98cbaa5f8fdc60984c03aca3cdee94b7ff5de818f9cce9ed166cd3b301aa90e1c5f3b2c0142ab34dce77477018b739dd745f6befe1eb518662b1f72da9c3d89b22013c263b6b725f5f6c1595f496836d2bc30ada874cc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85de1f95ea77ed601d0be3b20713c803c435b5504721f3d4aa4e7fe79727c0c56e2b30338ea2474cbaecff3af6b9226cfa0e03934f2d5d57edf9bf257eea1919e1499ac969dd1bfec46c36d5d1ff1fd27c023964afa2c9879588c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5a355e7141d67a4bfb2e19dc24940d32399fffe307adfd315af302a1439c824f61dcf9de754a7f5e1350181afeddecb0e5c20b84dc704562bf54ecf169db7fe53551b6fa9bcc6f1af6f1ce555fe60dfeb6516527d417142920ed9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6efb791a584a4e65ca7fa3d7740470289d9586b3998d47ccb3971659e145fdd9415a34f2b4f7b886fb66eaaaf37814dc8d0e06781ec6ac0141520ce1b53cd8752fdb5813f9573e848ddef3a8ca9fe3c87d4a8bdd7999974c86eafb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8230d4a5c7cb4bc12322bcdc4442dcd4d573daf1dc8990d359a9bee96b8661fd1b52eafc2a193bfff8438ed61d22c7fac36add6784b9ce3e268e828611eae13ad1b5ccb28afa3282139a19552b6d5ac5320ad4e9f9e3474a787ef0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2027158aa2d0acfef5f2ec057d9b786a4afef31915a195a98ca62c98098a2e19773d11adb665d35f9eb217b15d9ed1a81746927197db83116eae5f447fcf646178658e28a35a16e88a5c838030a1f8e196a9423a9742274db18a80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7015a0d6ae3180e708bd6b7692f32b3daa916837b52461723a3768ca6b3fcd6fe4421a93b65f5d73d813a81813c638e68cb54a6a4348fcd2e50407ebaf43d51db1608b51285921b0ab622853b4029ff4b5236c080f714b9577386;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fd6f5e4a5337f8772ad6f2790a4c84bafca29eaa317b9b01506eb1ad3d3d3c706d5631e47cd2878d50dbebb75ed8c9778446c4c44611260acb7657c37120a44a0e4d75fd95e1a2407f8ffb27e4b54c875ea70abea77da01283992;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a2350a343f732e40c8811130e939dd2b11e97c8dca1837fd95280634b6f4ca4edbf34e4b8a8147e3555d78ec6e5034b7121e24441b5ea6390cf37de3532f4ad76aedcfe706cd1d3253dfea8f3062ea6ed53c32db43b2f9d172213;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hedd93b48fe120a8a9408698dfb2bc9e57c2c775f3a8607bd579d704cdb3883f33f5462a2963c15c0c39139e94bec2ac6c5c6fea3268160416cbd7db53e42d397835cdada9a0b9fe0f008e63192418c3236690b051329894931e184;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf53524082b090615353965fcb408ba348c6745124f03a48126c0ca90db022d8d5793ff9b0e8d12d28473e52ca9af2b72b26cd141ec759d1f8e0c73453c61a271f62e3912fd4c836cb56c71566b05c6803f97ce177965f549576214;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc99fbee05cd046661fcd32d2d66d5f64091d65a616572fcbe35608b0755210c3d8ac913e7bbb4de034f6afbe69fb70f2ef07b0dc925c79464f5b86f672158ce5924d4a579584d05e7b5bad01dd99bad99b2b4f70088fcc47796c1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1356f2928430c605a26c450bcffac42021c199999b93d33e737aa19e1f092b2b810df4a0a9bebdf75a66471755317b37ee865e3198eddd9e8f559b7ba11511305950db951c7f0c66a6488f0ef30f801362c3baaf66158e67b81c517;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11dd9e98a82ec8abc04a15d48795b88810b66309bfc361bbc795558c33ce492153951ef4b211831d7d036aa578f2bd6c1989b347a0a1cf781435805affa9f382bcc573ca6ae8c75d0fbb129fe6271b8a32f9b02fba0359ebec0d095;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176cb3a4264034c4d5f5bc45b48466a199d55bb039cd4c9e5645b5c2e9f11829540fc7e633b4197402d616a4bc0a3102e449bc2679464d5c9ad34de9a1dd9de31822d79852badde7afb7bf9db581a28ca4741c52a63c7dd7a5f405b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2335bf5f5e3b987d33e4b383edf07a010caf49978269d87881ecf8e8af81a3ae9fd7c247f459573cdb50086bd4bd294a3bcb806f43ebd10133622b669b88e59b77014eb2e64603dabf961f615a4cae1ee9b72faff59cdb41390ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c941181e5aa5c2b6f41a097c4c2be4579e690ceb8d0c94c384cbd0a3b848573083f0a654d90d76f4b07df5a0c2d7a0cd1acc9503ca410211ac3fcb7136c9af7d1941b05d14f466ae91af53e8578e908836dfc7ed6fced872eb2432;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179a19cfaf7b17c0f913cefe18035f88f6627a11632f536bc4808f73a7e5e3c80075c0403f02fdcc13ee9a1901437274deb932ac62c69ed3f3cc6f797a760dc5f4cd8ddbc3947dc9af4302d5b8f83ee1e4021b1a04fd7809e35c642;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b396afb0dc9a689a4ac06fa8d082e04fd42bf1debc96729b74bbcceeaed6c04fb22c8f4f5357210d7ac030e3ce7b22c4f508fe000ec86f21a246448e946a084f13815082159fd1570aa6dd0b96fcd46918d29a6e92f71f863c5f69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190d18ae5d7be7d1ad4749a697c31ae382498fa6ccf372eac7732b2686f7957db46ec072b4fe733132f1412df902da71dcf40dd67649a3a6f4141fe5590fc602dbf0fd93b1cfe5d24aa704eff3a198b54478ba33de66515b8da08c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8554c2e270d49b99d8d9791c364ff2c3f2000a6824718fc76c7c138b0898f514cc993179b6f9ede83f0195e89ad48f7e339a4fdca9ff8ee68a54e39fdb553173cb232ebf2e91e866565457b60f961c45e043b085097cbdd3154d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb41336b1fa111bfbb68ef82b0151ff0b4c671cc28bba8fa25c24d5fe40ba2c8901bdfce2cc059fa8d59899725e0ed22b19fd25e5e19a390837a958f441f4d1a3dd9909acd6877a0f7ee428559d3fe3bd0585a74522aa51532181d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hafc889852468dbf46856068b3aed4dfc9ea5f7179a4482d06f0ab3fecd9c7c6517c79a963e8c005369dd4887ec7790dcc3ca0813441f4bec2d3d13ed7fdaeb4d4d82aac6be64d0979ca48d12aa984ab52539edaf56a58476b05ce7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1298aea5e42340bfab49c89150d0dc7781105ef3e3922fcc5fd9e6c5ec118515556afbc678ab3697f6c20814289f0926145886e0feec51452a86e4103969c1f809a4a49c734edc3e05bfa78cee1a3bb5444fee5690c748a6ecdbb97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2906d7ea1305d85ffef396da4b12a87e8c6d90a65ba55a2ae25428fead344739e512f67116b6807f529835138beee58dddbc93ed0575f1c3b07dae79fb8f51ccad5c1d0543851ae1e7ad52abd02a1d99841026d96d7f13b5cd4559;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164563026c2791489e2ae09bb3987b20c70f99d19b3cc18c7006f6032054be42104677740f1124b541c5a0d7bca5c080dafed192025952d72afa0df70d720b1a3234df83e00f03f7ee70cc5271da221d5f8de314d610b2faadddbd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136da34374f96c004a58a4df85bc6ab3bd86f09f3ecc227ba5e918bb1eadb9d8fa0f78a3effdd2b06fb8041e1f942a6c5dc04673c64a7401c011118a00accebfaaa28ad849cc690701ad05a3735df6fe5f3a7bab8e185c9bbf025f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b8a3f1ace8b3bd1ea1edca54f7620756c61685494b9456f73daea2b14982b321c447e3ad858c08805401b38323a2732d3de7deabe01c3563cd8050dfe1c376ea9711260f6d09ac3f878c6782d121cda5a1127d3eb1e2d1732dd7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha52e8b6a332a4e1e475e4f1108c29108673b0aa5d9f5a741492f047b0850f3c7c90234f69c2406ae8e585b3480988cad47e316f7ced55752099f82d6a2618e1503f074e60277ff9ce84d2ecfb13ac02595d47ab4dff3647cf0a8fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1266bca9ef3fb4c97b472f6b7023244bf3156729b167a6a234f5d9581868e14162729bd3d79cd714ac752cf8391866cd7169b00efb36abc7950b11187c9e4848a7283c7f9c971fab61e29f86a7d798969e2f24addfe5a6ecd49acf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h150b42440d0f92026cb232deedf222bc5d8ff8fb01494d72d8017f943aff689ce4107d0e24b5fad5b21ee63b0cc7752516051a253dfd6af7ffd1e45557a51e09f776fe4807541efd151561f896bfa3831acc84c3dc37969e6ece4e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124c781c78f1c996630a6b337a6eb0ca8aa6984d1d0344f36a3276b67b152bc73c40a8f3cc1403fb54b5d5a148508657663445c0ce0d8613da6c29d3044f0d226177d24cd23bb2b34d012bb3e6b512564be15c3d8e87d2c51ed716;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6deeda88eb5144404a62226747c2caf1d71d6fc4af54e9828239b03b09abf1d4b5ddd09239d55980cc9062f888511cc0705c6d4542a590476b168d063a05d138cb392d533c9184f173661fa4fbb3422d522c26af7dc37b55d71772;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3078b8b6606700e1fcb9b975c0ff2256011b336fb5dc95421338ae217bf3bdbf5ac87d707034cf15740f6d1e4b31393ab6c87e0544bdb57b6e97a961df257dc69a30810c4cec742d03a70e1c52e286a125310a7a771a707308761;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26ffab5062f397a7c25e6bccb1be5860b78aa90658661751b5e888fa147bd8b3d7ab33cb680957f98cafced51d05b43b5a265da15c898bd12732c72307b689f8f2e45af3910af02ab9022f41e1b130bfcb550717a9a148d2a90171;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc91d74fd66c05fb1005651f1dbcc1d4fb4ec58f8f63b7c98409d524bb58b822c6f439fcd3e17b43473484f8c89b68284efe6ee18134a0f8177de432c6ffc4f9d2a1e60cb008738dda39f25115075a1c8c1dd4eea75d38ebd57911e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90e297e13315bf3febe9d72159d30cc70a0d341f81cd9365edb88c92125101b01742d5dca199f8ca229174af4ea9b4854ebcce1a70121df11ddd05dfc65ca36788720602e1dd048d88a119832513dc6bbf86cc7ae2469fe417b948;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf5bd69d78d98ac7655afbf482a02cee494fbc18de7bbcf50d490a4dfa8e9fe364ef57a48b2dcf95b7beae1a1bbca05156f3f18883f87a158594c78fb8a8c97a23abbf20bea30b3432d87d7fbb4c4325330d74c027c5230be28763;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b7e419df9d4741b9a4ce127b38819d35c21ad0674c679ff7b3e806dd8d7fccf380e69fd3e822bbd23d8489a906fc703836515a3eda035f3fda527bf4ea4415b9dee1807673325ea2cd1080efbcf92ef9f539f5c66c005b8bb1d0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3f07dc7159895d3360a16829d38d3f4902465fc7534f2b084cd5d26429ed2e6911286f2cc485a3c74b850378a007e4cfa31ce58e24ae2fbb148104e6614fe7d83d611f9220e01650b168b3223c49586669b25735fffdb8c14b7ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h914a69d75f97459eced5f83a366d11e2b56456fd5b52f4fff3f8ac0ec6f8a828a5efd3fb77ffc35a71bd4fb7b626689b53161cca22118f289e1411b50308be47be4a3d6fff44a3ef0366c1347319a5e21c47a1eafc6280320b66db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109b3bf8c6ce402b81e9acc1f105e67aa51dd62d4f8f5a40771b246e80f2aa7e42d1c70367f13bbbcf8643114b78dac08ab056588a91b9332dd3af16edb95c1d73efd0ee1594da126ca3a95ab4f459402e7fd365c24247fd0191654;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cc0713036021834817f0875edb0b62e6ad012de6679259dce91b236051e3a8b9c9cd4bfaa601436e8945df56fbcbcf9e7883254ea863e36375869834617d8ad851f48cf122342ea3d884a283017f1f6c27e27d79c2fa3b5a7b014;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f9227fa321102a26585d43d1e5db0c57fd5e3c75a2d97506daa0cfb56d5146bd146afd3411adbbcabfd2da047c9605445a854b86aa0a45b26389c5dba71fcaf4fa7cdd56f10c3b12824028af0f21e38bab86556c3ed8a4bfaa308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd78c5482dd887f60ec16432e726001722f2e304d48c6da48b806eb2b4c73742e090b8dd2a7408bd45889a97d0f84e8c8fec60cef2661c851a3f973b71f9ca80dc3db47c7dbf510cd59f00a6cebe7245f80f5137f12b7c16ee8412;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdbc815f659a17fde37a8cb4305f195f10caa4dfe617849ab0e90a4c89ce8f155daa451d34201eac4774f0c47df0100a324c43ae25b6fbac55461b77da6a8e08a060505501adda4249e399e37b47a006c0b5de8074b0468da8fcb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9ed37c061f11ee6e68a5ac98a758b61991bbd27e33555cc571d3b56a6de5e515f45f8cd03ecd5aba87be343574ba2874219fec26d54e3b9f265826112a45b8d65a38c526b8dfca290cc78ebb73c358c3a66a578d43c1b6b419f6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ab822fd7d3d3426e34641dcc4b01c2462bb576b02dc9d6ccc75b3ee3e721894005529ece12a79a4ff1dcf0fe035c38c29fb6a48f4229c03f71fc3e93c6026f586fb7755fceb148540ddb25e65939cee55bece2a7c181e68067141;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab9e2a2d5e7217d37affb9ecee907400daac32494f95a2c07bcb1a660874af248d32ea8c8e441327e27f1480a3e84f40b9fdae27d0e49e9517e33fe63d7b7e1036a0866decbac6e9d78ca9f64b48ffececd16399500d08d6a3f24e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9c0207f7b9a71fd19cc2c320e126d05e4219b5f79abb44c1e74ef380b88e8368eab8b3d32be1affbc19ff2cceef17042b9be0905992e562f7a1a892dd653db6294c68b78c5cccdaf21ac29989c7822cd553cfd678076281d9be44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43e973d75d54aa67abb7173ff69afb5011e1da7fe126aa3e80696399ee9b6e4333d6613993fdb8bd1bc8879fcb43560b4e7fbbd07c9d1579ec0536b77a829317e4b9a6d91cabf92406e9ea95620d270aa3248a14bcc7d620f17c90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d8d65172718a4e6d59301154a4ac32d3a7c492d2f07e2de6aaabf4f9498afad3e4c85d067e69fd446d6d6002a69eb0dc0c968e534ad951bf9b7fdcb536648528aff8852326b4f2ad04a3fe9e5e624b20c347fba9a16a24bbbf26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc659ad7740bad5ecc4f70673b6bc0ed6c661d2f9c52ae5f379aa7af8e029a6184965450bd7b75791c4d02f2286047e9ed5f20c2582835e29b6c8f0e4a1229d2dec7a79b9bd94efe21ebfdad655f5a49563f7ae08ae68a0f400a6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4e3f39c8292089a6e3a696041bfbae15b999cbfe0f1eef02224ad2b0e9b2a79d522db28c18de6566293192026b67a5d0fed4195f39369ac895c2efbdc89bd696f02eb8674e7ffe1e855582f32cf16ca4708e9cc8cc2c962b95e4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102d8bdaa13bd3a564cc244d33fbffe028c1b0247281628a267d8e2250bd500c3313614919c4ea82819cf4f13da9a35a291984676095158c99aa36818d91118e3d31b5e721589aa93f7c5569a9056b9646739c80bf88dd5cd7013d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1634232d1fe10c14b6291df0948522091971c8760389f7f18d323ee0c50a5e419d92b1268506cb52918ab82f46b9ee70f8aed5e2db902ccf75c789afa65960139edc8dbaf0481feec7dc5927b7e3b06dbc4c2774bd30b24c8c1b5ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ebe2128295c2ce6dfd9e14dbf909b3221703ab1758b2eb970e8fa014a55f0d1e7bdc47fe4f80eb156b4dabe5f3dcf336f410c461b8b059e888a04f1a37d84f0102aa13d09cd76b9f541c910118c05b27279012c137724601bf828;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40d54243cee6b19cc38cc2b187560bb347b5640de9889a4f57d2c9eec85172707907288b1650a814fdbec0824b4936b282e88aeea6e0e1b1b9300dfdcef949b501c82ee4e64d1eca40674e8185e2557d49785e926c907ed8a04c8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124326bd8515ee22e5f8b6fc6555a52590d78dcecd872b828fced787929322d2fe104dd9c0e7d7dd32b8ad2f25df072b7018cfb36463596562c0747fb2d4f7e289a2496e6eba37a8472c339c11e70170afb20cbd4f7b43c27f145c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h506502e92a37cd8cd61777ce5eee7c3291b7df60a6760496891101b20a3f6891790df8707d85fddc7b4519ba3e555117b0753d768429d535629e172fd1093b5dbf383fbde3ba4bd3421564312168152feed6f04867982888272295;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9b188e8291cbd59eca9ebdcbe3d8f7b3982112c3bbeb9ff6063f3010aa65fdb98137133ca6201f6163bd58716161aa25956e60ab0a1ed55e3ee6244117f4800c006a8a5829fc51aa5e99b1dd7da41d20330a14349fb133476a0c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47e130ca98c9d00c3b0545612f022d396bcf97c97f0dda0574649a1638659b6c0c1753f219bebb9cb4c8473b88db3c6da1aba6af92c9fc40ebe708cc2e776a0a2c1faa72324a4d6023c0dcc3325d511f896c94c4c2cb0e821cb531;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf80b406ae63cf856173ab83e0e72ab4c51832c84ac83cbeb1d44b74f67958493f78e05d7822825b2890a920d3b40da92e5df5473691b0d24e520dc1f573bc7f1b698499517517d261dbd7f410fca7dea87a5343fb89bceb046979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d073f5c96b45ad148028d848ef6895115200eb5bc32df5c10a873bb2f4f9e5e223a1057fbe33f497959e7e3b4e682bd2a9f387f61b1532f7504f2e1816ef687db69064fbaeccff4984d71db800fc79ee8e374c324872e1d3b63d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144bc01b37c57c013e15366b8b0ec5fd1d7e001a558f6781fa674c364de0830ea80715833463665f27f86385a73378c8a71875f6f0118e0e686a7c1d16d5db7c230e6e50a80d39acc652380d2355a931decd281216a64e454ec43f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7ea33de0ba33b13f3eef73ac8dc6195da554a82db78cef7ae2835d86418640cff4186357a94ca58486d9fa224c2e9c41f1f3ba486774d4ca5f763bb488ffbd63c3ada481d5fb8e4308d585129c90fcf6856389081edc0c31c383a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49d73b8236ec44839e9da053babacc5011ac0ee2a6a9850f595262054d90a71ee1a507de21c5f89dcd749ba96f1d3c009102540d18c553c2f51a5a3941f43e7306b43f83b8864db38a071a2ac928543400783c3713702a73978298;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2918d711532d775f4f05a39adb0f7273a09953dde588ab988e3cd8685ca28ab45a4cc4f098267a0e4416a7fd7f31a532eba38bfc95c95fc2d57af393745ec2bc7355aa4d580d73b111ebcf4cf4f879872d802f2fa05f98d55d56f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h829bab9b12a02f9cfbcb40e18da89b2278e09da1117667b47390ec328a0e8dcaaca0b057a840f22f95acddb86c07120fa1a234d52fefa65ff021521e6d203d20c3a488b28fb94dc466cd91b51422e12835bcb2ae6f45c045dc6f3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfd20172ef17c82414ed6cee66ef8902ce06f6e34d14ede3b73891a20a0f1ae7cf008dfb3c3f6f29f6cb23f2d5a77c64052a8c12868813d52bee9ac8558c5f448a784b5238dbd14ba826b6091da1267e570caaf18c97872873923;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffc29bd68ede51ffe0a8ca76c23d42a9ab00ce41aac2556a5d7b07029e5ef4feac5a2ca87e225c0c07c8ab394740bf4b86b377d17e42b26491e5131a6c7c34623d209ce579805ccfea9257c5c6b42e888532ed4fedf428924cb6bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb226d1dac774e3f1480bd05a3e6456e80dbe8be13c7bc2fff9949d8b372f38fcbd6f49114e46913ee96481b5c357e19a189eb17f3e4d6db39f3eb68bd1ab019db7a5d2e2e33a3e8985a9bdbb0822ba9fefec023514edfe9ec48bd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb79ae7051ecae737674b0c3e43ab5caad15a332baa8bb1a5c08aa4aa99d43843c5146a21d3aae87660fb7e9170e1abaf5d6db00f708194e6331f2b583aca6bb2e1045c73dc8c0a06aebc4545739be24197417a786c196fb91da19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h392fad225d8f48e4eeee6681814665141575957ecccf4b3374fb1ba167b25fa6c22981d0071194b96337d0978b3640cbb55d40f7883751ef5faef4ce00e38635d4f5572c38b3dcbf80129c119a0249c1d1e57f956fa9095700b8ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0e6276b61e7e0ba950f54491a8ecb7fde76473e155565b721cfa999c4f1206eb133e591babc22fd8ae3c354b97084796c8d95c93d557b59d23562ce2c2af2bc7b8cf65e1644c68de97169e6f9cbb8bfe5d94169444dee8b2c2502;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19eb24bcd84b0bfffad84c90c840c4a92283e8e6c469044150dd2772f6fc9c8c1202cfdf829d63356736779728d524bca4cb40892c1c5461ddf41b64028068c55685fdced64e15a6d155df175f9ec92e372d885fa25eb20987fdf35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f456fed6f243f74f6f24ac6efca3c25bb7d3fb9efe994a08047ba89f61c8fcf5cf1c296b02eee7cc4f9c2960e5eb5db084d49703f97f3bafb1a5af3226f51a7697eb4670e474db91fb6486abec1feeb35089f1bf3a1a7e530c9f7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1578ca72e8da6526ff2fd91c99f1f38096e298f4a671a6f40a32306201b41a5491c367cf241f7307a4f0414678654790afb187ff59771fc734763cef84bc2006bb974b4892f238550920baf39602494bc7481eae92ac1fe4b7a5f79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc250409a13adad9380e54c4767370262335db46228c53419b0fdd4914b4cbd72424b25ae4bda47c467efc304e0db25250d8d108a6c1ba1215d358de5c1eacc02b92d9b764ab4c5abef38ebe73b04c152b09249f3abfbc5ab8f5bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b75770af8aa0cff883c108ae518691b56b7350c5555bbee5ed6ca606f97135c8ac263c109df3812cc4eafa6c2c06a9e5d21bfdae0bcdb175effbfa1b53d49c39fae0fc12eb536c8b9953f2d65866b68d9e2bdd456a766eaf38107c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af0ea92bcbc80cf55b3c8ae8032080058e56756424b9c298ab5a42a65ad23acd87356168da86bc0fe621e885b9caa4950e1ea10036467fc9cdc45285923bfee62a14a3c1c141de20cc729abd5517b308fc4d63a5e191280eb145f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6055dd5da02a03885dbf15d43bdd77b8f4324c0e68131720c1e53ddf644165291dd1aedd158e6a89291f719275f725e297c04440b0b11d6d71de5f62b810febbbe2e314e8b6e88e73e4e1f4b54c41463973846fb3716bf00e8f851;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed851ca902af200c27ac850f9116bb163e4d104c30ec77a6a861005ba4b397a58a244c494c752930ea6c0a05efcd040d4c607c6f94c92539ce7d048714c161e11a540fa6a8bf41f4c09bfe010e73a11e96250f786aea6472b6da3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd28be8912a0bf78b58a8e8d4e743289b7cbcce0e12f0f178be30e8e1533a9eee7af46c8045e10016ceb6de5fcf8593ff90233a0db8f62fe15f2a25a4d308a642468b5c1cb7a28caef28a7ba3ed63029605d7d6c71906917221349d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d56416093a24574a5d257bc47acda5bda9dc3a4e3484d45a3a714abc5fb68ddfbd571cbfd86b39f82073ee5e764ce8d706723a3e026b1b2fa764aa11c4fbb4c5926a6c465b9e2ec99ab8118a4055cd0bc7a7bf3d71b06a8f44cf60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bacb2197452321cfa3a1d1ae57bae9a5d6b8dbc12ed6e3041d33c926553e358701eee0cfbe9b8223a2ff668b7ab0be0c0e0232210c6c743c4261ec1c31323d55a6db8bbeb100affe1bc137a9a9b7f760e5fa3ecb9c32fa7fe07d61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h843e593973be993fcdcf14e5c7b0155dc0ba672f234435df6616c82187b92613243ebb6b020a2d1381e125efe5e7bf34fc235a33063d398eebbd96e19501ba545798f11ba9832cbf40f943652c94b98e5645776705e6040946a24d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177e176afe6e4623fe4f1d4a7b5be23917149c5b1880d709e6ec91b43a032934f27b8b8aae69d2aa5533f3b60584d0b2f61f2dcedc35a3229627c3a7c4a7713890fefae3587a91820b160578cbc5de7441e26266a85718beecff2fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1314e11d9189a3045e784a82441b070f9a8ffe5bcdc186a942d5cc23cdb4d4d681bfb6f268df69fa7c398b3e31a1c73f7b204bf5c818351ca29fe4f86bba2d590739ae599174d55233ce2a28a2c2850cd87a1c68fdc45c2d1f79223;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9acc189888f7a8df786f9e849e6b4de25aed0e9e18a1cfcdb8e0dacdfebc7cbf07ededf0b70748f43bec9fa01cd34e5f7df45bee23f74fe4a5a19e710d6c32b2455c0bc5c71aa82e217405d5ac8499d16e20a6260044b3271773b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e471dcd2af9208a3555ef027bb942b3ace5bb0ede2600f5945d7c6c402cdd986027bbd5e8b4914b47e5c69c7835dfd1c77f2219a5e3f88f6628d4fb3c22a0f240711301e26ccbefd144ede115327e948e9dec9529eaa1f863c77d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d03b36de142e36be53256e7c1752a5b4ce7eab56d2d2113796881e6e2ed860dbe6a2c29635355e545ae2e3e76b3163c9da2d680e86e69ab2b03432bc162e8a9bc56230479c0f53b7f14813a1870330e95f560958c5aa7f7e43ae18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcf5f2839534ba584f0617d7044e4f46c007ef2d960e4b28ef550c3ffa7ab52e34310bab0294a5be7a0c1d6a01ad89c0ca46b6997b3c11e8a537e5fab38841fa365466031e1f1dd7884851495d3d27b86c1fc84f3ccefb6a66543a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17842bef97f1096c41f7a3747a3c4b14abf1f04a164031a54f5bd392a5f4d82a11d8407bbf922ccaad6391598dc29fc3c2f07d6289956251981c164273de924cfd03bf924c2ba3f612aa0e38dc53e19c786722fb6f91f5e4f9d61f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f3c5e3e086ca4ec4907738fcf4aeb15d4cf60b8fdc525bd9a99379e5633732960410e3d1e222e7713d9f08562c283b014c32c4a79097f21a62181be7acb0dff8f6415a275e6b0c2f9cd02be88315d1027ab935b7e42bfc68db14d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b362e391d35222b895ff4e4b8fe6d40ac04aa19d436501da4f6ae27b36a27e926696b7d41881f74a76d90b750bf4e3101d9d4141548c9884228f2499eebcf9d4d1c37059e37161b889b648883edf49d4cd5bb36d6c171767d7b88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc46ab7747fb927e8842140fe89cc8d1e43b5a2131ff3d2a1a6691cdac91c209d1004cb07daa5f210a102d3723d1882890dae8f36b86b60d7c73b5efe035c8b37a457ce711db330a2183cf9eb5a3419bd71024426bade03504d71bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f5bfc2e2c1bf25faee60e496f258723c56fd34f76c246f047c49fcce89ee935f13d1a4879c84c838730db33fb09c140cc7d062c45015ff58ef4be594bb181922f0bd0cce34e4e93d2e0b7f9e89cb924dc55cedec13f725e6003a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df0b400a4af80e736689f91aff054a3f32615c8988ad0c7a6a0a6857f7269f3afd5d70d3153560c119d1bdc858e4250b0721fafc898085bd536c847c30ab45aacfa47614ca72f7bcdddde6c34c6d9725b887f03b779bf43f7c9d47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1249fa0e4e1377c28a5ed25ada8e9dffdacc4a14fd38867c0bb4578e3dbad9c4b613ba0c66c423df91ef1a400ff10998705eefd4e394973b2bfac180df4ba931e4610a00caf1332328fe962fcabd3a9f2fe2ad2fd673ee258cd76f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e2c5331a39b3266775d64984d203d11f542b6559bb3a06e9da63de2c84145dd5bc87dbc265ab77cbfc5755c728eac49585a2e2a3459a5d341f9bb430b321718116d99540e4126f085154a4209dbe15fc5c1c52dcb8fb431854b3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5559195c998e14552968c0f4abb3476458c9e665297e01cbca152df6639e9cfece6b045c27a9df2a3bdb2708b09016520476936b9b007b08126cb2c01fdae187dbfdf81b0732176ac872485ca236e4958c0a53bdd506a2e9c48bc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99fd9fa2e97d44158d97e85d320cfbd3b540ff9b2715006fbd56e6a68e38e15b8d0afb2a2d44451d5bd75e2d93f17190c131120c0ce9fbb1bda92e92537e6e8c269559db7a238494a75be45d8219be308d4abfa1bf18249dde10e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17672cb649f0a069ee9ff91ea97d1827e06dc1fa15ef48cacccbefcddb60e6344202a82e6a0373cb20ab1085ddaec02593017b20e5b0a9781d84fdb8dc24927ba07d6c6cc0ee5aa3cce92752ffe2fb2243aae21af8c076fce2f3401;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190c6a4faf2adffb7e0e06ea154205552be9a8feb1c0d28bdc29dde3462bb9aaa63c99b6b65538b4eafaaed103f391651465d6102eb13258cc649f7ec752262d7be88229ab283a205da72f0eae51064b8c635768eb1e2200efa5800;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b3ae6277b0413d27b973e3a473034e7dad45ad50de89a17917e1c639b445c7c7524a5547200e2551ad32ac543f4163bb01298a219c809c625b67f3192d708abd2b507f4e451ffd55d047932e779a3c062f03e939accc827b5516d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199525ab664209a24e43862619962794a952cb7006169e31e7116ba7f616afe37d4c10aa79b1bc6c29d5c9220b4da130d7452da142c8095500a4f4033173cddf34ceb84a363cc9586ac957a563fc3dc7510a2e5b491f7d6254a0c0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46cb1ba36a1a2b3f4cc803ed232a9a6b4fc3d4ce1d13d6c243d01a50c628cad1da087e37bc0fd1248671b7df23e422f07ae0bff4235b611994d189766c415d5cfa131955dd84677e6154897811026b8f1cc23e1f14982262f625c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e28b7f32406c4602122ab5fd403ad09677bbfa3c18dea937c7db8066c46e78e25e4edf16594e4817b36b6802f0cf5dfbfa2c186ce3aa0dfc97c35b1156425977155dd2b618768e9f65285573fa0c729e276ed293e7163c235510;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9a2718f1b44d507fb69612c9d8667774ef729ff43616815afbfe867bb52163263a14cc33c81fc486f183af7f4e831c8fbea7418e1bb82087f478773820b788dd99737e009b8120ac66774ffc31671cecb61109973fdcdc4263185;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18397016671f3d68ece9b804e12115f5fbdf98e2e1dc64aff1dde5ff8d821c7fcf2852101fde2c2bb92983edc165bf9ae8fedf082c34597df4bde301e465081cce451c4935b673167cec858f12a563f56c2577e902a1c02fd495ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9070375cfa4e5a1c02866e436e2d471a930808f1eaaab804dae3e43faa8256775d1b666538e9b3bb76dd0903f5c754399ee866606fd42e8f9785d1ce724c68c41eee70a71eaaf10f15ecc9b4f3a122fb25d46f97175620825cb197;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27a8f7edfa5aef08d66b31bf7f3c7d33d6b948b292fda5f72a1c9675acd3d10bb8b8cae4de273010dad8a7e635f510b4d975fcbdc37d43e14ef75ea577d65e3041801604917ee34e29014bfb1a1f5f5e10e49023e934dc596cf0b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8202f8f01e9269334b335636365a83e9be33f6147e60b0fef2889f29da0d6dad582642998f435f30c5e116c7498cb7c84f23599e044b083cba3eaef8b85e0652f35d442c6132217ca1740acd35cd8111710a913070b9bc9a47b56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8afa267f9337dc4c082920568e4813290c7d184debfba6e16de5d7a40b3ccbfe98c14464b5dd9f400bfcb19c5a7475536527a08709f47a3540b0e00936ba4eb88d6ae8fee0c4a5e9bdaade38eb5fd81f94d25e61aa699a899bec59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca0e775ecd6a74cd9b1c696299070ed172e8f9a4d0b987a05b34ecf3415b27c1966b818b336f61286175875c35a0497cea437164d63bb1c57eb54b9f589ec9c8e68aa0f1a1e4ce406e2105bfb3998bb6bde1d9edbf5fa0ac382dd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25c03a33226aea1caa800adf49e15ce30013528a05d88a594d29257053229f5fcf1dd175edb375dfadd72ca53338949a218c296a70c7cda6246542a7c884cc5e11ae349e9714ef5fb8f03a45fb0fcc63af7e7cf668e5f9c5271bf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bbae4ee0f43901a661cfa559941b8219b608e68e41e395d5b43af6896e0934dcc96fbf7c299ab09bd246e18d9de1109f693d0198df92f423e77149c0887b7adad4408c1788b1d15f35c752a252d5927c01953c003ce0b361a09b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cff4813af0fb19acef5d5ce054e0afaca2ff4183f14cac2a6b24aa83a6f9a8fb1aa8794abfebaf999984417bfa68d48c9dd9f2328f06d46fe07cd94616ed587c72b8197136ae73958587fe88fe2aa4d94f9b421f9ff41fe3e1a90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af91a4e82114162efca892371efc32524650ebf596d3baed7d5c1c412ed8705fcf5ae3736bf3f6a6b69bf2294c551821e0bc2951fdddeb2308a81310eb2ceb30a42650e913097a0244bccaf91fa0b5c57da26966b22782cf42acf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6fc69e26c8b74b31b9b900d84edc0f32b80f13cb8a2fccd0a087f54bebef557e4ff7c90945eb5db0197449fcb8d91abe30c67f28ca2c3e61a9dfba864a4f84ea635738e4e8cc343071504a347389664514df2cdda461ca6240465;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123872a4d2dfd90d58816b625408f3a1be1d679d51220d616195b27fea8eac3c05b342a2856c84b93d07e5abbca289102b2a3a429812048c8bb931caaff2d9bfb435b4f4592a1eb96a43f497649e4e91c03c73d1ac6835041fc1fae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106046a1ceb479612bc60d397448d822f6cbe5ad292ef0a384759fdcc2a4e08928c2fe841af777c28cc65c00e72582ace7cde16c84fdab4215ad8960b2ca9155c7749ca2382bffa9682f3296c4ef9711c8be83c09a3678c16f79ed4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5881cf0f1eb171dc95b4789b3b5af7820d1316fa26d5828988f10f2384ccdb15f76d6df06e55fca32d321f65cd928dbf8102032547f51b723ac80a10721781799ece96a664959eb8afb0158a23ed6ac8afdfc307e35138a929adc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5356ac20d0f933b0409a38d85cb90ff6bf334c09b4d8d78ece6890e8d605d14672f94e6153cfd6c7b90595ee222c02667a03335040bef2104035561c0214ab0e431ff1accc7b3d5f2e4145081eaba7c079ca642c45f8d76bc82f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169dcd0244974d55dbc14f8e1c6fbf632b6e723e70c77b5334cb5999c8e4f20c1dfb685e1f730205806bd25092b4ac6bff2b256d6722ed8cda2f680e128114811b0c619f6ff8f4a5a51496f6aad1b3396b7ee266450db4f26e96bd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6b90f1cb3a9bc4a52b71202ceadbfd32a77c897bac89ebec7a6c8f15bc81d66b96a5a5fdf7bc0c0224418e3c0dd12334b8bae2f33532eebf74522a5160fc473e6052bcc3b2faef1441d6230d67e9727a91319586091b7fcc1a3c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e58fa1f934f52e4d0d267cd6c5c02febf77a8111020920886ff01649b47c061a471e3ada56e6bb8365f2aa15af78554ae752c64bb6a1b9a54ae6c247375edbc7411cf9744854c6a7ed8cea537ccdddac364a1818e23daa0ff4c6cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1e4eac9dce155e8efeadf703ff0e981c83e6068b1b4611b428a72bb8aaa322dd7ad65f1ff8d2248d284b4ec8760c411d0862fce82d8c5e3b39a9563e0ae667d45494c50eb57848baa4dec4f43fcbbfffb2561f95f58232c7c8220;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a84ad232e2d44dfcb328897f6e1db204150b4484e2e03c1ed8c7822d6fe84ecd4bc9175df6f6786ad89f92bbd1020ef90acdfa3374f8cf31f51b3dbf45a84d169bab2c0bb0c801a7e115704c2bf51ef7a19f92304d82b9d51949b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c234b5c8ca6f023fbb3474aea46b2bef3c07d984c5f13510314a2a47c3bdcc6aecb1d8f2a8abb0e59086e5491ace3d7df6c852afc360e48db3877dc8e457548f8126ee4e0791975ca666cd221bdf43b75a814e72f01dbab5946ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf44f3098fe7823631f622eca6cf2a6afc0a3cadd18d5f8d203da0721121e57ea4a3c6ea051fab0ac724aae2c910ef6602b7a84323db9463fed6293e39f5c048c50885cbb3cc49541e6e97e7f1469ee46017eb8180ab06406085db1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24baf4007840215ada0a08dfd1e5b188888a9049c6a9d0f125615f409a8de379b9c370edf9edb753356eda28900dc8b2baf6127602cc9c5fc1ab455ae7913f7b827ffcbe38e519d7660a36ce071a44e95c0e7dea3a8424d03dd69c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53ec3e87758ebfbbf2941eccca880eb6108f399b4804ddc0037d479c9f68ee19b85b19efb6446b01e74bf53fcb4dbed1a6efb49cd37ea216ad105e14ecbdb8bf0fff73aabcfac422317f0458dfd0301e9c12abc35a140188058686;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf290625034dfcc6ca59b68ddd831adbebd50729b27c2004c9f39ab2bc0eb28f1a4d145d83f59f7e35a649e4c1e4c0e3769e33c46fe04727fc23b672ae55377abc5c67b8024290d2fe8c343efda7e37f568459c6b45a2d1c5df7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f15135f9f65a7d40db0c50b1ab33cf2d3c5e1e00422407a0179821202549e5a7487149616d9ce0825d9560612f1d96bbf0e6db1c9df045248de1485c118397bf1d9b243d65dbcef1b5c3e72ac3332464924a7c6323b3ed840ad8a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c6c02947893f2ce2662f845f65d9d37ab4304f138659033f949ee82698f6a81b568ccbe6eea97bc6f3d904856618013762f8e8ca209433c9536f045a78439d4272b6bdf6b2e54b49a95d184758559a87b38ecb3e4ad13ff18b23a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd71308790c6ac7301b019662070f23848a13120e5053d47a4c87eb38035535976e4ee7a9bfd38fbdfecf20161b154942428dc462d56123c131352b5139f584ddd8e8b79d4eeee0519a88532b3f06c49e8f2d1bd6f4dc9cf768c45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72fb50e111f1137e4b710db099eb0e787c92f58247f1302c70be44c84db92b3f008647dc4a4c87393e2ed892b6dfc26c7491d99cb366f19e5598ec98065b82bee4f17472a5cd39ebb23949d4b780de7362963f507642ac3a81ea48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e49506799b85be00c7b4a9e41306e42a90c4ecca92b1123f15b0213f0016982184f76b92074fdd16c4f13c0fc411242c8509929484de74f59b3eb2f813c08dfd417924968be93e0a9d289366f6b3d3b17cebc988cf120b30406a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104fcbb602047c10c24e2b817d2d94d951fedefc8f32e5f965c8aef29ac553bba15a78382b965f9621362ba83090b9791951463ec50c4331b7c04c2358ee6fe85c80216fb5afc9159038d3e1f0310190a2489d07994edbb864ec6a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba5e840114bb12ba2ad69411b24e37ce9413cb1ce9857b47e62c067845ec098aacd01402721af0ea9f239afc43cd5fb616cc1756a2f37cb4269de50a5a798b2b1008ec4d82fc41b73ca11a4aef9f7a177343682eec3748f278f8da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a589e959efaad8db47ae7782c1c5b0455c89b2bb7cbc0105bbe444836ca0cce5154aede3ce92e0d5207f3256e85650b70242859635a82d8300a32b8b602dfd2af699146adefcb8f75eafbef2d97812f9bf36daeaad2d2e19439c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d3b3dde4e87cd2a9528ec0eedad14b6a1ee6d9c8ba2a576b7b0972373ad8d0d35d9310f98f8cd8ebc5399b80d4c580ce58d2e77e65e1c6e98f584c0d409af33653949d86db4e5093a81c49b3a520d304e1950ec1f37c7b0cd41f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7150edc71b5358de4b7263f962b6462336ccdd6eb835302a1f6c39afb8657f55c34d4607efe8987878ca5e491a68b37367669b4708817993827266f339c1d49df96b4b6389daadeeae4f4a69d8f7fa82cb522c621f68947a6f9c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123009fe3c7e62282548a9e1a2a63b603a9fc25386b92befa7eea0b8f43efbe3715ddc441c85d81b3544f0ebdcdcc706a157f832cdc5285e98acde3b2b9e0ab17f991ca1bbc7e91a98c572f7dd2329e8bc4dc07e063a92d54b9ae4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f08e9d933ab2af79a72f74130e6aea0c6c3648bee97aa1c08c9f583d9d3150d172d5418f3315f55751d3cca52a98db75fde14aa7070be3b255906ce31737c8fdba76608c2efc42d11883f335e57609605b5fdcd55512d5aaa8f251;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba3e144b5e8f2fb856275e579f8384eae6e8030510a2c7bd41917114300c69b8734ad7ef3148df9724b11c67f2075ddb65e5bbbae06d8cc2c70bebb089ce382cfd92072dda51fd319c4986ce05c27575b3617564b2729870a0309c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5c802f480d1649a5828bf6baf209ca7240b53721a817e66346919412a064dd9a92e409ec8495aef4c3cfa5cb57c806493c0fdf5261239b10b1110670572562fd4b8d781ee50e61311d9b9ae79015b4458c0e71b1ab72091254729;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b77b8ddb21b2d0f7852a38a0ea1c9ada9d8a9c5dec95b44a6ad627f168fd886c8bdbe6857e301afdd1d09abdb73110f7ef07dd37998fe4d23144f308f7fdd67eb2e434ed45f5e0041cad9015460330812239da808e07fe05d8489;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e27963c21831ca15b5b11c6ec71a1fe4c3aa5d55c16c0ca7e87e9523b90cb3911876b46cec150cffd5eba16f12013c3430b962f32c35f79ac834e0cd43fb2efa42ac9b0155dbd04cb918492e942dfbb6b499917ccdcc54b2a1c84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8031257c996fc4f49be30b1e211f2afda77d772ceda8e5352c289a2d54cb55b34d146c4efbed13ddb1018e4d744993b7a2e68f8b3ed26add99af0493439ec1209602dfb0830a0a58a71011fa03a98652b6e690eafea588fe0ad599;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdbcee2fe2270f56ae2fb67edbbc660775e8b93ac098ca89461e331e960eac05059d243d9d268bf93bbb4081da7a0b8f6926af95aeb67a86b8099ba2c29888b021906c470eaf8cc5eadc45d0eed43a5c1117596042922811135bcf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f495898d0d8348b02646defa7043f093e91696c63b72f8a65dfe7a8972fa618a8a50f7f0309fa483df0e07e8ea73ad65489b634771076fcee68d313fe35d8db45f40e88ba00ad26a5a8354eab3683497eb7c21202c16a8d39532d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda79b5a98eda95110fd9012e9168bfcba564b88e934846cb9a0c0c34a28b32fa4b4f9eb02005e96f284b2fe0a98ed024007edda378946cd7d18a845f1d9cd994317b081c46b111f7e20a3cafab524ad5a4914399c90f494e8c110d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha16c101f005ed01a92851d3ee2daada8a76c6a8154298e5d39619cb227f34dcad54088c7ba495ff6180a6fb86497345e6cadec1124a4ff884f129364d087bcd399646f17a1d5d53cca68d2a1254570354f906b84390ad417b1b172;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153286b0d79ac7d6629e0d92d657c2ed383c7cc36fef3dd07f0a1554b29eff12c93256c8d3bedf9e3786747dee24188525f133a2646e7fd603de7b5079ff43c49124ec018cb1ad589aeba7dce61d6804f7f43efeb4d3714339526b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb39857eaa849f11974bdcb503f31150ce9e18d9eb27a12daee65ff27e877f47eece0dad9e020e70dd881aa6b8548133fb2e5ec6f989f1f4e1eaa70721620663c1f2068db77ec47189b5160c74ed4b4937506b2e309a34400d9784;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6f3217f58a76a21291307f692305fd8bdfc0bd062616e05992961f72e2c2c62a2ab459657774435721ef3b99f13fdd6d3920207d65379b264965ba1f64a336006d36c3417390f8bc075a089ccb54f9423cee10802081fa4ee8797;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6311b784ee8c60521142de933f6e3928c2342474e39d273bd84d966b047a1f20d21dbf33c22746fe26b6e55d7ea341dc56ca386bf5f312724373fe221fb24d7e1364cd02b152cf0593aeab49b4a2cbf02fcad23405976ad3bb8f22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a523e5edaf38b50bba3aa3108570182fd8b2d3f052fcd160c542480872d999a7f29a3ec98d914aa90186acaa2648c0eefebdf4010162bad732eb190f8a4248c5c4301c1fc0d325b7a424057bcdd8389b1c8d774ec9eb9433cebb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e20a5f2b968ea68a9945a8348fa41fe9729d2c176f2f91cca9e515c6fbe63e7c4afd181253610dc3deb279542b1e1096fb0cc32fc80589f31f29bb234cb06e18f577324f35b5e9940cc56e73ff88de6404adab96ec2f3d6e1d459;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186c652a6c757cf5a0a7f46349197d2a11a0a9a6d936e15297d3f695c82217ef6d78c2e162bf18781b9abe9bde463fd9be9c1f6ca2888f643ad823ce228512bdaec96ab11126640dad02adbcd6510b19ade506815ed425f03b90867;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd9cad676e6184b03d147a5c6203d257c20cd416480ecca4dff3252c1915aa96b7fb6e1372e84dfce9ccf469ee7cde7b845bb0b697eb9e95552d67e7afeb9806bb428c1601cfdce0ed141db25c61d6d0ef94ce8508f9fff624f51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10142b659e01f343aec02796ad4a6435cfc9109b592853f39b379a838bfbda0fa14ee8a064c96ae8e0546da0d1c20a7dfc80679d434f6a60790d5c5c5d682777044752d16445ab4494136bace1e7d8cb13abdc22e705193cc74d43f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8c2f4cb87d1142bb7a6eb2ae7be08239f68361f0217cf00a251f9e1debc0c083c45d57ab017d97e0f27a699516cd86a197124d0e1c1ee1f2bd59b8a1f039f8ed77d861115872528b82eaafaba7f90d348b4270067135ff7a388e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h298d08ec290dc22cd41bbefa1b7d4bd8a6a44a0ba9d951a4a6bab9657fec7b630eb073c21f10ca754faed30eb899b6cc9784e22498d25a3037bf3a03071c8d16ad0e412f0a270deb8f74fecfc09b32c50eeca9d051693966865a7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144f418dce9e8ff67f3e61e9a8602789fbac01de2ed9f866c0fb1a875bc9be6d90f20b27f0231d5d9de3ffbb2424b210159ff5fec376515cf58c652538bbb5dc96912c8785c9362c5973d600e731066d9f4400f79a7fccdc041feae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc53d6ca60f2a61fc1b9787cbd9bdb9ca5400b7fc75df3b42c278ee1f1f44fe4e2def168b8880a19f69a76f47df5394ccd839f9df679cdc937ae434ab29c28def3df89c022edc51ec8be634c189af15d3201cb5fe270b6be6c329d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11df35be4f463ada386d49a74f0effde22ab8a8fbe4ea748310ba10250c23ad64660b518c5b012c3a7e374b521affe224c3bd807945a0f527df8a5cd681194d6ffd68e010524d373f5bb81e13a24dc99e1568b4e0ac82a96530b3dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e37c01a7cda1bffb6ffae2984947cdf8a0537224b7f286a43c7f2a2c13dacbe07d93a2b62b7a0d168e41727bb85bf23a9ed578bc93b1f43475d472f0b4e6ab45141f0f5e5f9caebf38e8468642bdf87cba5d4526db6af5eb1920d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b90420130d6c86d5f604e80be0c5ee22cae91254a18ce639eeecf66815472781c3d006f1df658b1e43626f97cb1a32ee271225c43c1d40d6803e13df8623309ece62e4af3bd158ce75d849c21a1d56c55bb1c9635839302768534;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ce8357198c95b23db0d6a99ddfc6c2f8f8ff2271e9758c688df392729b02ef618fe5162c18d25cfae9fbbea8484989f1423a52f16c0b3ea36162f1846a0292c93544df1038ba45d62d50beb8984fd8dd0ddb89129f68f286005c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d0a4408224c3f48d4dcf94bbeab02dd783a78ce8d6f1c8f48505194c22915715def0eadb52debf093010f81a45f1dcf0241f3e2611593036957e4b3ef7484f59594405f66a723fd5db6dc94448ab7025201f711f98b41bfeb04dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf624b9a969f8032474739ae66b54c6703d839fd26485a7f75c79f86f925cefd667622d441b2fe0314e2a637786081c5052b82b0105061ab3ba520ca59d2fb4762540f4de474c4479490d8e708c9ea2cd7064f1ecf633e781d16537;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf55d0df42937c0251070e130468366affc90573e177b42a8ad4eb3d43bdf09b857c9c531a205edd4e11614f55370af853149544f34191ca4d4e49000f5d075fc9ef5006fb02866fc66af98945fdd1577a52933f0fa396233621aa7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2dcfc496690a963fc4869b816f063b97907f65738565ce68e757a0af19b0260d05ab446f45b4ec3c868727c836083b59c53d830bd0bbe514f8359977b5a9df8bd8a000553ac962e9abb84a2a72fee10d8350e6fcbafa063073f8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ddaab1436273397c7db08e0363cb0d654e14382d355026d8e7e560e079b9468425ac6d3d810d53edb25aba3b89e9e51862555935d9751b7b923533ef2452413ef30814de2fa37dcfda194989cfda9679ae7024cfc506d86b0dd44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7854d08787f2c7d45486a92c418cf2411e307ec11e0adcd1f3322103973e94bcb6dcb694fdfef244accc1144349c31498609a4fe1f6765a9fdf21ebfcd023c2802f98993e9f8398d4892ad3a7423b9bc8cbb12240cc3067f3622e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h485ddae740494f3bd58a1cef9954d7bcae5866910986394b9d831f60d860f24b1868318f11116305b42790bbbb436e66a4e9d8fe6b2600795baffc8ea60e357a861ad6b01dad59340c1dbbe5b7f86cb3d6b8841e7c706e82a94c85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbad43bb6d0cf8cc0adb6f73f75384fe47f71b40cdb5c73b6366b2dbbeb75a7bb166fe96b1a4bf9ca43f12ec6606f80a8a40fc27be83c7eb5ef0ee56a49f97fc3fdb2005590ed5570906378608b467e330a1fec5cedd99458c26104;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183c37a427f298d318d9e94b628f20f026e654db82d99fe0e8b751b4bfda7a82177ba39fab18bc8baadd9f01b45510559d6955a0317bdbc79593e545fb525a6cb7f49a968731a6ac8589ae54d2b28a49d707bca9049def1ff50eedf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1f76e9f3b861c13a0638a182ab3c80386fb8e7fec5963a2e8d6f21615e066533a56110f342bc988ac99923300a5f6f3799b843773af8d1a4f99d3ac95f109e4b518df3c3f79b9d0b1eb303d42e6489f23bf76853ff70e157f4b9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef4f7ef6ea3919fae1e3f8f63e25b2314862cc80fcc00c5e7e00678d9619a22f1270b68075567301730c2a891cac4c80f4c8e7d0049ac099fd44282a6c3c323d6f392f8b983bc790f5e18e19720e695ba2efa0e06cbefc69301caa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54c595c3e329b5355877958375e5e8493ffba0f8332edc67ebe8b25581fb38b567b84db7583cc8b5a2d8a38b5f015ff52d6b8501e9546d467d9c797330d18de871e4769aa14436875775e7c4ef5660fd38151e10a4449bf55569d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b680ea4ac280d06a7186ddae9c93a9d197f42789a627b387d0b7fd33f4dc56b821f92cc10e3eb8596e104350649dac0d9aa606e528bff6f94a7899d30eed09f2354d84d06540f1c05e8621ae91f8ba3263b95399d771212bbe22c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb82effc843be28729ca0494931bedc13ff0bb0b54a11c0bc955293f8a72eb89aed6be1a882202442d4e3ee54357a4dc031115413f65b5cfc3b6699c5aab57474203ab64d34e5b23c243fd4c96c1c51d424f02c113ab74c3b2da2ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119588bdf28ae7138401b5884b4a07b23633fe6a414eaefa875617dd44788e336d160969b7fd5a7e6a69c5c98d4913784a161ac8f4300a0ba8807bce51a404cc87154a523d7f18fb8cdb9fd09cbe4e7c7a1cafcfcd9c37c4d7e5cda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7749d2238c7ed34e7fb72d0cac7e7cf873291476607626cc450b7683a823093ce8132bbea779b39c154acd73def764dc554e08cf080cdef9a2ed93096ced2056ce09064dd5479e2e12a757b392e570564cadc657dc3c6dc7cb0d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4e7abda0b139fe32917b1cb52145c6abd380fe8a5fc34a886753ce7984a18899495d713f028e7736322988d64d8ea56e3c43759584f1eb5f8c5db0019362f171261f62e63bf6cd46ab60800602d6f11d88d1682bef47ce6b8bd93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122f2717034a01b5d1bc40f005f061bc137be7d395d3a5dd8fa3be804fc5570fd91ba500b8e5223cad85deb0fe5c0c8b71104fdb633f5ffeab0e753387936ea86ad99b630f8622e5a2266538cd2b520ccca6c6706661d3fb45d585a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119785a20931423b173ae7b63be717d0f43e5f366224f9d16a76c673985a35267b13e8dc77b6f30ea90d95d88d6312385386c8446b8682b9b7044b5a44b4d3ac9c112f0f831e7cc05b4f1fcc500e4d7d0715ce6a0a35c936abf5e36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee1e581ad3aebe43c0e7e3fb2b96aa23b44297315a81ebebe972320a3841c00ead637a848c73a68f573588391e39217b87313c7a17e1b1e86de85f3d3e7f123e528a032a0b5b4ce4823fb252d6402fb1c591f657c8de6d453fb4a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33a009bd3440e19ec1c37ca574869712571546ccae0c5ed15c2501b33d116a8f4b5002da2bca148c9e1aff53bab7b079454495ff042baccd7e17bb9d599c5e7d04e997d34f9814d2909fe98031f40f186670f65615bd20ea23b8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5675059f87ea46b6429135d0c8582ae12f6448b3cdd52b5c7bf18b6bb72fac2b804ff98ee4111d846fede47fc2bd858231ab76ae4cf145bc8010e4cb03580f74c928d4b2174aa8026aab2cd50cd2730e80ecb5a2aebc1bf5cc7c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115849b1e5465059a2bfa6ccccab4e430b11d59eb9ee1ffef179d7b37fc2e6786dda469468c4edeb373ee14f6ca44c675e6ce804a3b6af1394703a9847709f685669ce917294a2e12e482b13a3d040b5df7a339bac5b2c69f9320c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he41df5b169f332e34bce1f4441f62deb49a00dc07f556f454a5cffef6b7efa1ea9873de24a507fbdd8884f484319631c407d0307cf336782f1765ee6685672e1a49c3b7f149e273e7d8248930093ef7f998a8e048a75d6e5d4e7a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a583f28c2c50d0ebd4887928faa9c46a48a154a6e01494197a8c4f50f6488eb13476e4daef2436bd17ce3cc1643b1fd76eb1ff80ec74d7187739f6d38c7c2edd100ed80b0302270dab575e7676cbd16ee55361e4749cb9968b25d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ab53d9665ae6b897aca521dcd82a21610678b54fecbd1ef4d5449ffe821dcedb18339bfd4092fe6c627cbce5486e33d8cabec34721fbedec9fd7586ff58de40f377a8fef58d25c235486ebd8879e80c93cee7ddd8657333434f4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc139941750358075e5fff56b4d9b78aa6a818127f024b0983b5ae79632401df38730d0e2208fac67979c81858ca4fe1b001de6fd8da0360dbef042535311ec25da384a8b1ea4d90503bbea92b7e19c20f1d9b98721fe61adc356b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188fe0778b675b93c6e8c6714559a8e4f95d4cb2b9a57c45b438a1fd2b2be9df69574cd21918cfebc7f3e3503a085517501d065b2b90bac80af2e7d56e279f7dcefb7c8187ae4d6a478b89c9ff2ac427a46f8fe3c7cb6d609278eda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a32af35d78b53df45adeb1e30cceb5813bb7d34157861911e653edca86a923d81279127c869a68c5b9d259c9909bbdd9c539affc0c92d727a60ef6f108e702fdef343642543054000c67a3a873341c1b8ba99c7d7ef7024d909251;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187d13afd7eb42ccc6a6cec55b95bf0e50bd5360ca66b6f0eb1aa01e082f121c2312d5fbaffe9202d022ae02665f640feaf51a6d933673eeda990bbd14acf99c684862edf62717f45f085d648c6560ec6ff18487c764673a41c1d92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76c9f2cadb8056ddf40becb8a53527a3123d412671c6910c69f10ed1426a2f58fbd0aa496c1b7fcb56c54c59af4911aabf8f6f7f88e130fe7598c1b5de8169ceda8bb3cd5011ad9996c3980c43ed58496750c7ec810300707a089d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b74cc2fa026b2a5b880fb80f4c4c6b7666004cf3154ce11604298cf9ff489607cf53f9390d2fed5ad46d287afa488a19db636a4ebed1de7ec9fb56c580208f4312dc13f025b4c53db3a00febb6c6cc050c5e0718bf5842c0c88271;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10437753d41e768a32432958ad4d0e5904642178ab79b3122961170e38c4e670bbb20f499c97f9edf51bd8c5d5171856128c536b98d4140a343aaecfe775f12e3139306119eff06ed53b39f6645a447b06b1660cb712260d2025c77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d79a74b0bb9bb9edd7787ee89687371bc3f3fda34cdcc3946e1f1647dee7290404f231432264b48d8a9f442888c2d9d370770fb013749d05be0e6337111ca130a6fb34daa479bd51eae01b30834ade50d68244f742793bf2ae4ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac9fdb63be489c5618103a489730d97abfe8b0cf13edad484ccd01806eda522df7ffb6c05aae4833885d6aab081d5cca267e69a67c210532164e468526c4400e9a62d4d87a3bb443f2bdfcb35292d02db1c73ecd7323ff3586958a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea237ec75b2e86a0ee9f2da150c0a8423d0e27f0da6e3518ce27b0517360cefe7ddc0511d8379e9e8ce1da47bc122b66048967ca11cd0f4dbfc55e93116ef2c221c36faa4649027929f021bd99ee77c835230a5c107e9f6cedd996;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57d23008eec3f87e35d7b63e3c8bac85e83b03460fdaa3414189272de366b536f628dc5aa68b51cfcbc8321ed2c29612787117789c433cec1431b0a792b0ce5df50b604f11241923ebd7b3e72c67489b0d52032c8906ee2d839a0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b1a82b4ae4002d639ebd48552499b6f1fe3e971cab1d5bda4d6774a2be08b8842623d7485de2cb7750fec1c45bd21ca834696fad5af318af2435fbb136c7e5bce3861758d040d841891a84451d7b887aeb905e5fcb599603de936;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90f7684bdb1b2c039574fab9745dd35e42fdc4e498193168e3edc1f6c336e2850a646dc6089c11d08ed4a92d6307b853aa1ac6be554c70c5fb7fb3df441bc26523e2416ddcc14a05d083610cb148529afcf97d03adfc65649aae8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170a869588e9eb552f3e5c3de873fed3a9ffb6673333ea1e9bfb86e796dd5aa4b8a02b31c9b9846c9a7d0cde3c50bf40a49d1705747072ef61ef36cbff53ac2f44105cc199019eda282dd19d3f532d1e8a114c77861bffae6d15335;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h770029100338ac6f700abfc4140ab35c387d8476eda347475e841269a82e63fed19db3f2f7d03c1c474b227f3211d316497218dac73c530fbf3ddd2e52b9e03ca32bd8a79548193ed5c7ca2635986cc181c38ea7964b255641c476;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130ced7ea9339175a7b204d2e9635474108fe667eb387593c871cfcdc0587f5852a06ee9bfce6e617122f80c189252795016056597a3f38897d23b455cc2e24e1535b0b52ee543a3bd68cb25bd6eb773d961c7fd0304eada59c658b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17436c3eaf128845fde3e61ecc089ba9af088e95387e303252548e160762f52a7dfdd0b2621bccf941a844bbeacb68003b60ee436426cede964b9d2683d82be8fe5edc9b67ac035f77e3641258ac74c9a6b9e609c5089ad0a4b140c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e01c4668d4bbe7b3ce7f5b4cbeed3de67d2ee593ce42da6553a53b4ac02d7d0ff2384b5748deb585db95944a1a3c4c6b465fd96dc020442ebc01a9521b0291a42839da33e181f86ec426e66b5e7b217a0aa89de648214ea54d583c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcab3ae930d0e2c376acd4c78b57e6e68b1cc512b72179b83bb7a9d2741d000b2f019f71c37fe68fb60ba58b61ebba9f407d77041ab224e364f088388176d4dcc3978aad04287cbe0865ec51e1ff02ac116fdb83268f711e983a97d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he78843036d04a0e151673c5cbf1505a5d0ef28416acc64fbc681ff92fb36d2551d7e3845e6469dc467ddce459322df970209a6328e06ee583604a710d402be00f69c5bf5ad7c806a4850db31cea08865fafe6441e0aca9850177a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154bc8b9a3955a3a3422e6fb142713960ef58babe52095c21521e40f9fa1276d487678b9505051f06d1f0a83bda876f0b66e05ccce5eeae9955e381f205e621ae74ababdd3d43e63fce33b0ee87d524cb006ca077a24ee01cf1ff2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1656360fc0e7f5c7fdb2159d13b6f0a8c1b80e440c1db74f39212ffef56f0e6f175cab9aadbaec31b64855fb5388270f622acb2a7fae8d0bfef70a968aa256863b53c98c423d3ba0de5a723e625d3c829a9cf5116251f761b4b9433;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72b02e68297be1786064f11550fa4b27d967213b7b6069684ed096eddd202fa66cc423f02b1a627330d6d995c5c1f56f82381140bd54d963b1b28772b5f2c70d588a5adfee3dc09cc23a447a7935106e3eeb8570841155cf857c83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a46b32c87eec3dc3d0757f39169421d82949d897d0b20a571653e46c40385897af049627c46fb5cf336a6ca5b9ad4577034fed906f1170037a7a4f59669d0fb6120ab292673235c2df9622a72d1946ec1c7001d97b2952fdda9f30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3fcc53fd82f10b725dc7bca01dc598a158d22073f5f90bbcfdbfd4765a650808fb75125c3f6a8b785508b073d5ec8d5d3de005d20ee1ab75f1bca644f5322e955c784e6306d1db5c35e3272d0f2548cb2ada8cc61cc33e2616695;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2f72b8cf62b0c716409e69f049e416aefc2068b82efe3c12bb6b72d2545178800ca0789edd8c5c5c88879ca6cc8dda204d5be567dc0ed6529b9660648c7f1bd68c047f13d9cab226147c4f3f2dbe7b25986d7b7f71e7628d2a2d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57c7ef63212b7ca8957920762406487a0bcda6c05e8d50c28739b7dc906c74a02c13eff2faca91283028aad79580e9fdf2e3bdf46d7c2409a6c891e48aae69b8c699ef4b7355f97871175aa202b387f9541f7646c4735f7e2bde94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1349aa7925f71a46713368cccfd1985ab312de3ed614e03103aec07ffa48d0d0df3fa7e24602761f5e63f7cd6fe075aabefb889c28a7f8f3561ba3d13627ebab9d5dcdd01badca34c6be678b58c56b92617b851bbe833e266da3437;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a031fc12c6f2845051ba75c3b66b921d15d963ec8cce3809e3619bca90304eabe590326bd3be852b19e85fdbd9321bc69a38ede971aef9545bdf22fffb2c3ba685cf066d5ec81aa119f10173024b131b4b356462754f989f52cd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d6bbc10148b7586176a4d29e4eb967cc70ff884838ba61a0f6c243dc086a223a2c0866a587e781e0cff8e0aa94b6f564a3506b428e5d911c3fb6afe73750678fd27e2ad60c1796670c7f45ae6e5a6c506b69e4759c0a1dfb566ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haed8ed24adc04572324f014be6d80b9434debbdbb469b664d04b759f7cb42ee7e9e420a0d28022404752a142f4aaf813bd69699813c86e6a0c4b6594be269c75dd2096bba25a8616a856d253722f0766ae5d9a402d8e3bd13019f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c2457fdce0fd883cd98f9f541668e78f9a6c479dc02c46fd6b4d5223364acf153d6c6b0eb34a33bd35020c9c41535351417d382290774a0d9bc0fe5f6624a55ba5786eebc2deb47607e3a0a8b147297297e8f0291045205c43519;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14647747d50493e30fc8ee73d91455ec8535675f38f7ca158c603fc9b657706e1b8fc7c0a7dbc6c3deef466dfcadfdc91e5d2ed0722dab196cde3c32ee90072b13cb567a5dcc396a83a5e1563a9514601aebcaa2528d07fbf64f143;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8883d9c815521f98511a31a7a4bf39a3b7bfeb9f963461430de1c311c494ad7a69bbadb24bddc6b899420a52125245231bf424e71dedcf577f907b372260c518a214e4512437e3b9b1cdfb6d8cf98e33e47d397472b27b713d9cc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2543c93dd6bcadd33f1b3a909ec1c37be41ff32fde16549a3a6d5486533b8a846b7eac757033aff33cd0522dcb600c197021b9f9776779252a5567d1286e0bcdc7cc6ccbe4b57a28ed36f67f424429fb94b8b7c10940b80534986c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176d19ca9ce72917cf7ed1cc2c29d56872460ad696655c081fa99b6be8328b0ce2413735dbbd44d0a7cf44b7c6248d224c9cfe9202454ec252df2b6aacf5e129b2ecbacce64e1878a6979e25b962ea796a39726cb7bb0c6f54a45d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c3a537c1a5460bf320333ddc3eae12aa75e9aa46874d639d0bb07b408b8641041c651276463f21b752a44718f7f0659ffe57be704049cb269fd8db2e4be39818a1319d08ce8727876b6fe30bc5c76ee2e29a203a1299305044ca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15bdaf3062eb9a5c808e30be955244ef1c87d10d52eaa3b1cb9ecb313d118c462b966f6eb030245b31ce41929087e8692917d694fdffa5a9362978070e06486a12b5d7da28420fd291bfb7eb1605c3cf77e9ffdf5fd11c0be62378f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b3fe6eb0fe3c61fd01fa1e6edbc9597badf4ddbe0b965225d00179be42235f35f43cfaeb4b6ba8389b70eeb7a1b5a51fb4741ef47e3094cacd35d03f765ebf612c00a8d3cb7c9cd916bc3db374eda061071932586539aa928a68d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he566fa5e466e7d57e8638c211c653100f47ff39af06170d7173ca8f9d4da455d49ade21d3f0b956c4b83c26e69625ec9f66ab93795b0176ae8aae4a7cfbd55fcc3de65d6ba0d0651b7b83bf7052b64ce6c0c9e34380dea6892b858;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111580c2a6c984069c88ea8e9e5fc063f4a62136a80a1b8c343ed831380f28129edd308f3014886d6c47ab0ba8493626b7b0d25e568c5ec5e0722e414f2808f6b0a40a52a9dcf8cafeac0f111f935e519771534f18126e96e2ea847;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h317cb276b756a3bb49451f55125467bda942116920d17132ad4efd5aa6d90f7745b7f8335458e1ddbbf9fba0e77110cc978188786cb513883396bf33583b021352bf313ab1f9cb1f3f19933f2599471bde1b80e198e132040b10b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadaf09ce733a0d136e47db4ce7de5f49e49ab850afb6157dcfb9e3e9fea4555b459edbd9a94bc0b822ea3c5f9b2265c08c34a47349f83f9d99463bda2a29c0d3426c69c37e49509da8a7addb6b7d4d9a44d3bfc9b4dbb332c5faf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfca5bf943dc9e742af85b1bc4e034510fef42e2e94940d8505895df0f51f578a5f87753b3e954f410fe2fc0304c9f931eeb8c458c0ae621dd7c1acc76acff9a62ad1a9b990fccccb4a0b120cbc72e3a1e328fe08c88548b254423;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbe3be2df15d244e7bd933387ac72f56973de00c2a9ae460279bf5204610e55a819b4de6f3994785f6f08af504cb5a26502026850859c18103c33a552264eda7d89a33842ca6887a7edc678985c9f73f979ce4279655037e581259b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104a2de80cb5f89f5995bb65e3dbe22915995db4109ab1014b65fcfc7b67be044b6d7cf3d684a3e905c4b1acb6686089665ff88c22643ba17ac35f9470881280193bf60671bd0c511b61b077708e02612728bd3bcda7ef217aa08a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cdd88fc5a7127b49f956dde9bd63ef310098ad25a9c7954a3b1b4be051e7255e726c531dce0ce6b59591cc5d475395fc74f10170abbc8348eb26d50ef77a6dd182434a54bac35b74343112fbef8a9de8eda92703a93d9b3a20056d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3260b72612ed62d981790be77a386957dfd140404fe6715bc4215433603f45e075dbeb2b8979d824de02caaa38a73e2cea7bc96e72b1f7dfb6fb4a617e8d7cfb7569e999189b0e076e6a243be46d0677796a8548b1540c14590bb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdaaeddf3efdd360f5979a9320114ac3c9b0b4b95306905e713ae739ce8264d668fa99ac4b4af59d8500c3726d3fd5edbb6c3d47e7ca1b468bb201c5d8ee39f9b402c8760ade538ae6f4324c1034c136b3891b11415ac2611d0859;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d11b5649cf6919e24b1ef670aa1dd3ca9157503b9963979a2585d87a4f3756a159048ef78bf0e4b8f952039e1eff17ffe6a67025aec8f59c16c3daf193d5cde08a1109514d9cd1af2f9dd42bf305c40bbfe588d861d4c80891c02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed9accfcb358ee45518d45ca01f621e9091a8847148f73bd41e643df5ed2017091ffcfa437c98272abc5f08d5efe0156ffe6eb4c0aa5231c981acbdb14441abc3a41f4a058cd9c091649881b25b8db213de9cb34c80abe571f789c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30b2a8884bfa85dcc4673f96bea83186a5df5979b18d1fe0d36c9a76285d8f6955b651a3ce97b405835841bf569e3bab56246a2c0a2a10f0eed7a6816cc1dbbaf164d15d3f95360e108a3d5168b3bc4dbba612993873496c355ebd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73ba536e67c0a1f8cbfaebcd73d7d858a2e8cebc363e06f88cda288db9c7022ab69bdb22415637c7bb0483fa00143a1c0f43158c0716bd704ff207ac994240f5513f5bcb1f42980879fb3960bf498aa8092c0b5c8e5890cbea7992;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc585a10ed2bbef858eb6ea5f2b750f9c67b57ae53a4f6df19e781594fa658bc617109f197b6b31869b93fe97b018c332d3f055cbd128dae5e9f3646bcd7a46d021ed3a53d6fe559664740a7d6c2429dc3296956ea3a7524bf3404d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a0487bda4562a64685328393acb7250046aad8b5b9d9c81f7aa4b326155a0019fc18e05625b8d47fb0dcd94a9f37e10a7ba51a89a57131fb441839ef0e56d9bab4c3d155b389e2de1cc2343b4546a20754525c073b1b8b2ff5709;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14fb55b395477e624380c7eae2e6f16a50c6da152b294fb217414edc754f7794cecb910f93f3779faf7191175dcfec7edcbf5c9fdde10a6e0daa331d097bb6270cd193df982a9f8ad5c7d05a1e7723a7336ff4ee41850e0f0e6d859;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8396951305b921af81bcec87f298685cb3e9d44930c106c39a4334ba0abb41fe5d3f663d43fdd5f74778f89eadf588946d4f3c45f91bae7b8d2a5424bf81e0f81c2f04ef4ac9b54f372594fc76e1d192b361b03498032693a2722;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a99df596b80f14587e4a6fbd984de0816bc197e686435b7a240ac0bd878e19a023067b59f9cf6c789c72b8315f0bc80a996207628671e6e4b8dcef2a7c6f8244ccacfb382ed7763d59445dfe00cb38e1e7458bd02a2a5509a40f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c75693562fc0c48be24d0748da9c02db42b51d73382185ba92e411c1e41177da9591546b59afb9056fda7d22aa420d1217b698fdc6d17fcd777e757a1576afa079a6451cba4fb6bfb271da370eff9e0ab23d1454002f91fd84ef2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85f3a876a3d9a70b9b9651a197b21807f39531a3b0ac9b5ee90d4cba63471f9a94a8b0f746e7218afbc52e6cf9483473a862ede51b23904a2d552908c6aad7921b5692910b43b00f76d4a380d1d7723b25f2b64c00f82d6a252c5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cf76b5f6b4615d17a8377b55d696f1587fac2d87c72d8a523756f780115d71e428fe07974269676fb22cc46285b90fdff03ae0efbd1f60ea0d98f16313b8724a5b0fd393437cbadbf4995a401eca70a918fce3161312f9b8e5b65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f730c7de9511d81075d597dd3a027b0d336425faa04520f16887610143a9464d31647d4665ebb48cc1b81bd700beff991c03b89b13d8949b8ef63d5c106c7b27f123a238441edce4d7cfa5febf3173e894b8699be2ef839cdd187;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67122edca19ddb4b528fe066e3445235957e15ca2e66754dfcb4939599a6a8a3138cee9735175ae0186fbfe16299498a8f4a1ed4162c5682bbc055949b0ce00094377a73ada7c5708a63e7c95fa60776c172d7c6158d9e80c42c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hacf290b583e39c6dff574b2a06b871d01ec64efa3b73ada6a965fe3763cffd4aa8cbf61f3846e2a3078b570c1e9b12fa9e99aa45512bae033067aac572463aad69495dcfdb8f29875559d2f37a1f8319e51dc8760b739c9f7d64fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e50d6d49a966b8f7345c8ef1040d5033f8a13b1bb568e15edf2ed3fcdef789c1f0175be30cd00654f49f5a6265e87e457fd33acef5a537ad9d551a9b0f6656c20b9872a82a93cf7a89d3961787e31d69a183912ad629e8106ef09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d10648cc8197834de40392edf1e4d113185c8e71f58da09c7a2d00d69a4e033587ca9b40f597580b22ae442a0466ca99a4500fad7d94f0315595dccc5b15b553909eee5aaa795a96fa9b1a3c66d32e2f94cb7fce09a4cf8d751afc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6da3b6bd59c12e50685bf3d07ebdf656d2e9a172b904e693b813f5802fefd975a8fc2a6c7e8d65d1f1e704dfdd48f7db9e472a35d2cf32d6ee553d924e47567b07ceba530d1098b10973331c108f101563929b846fd1e631393464;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1500704eeaa50a84dd3e28b7cf14d3fe1213ccd3ff72d9d9aa9ede5b893c871c280682f53f2a110e07f285f2c8d4135c2a5a98e6bbc5a0d49594e4993c8e2b5ad209e629668676abc4b5a52e4f18c03a801bfd01af7d45826560a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h766b8e2c948c2b7c29142a20eb5fc87288248b78ea8cb9434e065541c6c54fcf4017e035427e277a00c9fb86bbe34934f31e494da8d7b4fac0adcb9ee59ffd28e2908b8d183d30ba279dfa6fb42a6d07a59734df9944e9000ee574;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha77bf33599512a1b0032765c51dfc2ef7135d2fea32db7e75512f423838c4fc0ee55fa2ab92b33f6bfd0b60b0aeb015ffbe3e9dc3b4ab0551e885aea9b3cf62fb1fc3a0684468582de67182e920da5b8a5dc94407f7adaed671019;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff977bbf1d876893cb1de58acebf2c04b8fb62b7fda6c051b72079bb830af0de676471700cbb6ba07e3a9d7351858cd269ca7ac62514c672ab49c286207a05cfcda1fff731a5f0518b173e9a70b2db85d55a746c9b7d38406c9b1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17359d638159627f2a6fe05f87830e70e5f2a02ba323db59336a8b5e449eea3722c73fb15166d619c7b7075c8908fbd84f828f4966a09d03dcfe9656a977ef6eafcf389dc3d271c86599a4089d46fce0642ed2344df3dc60ba46394;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4326e831216da34b9a1d2338524ff125c582bbf0aa86c05b0bfd618d605b7c8f48ac527e0b14d524b8d83f1cd25e9fd29fbcc569d671b74c4dd0194f687827e20b19b20e601c745cbbb714a724e5644dbd6c17682b7cb0988b56d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f685ff9bca16cb45449da98a87001ac60b81490b3e7f8a47fa22297cd1a74101f316770aa35f97075cbc29b6a7dc1ad541fd2efb787c77b7cf6c7050b711e21754438e5c4cab99cff9d1b3114826931e93ceac5bd46aa552f59f36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146914efaf2ef0d61684ba910de0ccf5803e44680e770345b98590462cb6147e93a33b90a38fa9f8703251c5fe5f394f2b86978e2a1680add1f514dc960e5eb3d532b29d6210715de5a9d5e65cd682b72608cc016a256ac8dffe9df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bff0dcbbb29218ba98882624d40ae69a2f72eef8b01236c128e06b30a2d9ff52ae916171dc4cbab791bc3090fac4978d6495a699c57a03515bc9ff12dc4588de7d6d5c54f030b228b6d9940f7486502c145aded4312b7c4dd9506;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4e5e026678fa5ba1280287e76fe808f1769abcc9dbf76790560d69264a9d7523519d39c21c3518d14e6f519e2bf358cf223cffbd77ac29e0db3ac41c0cc41e19c99300e8bf29e5154f7653ee2bb2c25a9eab45392b93a88670a27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2b41aee0851b59aa86a2a613c8f105a2d8d0081ce919a5b276fafd8401ebbd83c58e89ce3b91e6fed4a9e64553d2e125708b483b889d2b46b111384bb5e0d88bd0d94db51fb037bf8fb3ec134548dccc5062f7001fd71337630b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8b4a08bd5c4130f909ebef57e9388ef1e6d9dd85472bf6f7bd582fc86e67c1ff71bba43424a4dd1b86b94dbb25453fd6208543fab056e2a5a6be6b46b2ecb080608227fef3a963e6bcbcdce111219cc7cb24e50b5112149a5b7b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1230c4d1c62ae642f9ca55e26e4bbd4f89c0d71cda952958f15cc1141db28be2972a251b4da495cd61aeb1073d01bf79a2dcc4956b0b399000df52bcc850edca295da3c5c5b50c5236204d5bb6b7f544376e7255450e60476dc47e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf1c9622171905b4ea68d746b2115847259cc0ea669dbd22e536e40ca2e17f2e58ed08431919c9622b3a6eb747e259472412b8e5bc55c80a8d964826eb0e733a2b6469e57be49462c465ede7aee98b1026bcfaa3a3ebf01364b24d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba2fa5f5f9cea5987444eebbdee8a903073c3ef001ad72df073dbf2e864f5b6ef6a8136f4b20226294b19dfaf2902c8ade1bde82acf2b6ec03c0d65fdf3d34fa91350e55bfc4153ae9aa7833365b8961e55c63c95afd681bb7809;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a33c67f09d2366e1437594dc7f505f1cea51d042840055e807e29678ca41382fa4a6c89bb56e4bf95099a1ffcb8f5f446b7b2f4e1e9fe2aaf15bc0314c7c2e13652f5fd2e1c233acc2c573e55e1d920ee6c3f10fc0750b47c9d9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3012f49bc15034eb5d818a2bf335a5d5a6a8b2ccc9bbb52d1ff42c37278debb61182a55a37a854b4ae9679e38f3d3faf0cbd249fd2ca9cbd1460af014f380ff2a3178e063524f41728d2b99b1b989264c256503075b258b224bfd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbabaff913e6b0b46f3b4579df50d963e528e7385c949d31c515d98f02d3c9d1c7a3b8ff926429e304f9b67b614a88665248b602a80d1b723e0c6187ce60bd366d6bc8f4161c4409e14e488b69fa6bd06bf6cc0cae839a182f527d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2ba4ee5095a1d2c69211b4e2975ef043a8348bbd1193f15b12bd578858bcb6144e3d085b19344cfaeff94fb7911e53ee135078c58857674815d647e891a3e64ad1d57789667f422a4f181279fe9e22d3b38086d99bc342b2c422;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d358af3bb136535530a838878e51113e156ef5ce7a6765e9636a2f4f01506c444046768a710bc9ad6badf0d0c22e4704cfc63f2bba0b1800559212632f3d005f94242f313a1ef7dff7459b90bef59f187a6bede3cfa04682eb0079;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d00ce8e40124a0b872f4689f940a8bb4102d7695f7d511850fc0e5a2325f1ed9071bfb03c90fda9ba8ace95575d2d8109cdb3396b60a8c849807a40b18638ad533718ee7b05ad7e57d618b90dc9b7e6a56961fa0f634c7d184191;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1026e31c083b89f271a3f2bdcae3f9ac4b3ecfab5a7014a48918c594bfa40d23b52c2f801ddc8ab29c5da198c8b1aff76a9a2d64032e90ee7385f9670be9431af1655e1b98e20a8e0bf584510074d47f0d2b4223f275f8fcb2f2d56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h394cfbff5fc0844e568de01f9637905510b467732bbcb75231869b35894546203fca6b127e90c86b21a79ada4d174d048ca0ffcda685d27f812dc005537a7a6c25b9d6c8a1c86b1ca19590c3929fa8ccf01b6c7b9cb4e0c15a4711;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d40a3a5e382f394ebdf9d6e6b7763c2c12de1efeaecb896449fc4a56ba73dca42ae9f24c22001f7268cf3c946f7d632a7d30d2f5e1c63f85f2289f745e92add52c19db7e1c59282407bf73e3de0e4e37d9b1cf0752788e58bfe23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d04731220d60ff4ced41ff628086f471fa50a382a73d5a3e89c8d2828fe1db9370a5fb8730aba0e591ab1be3fd2452ffb7556947478d5b924d09f64d501d57e3e77ee08dd9d0e191f9d3ed1796bc9411f25b5666fd15e1ca1113f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99f84d25ee0c7d504928c8e533778d134431e12713b7fa8cfd0cdcc616630bcc6925ddf3254cb997faad47132174b5c49a3928beadd200e25011c6beae10f1e252a9e71baa4ed3994cc4a3ced45a040d50f1a1f2288aa2af16b33d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199f371f07b1dcd21674978ffb6480ebf8494e1ee85f3ed6d7c85114dfde3534de865a3e5057bb9df46d396c8b71638f6cb359620b33cef757719aeec5d3064b7dfdb104138561d62cd5e6da8aaee0724cb8d85360099c4177c2b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54a8a3b336572e7e8094ca8bf2f28e5ada6b0f1096e37de90baa38b43273d35be1fc4e1f81f6b6feddb2723dc56606ac400dd384db8a93431bcc14ecc2b88c72135830d3d5cf92d264484b94ae6f35421727602ab112bfa12f0881;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a41fa73a27a903a903dfc78511ca73a62eda62c240555441fa1dfe763b5d1afc60a8ebe85ab6ff0447e0b64073c928d82310f791fea10df32e493d6415dbeb5bf2e3f7a1f6f00a69bb76bdef9f429384f16fa2253f56c704a3e7fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd1cde7e962dd72af2f603df717fe1592d297fd6fd6529602b1dc07e1214eea329c19921b530ece8012956e79dbc2128357029b53dfc4fd43c1d5d64460870bd4740a9ecb8d4638bbf33a34e2925def873ca54914d26d54162124c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48e984ee201b8b28eebd1bcf2e2d5d96497563c90115fcbe5d5396462b091d90af1b1de727dcf4296eaa57590ab1a75489cb8418db42e1913431e4a99e210b183f43c46df95091310d4a73ad69c2e3152957822f4450bc7558e651;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18776271bfe42d69cd1104c48d4252a426838a5c40762e088a8418851c9228a75e6171e7fedcfc245bbcfa667fc89f60cf588d6fe87aa6a0a224b16774f16eb130dcaf83328843c8ad370c0f336fcf539f14885366763b8dc919f2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5de1a7d2654cbbce174ac873db5e19aa767313dcf4b0a84d07e9335a09248abbdba4533760d1e55b2e71ad616b79dc2abcfbef09136c4291281c8904f5b90b9663c4c910204a12ae7b6ddff6545230a29d8caab451bd5d1441a87f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118a4b7e57c3e668197b8b68678186a24d6dd7c1a88342536aeec7c3b7dae33b1d4172ac14ab6d485020c0b236f241bd8e921f0b9d0a5ad59df38087d1747927909e9446053515f71031c7126b865d4d4e6e58a4cba35058ac17d50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ec8cede15e8c2324ed3a9c073690fceb49245b391d06a14490beea0dc0e5c5d184cdd960af802f3c9a5546dd0a2a4df8471d9222bdb5aafbf30fe79a44d74314b3a40b80d11c2639c72f64b9dffa6243690141882f38c16d4107c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a08d717d9e8142091619af349d31c8ed99f7412e324ccf70a0843a261f4371c1febbce0b05474b569d64b2167e5c6d8010ab3e5f81ce9140e043694d2b1e398dc2c9436986c0aead293d1d7154b50ae3964b0d3306112db924408f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7d042dd394bb76fe3121b10ebea9a7902dc1dcb7014c7f465913820d4bd10e20bf08626b64e377454b55d8d3ddc278b4d7001f9d9bd9b93ce28398d458c0998735ce46b29f3fe6733545b2d93ab20bdd86b09e8e67fecac5253b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed52d011878ece48932738aaa733bdcd32a81ce59dd9ee6287bdca032caa09d7e70ef9cbc94d89d1da81408d39c1a6d10f9509c1daa6af97c4c191b11a5b1162d1db24ae314294f92eda6b20659bac0d365a4beb2593dc2f29021d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ba835a5eb1c616df28d79f3a7a884cf2a33d6b1925cec1ae9221e4a3892b0fe034cab3fa0dc3049a2c00f52f0abae2b2c094cb730f0004b3833330ca7060892de033a6899831910238436200b99c4044a9cda5dae0304554bedd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e0d4ead187f1a830f4796caf65714ba8be2709641c10314e356502ae62927e177f18697467ac7049051b753fb09cc9445f1337f33b53054bd6b9cd621a53d8e45324103deeb9fc5277ec2a48559cba1a3e895392e4b10a3770429;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1773b7e8ce1a68f88a36d5a9abb543e67c5753f336983e3ae90b0c7b213d35870fc8ceb13c7ab971920ae9c909cb4cc30ef4389f51da95febc199657b07dc4be99f9e5796700a7ed72c31504276e94b3cc9d6d9d4fe2c65cc636e21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1954a3ad08d1b7b5c055a6ef7dfcce0d3c61b49a5b10a862cf5d73fdda506cd7ceabcf9b3e8d195df2da6df9275ef252027d331255878fef7397b5e295fda0012957265a92d633def7b7e528584ef9f7139bed0303aabc92a08c5d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a40ac7e0dea81d52f3b4f05e78253684b41c7c4b7b0b2f41953cfcd65b84d1735fffd8665eb925642c1eec9a552edb271bee6bbe7f64158a7f7f4cf3a67fa54874f6a36d78f554c53832157accfd0e3820097d302b961db3afb33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ea7160d0e6051ed29ccc0d876b758fc3cfea906f66863f0a8226c3c9bdee1111c6081be8380792e2b679bf9e0679a337b31311209384bebd62a385f884a9f4e482a53bf6e73274c392874e6e77b96836180ca160e658118e29034;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c62e6ce53cd04b1025cab3429fa787f62f5bf9896395a17516bdfca1b048ac8d230117b2cca4da01be00af877532d23a2071d8f033131b893d9039f991bc815d3836c52deaf6ba612aa7e9d8c3a21ac7bc42409774ac2a8c96851;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9b3de24e8d1b5f23007c6424599e038c009604d37f8e41be2d2980ea5e7b65600e0b7d4c89cfacf4cd1bf691105286295fb057a35dcc07b752d271c771df6d1878b219c42e78a68007ca616a17b12279f1e4ffcb85a1018e48d1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1781e96660395a28153b5185269aaf2f57cadfa3fd106e343eaa558540f475cbbb40b1b9d71c14caeeee38e5ac6dc9d49e5a6fd36a6cb2328ca1c38da2693eec101fa6037d94df378c362b639135c0067bf905194ae552a1742d0b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e711c1924c764574cfdccac9b9fdef3926b9f528c779d636a6cc41a6537c8c77cd2527c81e8d60a02cb41ba1ead4f20003e06968294877e0699baedc628062e1e9b220ba8ce1e0ff43705cfc30bdbd623d177fbfa12cad0b295529;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb0ab36805c389effc183a927d1dc41e420e3f6173f052400c8b299c178f971d3e57120956f1729f234521b17726acb431c3251109650aca7469ab72242ac08076d57686eeee32045ca9e882b1ce85cec41c9d86627bbfb861d045;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ae09fc880dafa898072a19d5de01779296d2b93113f826655b7deab721d350d2935c72e45e8e123752e216b62f491d2479aef0341727bb0aaf71a669fa7fcfbacdab60e660db540f3c553d02de18bc4d349a1d1ae5474c0176387;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf3ccb753fc319eb086f64cb4492ba803e4571b09256cc700184d519f3c707e1eb80443baf4e1b8dcf5ce5a36d10ab859ea604bb6369007d07de91553a2dfc38bbc8d462ec765ee7e6064ea0f50c2713da229aae6da3958a1143a44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10496500832c6be0b818de53b41ea5bda6acb3eaf9ff9db516f200cdab4533e2f6c86177678bad78ba13d9220eeeca0d567e32747a79f672decae1400e1e2b47cbfa47380e0ec365f47bcea409d41fb1e9fc584506195a39901a29a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0f9a8f4b978dfc20bad7b788cbf5bf0370df4898448d0e3e8fb0beb026889c0c127ff2d0e51f8624debcb7b5e9550d2f9a13067167b2cb56523a435f417118e43a404aa681b710b7c54f47cc7b3bd3dd17b2edfc4e411b9b113f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1530d4ea8c310737d30b8dbee4f8a4f2cc036d1f0f9d6323bd47d3093a19d94ccef30c69fc71bb8dd854d65b2cb5cc7fd5769fad664300e591ca00f16b0ff2cc1e9734ff38519b56bc78547beb66368655159faaddd31f0fd815d6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb06ad2368ff5bb7d53171f0e1c43e84129b6fe3838482ac70cd518a17f37c40be428a5fd0fb85456783d29c8c0e808bf13639acffcca34721b93bfe3a8f3067026075183d42a10bcf3a13f9bd362551282cf4bf28c8b6cd684acfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152f2f5f03986ca3d55f2c883e7d5b25a6ef59463ded0736762fbccd516f2aed7cd9edfa8585cab5bfbd74dbe0297b90f08c5df0c4905166eb27739109f0d7ee404d1f7fc8202aea1aeab2253146fe04b1011a0f2c147d322d893dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c4d8bd0c607980a357af9c1de084d56f11a8e44b63c541d24cbff57c0a6222b7e81b96dda380643a7b7857445d0e03ab573275e51791cc9a89c072f82e777ed96387f727776f7728e521614581e0e49ad20aa2818910bb7275e22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100666f808d591991647b3c24146826fa339bbb14fd3a389251bf742396905cf1847641d9fcdf80a205be2fd83f6af49beefa0bc3740619c4b27983ec6d03fa7b21e70421390a2ef74fb2c68a0635c08b1fd5563724f1251f681a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c7923d04f0e32320333cf26112234b90f1db10fc7b299fb6ca81e5271e4cdf6a3e9c438096be19a21fe24a8555b24bcd2644cc5bb4a274ece852b43949a8c3731e073c7a9360486e3eb9420f923e7a293bd0e9b026c86d9a5c8c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b54b6706172639d4db1cff64306ccd993fab4e7f15b96d7e8b2990c563175355fed1b2740cd86572f8ef57fe636827d7bf2a6d4f7eba6d1ed1ef5fc317568f86bd495708e75afbb9a9c464dc620400ac00f95edd1bf0df7bb750fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a1d7cc9d78e2221f0074d1d3ad67ca5ae014c4b0536f1c53fd2874516c28423399b712ad6f402d739e267dfec72ddeea5b5177adfa9fceb8806210fc3b366f34b1c4237afb2d0ed8901103de2531bd656b9d6aa7486097b234815;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ccd6c4a7359eba9edd677d8fb9bef47b7d69a6717fda0700a189409c92e2584f79441b95824c79b820f4dec443db0b3279c6f9b8b93de9d6905c30282cdb77bddc3afc44ae30a61bbff44e2d52c609936eea6445044a0a1d6867a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164b19f6d7cbf847f9e548e735998576935f9b89ee0af052f5bfbcb3bbb118f4c9f976a893977c097fa497814ea6ef82eb748c6823279cd149ecaa3ca50689a9b3001fbd6da448fb3e39ef995f3f7fc94f75070833973ea7baa7434;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6fca24775774d447f0192256338c3625c2f872819029a781fcbf60a9153448a51bc6a0ce4296b067e4649bf9821a150ef1a3c8d832f2d2e782c443443480157ef12b06eb6eb24a75bbab5938e156fb16db5d5da0656679c48c68cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca949854139e5c9302b0860dd1b46e69b386d098dc3723b2da6f90e0667195116e495e3ac5957b562e2dee2a09992ae4299a155df6ae32753a472c4cfef64124e3a318d18a64c8de36a76d0d528fa01294e11902c7dd4455c14539;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd59dc4c48715983272770c57a68a8737916424bbd06d23df49b901d9b0b327f39b0dddd493b40885f90b539b9cbe97d2c3d767872998a06ba276facbe26e2551a71937fef94048de57bd22b5193dc59b8726d19788ffabd321ca9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he938ceee2842854c45a941274116b5d63b079a54c2583e2a9d103efda91164b9eaedc6ae3816a1eaf8c6e37564cbf66cc599eea535b13bbc62f08609b68be9d527828e5019151e5842b21fafec500df6ee7c57c02db3e404e50ca8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4a509a5d47ee5921f648942010f6530ccc47107a3320340fe1513924436c42026789ad44bda518123ad420ba1ba450c33406f863dac010bc76f7f8e43fca3d8ca1641b20385f10fbdca451c4c239104609cbcca82ba0f58f80b0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7dd0c979048d331ed3c13c349b1d01469d3837089b28f6282e4fce4d8f810e4cc78dbabbc000a56fa3c9f9f6acd0b5b9ae4c0f6ede0fd7e9bebae543cd9f7bf91546807e9070e9dd48b3bfa52d6158048c6be99802366d88753538;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c64d370ebb08c46f4315ff9017eb1ba80e410078e2c22d0228da0ba7475525526a50f98eb44f5fe1a08aaabe581b331e4d71377c8b8e310a560befd673f8bb073ea7a387b37ba866e8a4c8c9c1d95b96db7fddd24fea13b353b6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e6fc5d5f863a3fde79813bbbd52b87531032125eb76ca271339cac083a8ae96fc4ebf12ae05033c8414cec41b99b690249a802d08b3f64bb8350f14cd17d680725c82095ea97e942b90a6c10a4d54d51d64417193e68212c71e91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c0d679e44d9d9da0ff8ca0385178e463706704ed24e7323586f4d68633d9f4a14b262f07dbb8ef1bf6ebd5ac416552d781b6aecf2f3bcb83bf42b94be5f4627b73000ba40ae2cbd3e9bda6171b618f4f5f1ea25f385b8d7e0e3b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h66a24544215b4d003f539e14037981a504677da8941b5d22fa3eb6ddf700e3e61ad1dc2b2edf26de8ba9f33254cefe530c3c544cd0eda2a9fe6c73fb4708696d97f64535cf44b9ef377fa38a90baf3c3aa5f4850beaf2efda3a263;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7bc4c52434e74a14ed987d53eeff1be5070e446f4299be97732c5a8c26474c99bca424da7e6e5939fe53bfd0467607369a156a9d25e1effac779d155fa00460495b1b39755257682c7edf3def012386bf880aad5e9d025b975421c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52e5feb0ae8d5a11876c18a3d675cde12b90abe30a306a7433ae5efee07046fc3e5e83eccd1ba0eaa05bd54cc160bed81e4286a5bfae82580cdbf973df32126832e5962f8d37f9b92a0e5c06762875e45ae707ff0474881b96c618;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d0a866bb1c467b06de0a1fb88ec10e1193b97bf827dbbffe5916bf8e282e46cf0ab3e5972273807f23d7e548c5423d0ce5e0a794c815750bb95e2f5b78d28e9c2a6586679bdb9f42117a8e65bdc5e33f70a60fd89d4fcb6ac57fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172808c43e39f914f4a6774ccf85853994dec78032c105ad5fe4498edbbf52aa14a4e4199e956ace9f423e0c184e4dc753335c2fef92fb2e2b8410001426b37a800281e83a916b58c6c35c9342a0d52766e24236f0ac350ddbdd12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1146cc5321cbbfe22bc1ba85b11c42e2b39aa1100789862cfd108eff705f76431ed327b32cfc8e6edb3dd7687ebe0ae4146192c1ff476fc796bb226078cca6592aad0d213d475817602647bfe88e201a1444b1f76ba0e2041daea6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af9ed4e6d15028b14f9f01f3dc0cf7f190179259d258c4ade7a47018cbe9ec41d9824e715c775abc7e765c0bc2546ec967c05deca2c8fdf5ab085425ecc8fde3b362a86b7b04324c5387899a83e2217c3d8d983b9622bdb2ea64c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134d5d9a1f7a759f57d21b19af5bddc24be08fd7089cf41edbfc6fd582925bfd35278af91d60b0099dbaf08721850e4fab3f1125b25063df2e64e3f343ebdff0c856d47f2f47d703c0812d59a7998509cee25f73fc689eea05c5924;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be9ba0f0cc07fcade214a8eac8638954a290202f1e1922cdbfa499e446230d0ad188e261df93bfe385baf56a90fe312c2f283fc1652ce70d8719711f79a6f136092494b0aa3e0cbf5867379de819173e7c83e3ce76e62ab63e5a6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4773e6571d18068f2b0de08ceca96cf1fa94166479170d828c977fae4b3ae8a83044d46ea75965163d53c474df52553227fbcce7c4ae2ac3b52e361ec0e9fe83c0c887257061d23fb54fbacc78dd2415ed0af20c635aa6f4e9b1cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12275c146d514fe7a2a14b31fd604746cdfb49dc358dc92c7d011c52fa5ca893a785998bd3819745766bd437efb4d7c450d05e0bbbe96274f008811408acc198911c29bf572774217c7c787b1e9b4c461b7690867ddefd68b5b9fdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a700b362526798b4308704acdaec8903e40f515e8f5ff2cb40173980506ff9f674a5dfbfd3923c401a217f19f916e8437f7097b9fe1559a6346edf4cd8ce68fa0abd6eff4580827ef9de8a05612b1a45372945b7a4f4fefb38cb9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2a8679b41d45cd6c74c4b7b4795ea0f681ef70d669b273e75edace907ae1ff5a422fc5c79b5a0e0c91e5476d2f940a88968024fec2afd459da3f5243901ed1403503244ed3d738abc31e4014d2742df7da14c6cb6de2ec060b106;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1508283f10cfed3550c5ef7b2b3e96063023f2f596bb77c4d5d0490009e48c562ee65a6be242f4f8682c2e39c685190bd10f153748a1ea84a8a30635e9430081bb6be4e00014ccb80273b363238263134d0ac228fe74d9433b54e02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eabee803f0e97acd6b9b7b2e62d94330d5fbf980ae51150641ab1a7c4dd9670c434b9a99123acb58fdec21264b5ff6ff1bd9a21227fdba1b96c5ad24134123098a6272f880186c134b1fbcf9729f9b763f78fa0e7752b8cb52fe0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a42ceae7696ee4660be7096de925a747c51945c23d23d5684d04831691ad46a9aebe2377d4048bd5f2fbc1e02507aed9ab772ad749644ea75b75f19c36ccd28b1d6dfc7110a5ef3cf08a6d5ae0a5275bf58e9063aa2722244a7fff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a527a4b8bae97386178594e117b2e26d3fa4574d8f51fe02928f86e6e2cfa6294c77970d58a6c422b26042dcf1a82bbe93ef2bdff5c373742c7601ee1de10f9bd6ca5c2ea8b87271f39460a98fb514232614ab03a13a8a5ca46b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9413c0d1969741fa0a1416af72e632069f81a690f20ae0b018b76866528536450c00152a71e662789aa733a7601ae78f69567b417e377a2607841e6d103a5b16d726f4c84c6281cd6af73274d19f63524e00622a6b1d0993b29186;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18771295c8c79ff5c778bac5dd82dd8dd847d71cbcd9c9602225030635d930990ec73a1d6d86bfcd7cfbb5cf5c00feac58fa4dd8b0bdbe4d6e4c157eb3dc67dd796dd638659d17694b1e53fa7486806140155314b8ebea7f62196cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efa6c5f59480e3fd93b0195d479c3434d6f3003b6bbd1586c717c5b682775feb698211f9e24b2be92ecb9420bf5f83c3599863a00402c0ed28832d3c1ea5687a90998a611594deb24c5c4aeb9eba5024258b99aebb82f2bc6077d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h236523703aa39d74267158b2f9fd6f6ef17bd7e5eed8d6fc9d8d226e587e9bc785838ec8f5352e21a59c1056f1ae729a6bada68a2db39745b81641cd948ccc182bdd87c4d66fb25299a7c6f05f055b0f63f2b1b636ec6066ea4fd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11db33f00d4bda5989f5270e7242c26a19cf7c61c6ddb2cedf19cec8e8db76409729a6a9d6f27ee739d2f21101946095fedfb1f4671f40eed9d3a211ca46bb785213067071c9ab4d5904eab38f4fd87008dac39bad5ac8711201d72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae298edb520e591303c59943702f75d7c9bb18716e9021eb6174607ecd50f75fc72d5bcadea12ed00f2ece27245db4f7850d3f29ab8a0a690be2c320d830bc8b1f594714da3cd0f9095001d3b86a567afa6c5c29971a4ebf8248fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ac1b64fad44fbd5838bfcbdf0457bac3c4e07edf9561de6f9256dd63c2bb63f54aa26fe26986ace04855e66d223d764201854ee3dcc7d3e0e7d8ac6ffd0c386ce7e7dd184a5b2de9405563dfcfafbdcbc9ea01c3babc862167ada;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174ac92d0cac822f209e10f9216ff04ed933129f073fec64ff73f54c582a6677d6f687055630341dbee48e60b491b7bd0446a779743bb54676237dc31e9fe95cfb04c44aa8bacd02494fcd668d1b2a0ba8cabbee0fc3497ac002c47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1e039a32b0fc679f23ae9131ab2fefdb54352358a63a7b4107c09fde48a6bf4a5351a1fc6c1f2831b7e26ff5cf4a662c3a5c1e45492f1ebea0fadf8f0f0b1ab4ab509b20bd5db1ca476899683615973146443fb0d245ce11de70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ce14a202c977090ce5ea525f5e966748b73c3106d579b1ce386960e94a1e35e2c1e26fb12f7fed64e2d7e8bfce10415c0e4a0f393374c70cf78f6cbeb701f0dcff0052c808b851836c2bc8b2c4ac9ee48ffe43abc2b23d08948ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e197d5f38b5c7acc8f8d922877a732064ac1c3e00b87afd8e990a79f0199d0699e6f4fe12e70865b86d20d4b286ccc7cbf91f184d95a231972569f9f22db4c0e1821b9e68bc3bc626d32493497c591681f9124acbe8ba0489b517;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51f64d137805fe44253f7edaa7d272c0c218db1305a1af0e4fe9209760bb91c561d9e648afa5fe3c5caae1385b92fdada20afca7fd555af3ec6e782f598d6af4041b2e165428d442c049520444176cb8aa64dc18a591c9aeddff3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c9bda038d0befced57a4ab880c876e8e3ed8db787a5d5e17d6a0c21c84d6b1ea178958a6b00dea875438b756cff35fda872eae088965057b2f7aefc1ce9f3de4ab6277987bf788044393bfcae07c6316f1f6a134dcc79df10870;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb13e8286cc26d4e1e1e0b3dc1bcc306407b28821f31a12ef940ef47af562fb1e34af13c259ec3029eb3072d1eaaa5f9f398629064634a5c795e964b6f6c491d029ffef990f1d2a6961eee3bff428031af1d3ed375c662c8ae7d7cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104b546ddbca490251a73a106ed729d26a2d4174814ddb064ee3a8bf7f0ddce85e60b24254025852e9a2f376f3cece1e66961503b3ea6339ba3276815fc90b2e6b5e88274d3a45f95c20c209d4412c33c03d234c39aa564a0d190d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cd0ac6946b3e2c541f0c71199251afda9cb1a44e5b8315b6968e4a719629deee92f57ef79c672ceb86123229277fac7943aca275c0d002d09986321e01583649c0882eae8f20a21158aa65e8fb4230123fd1b01f01790c7d1d1e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f9666c29ebc0d4193633191b7a71d26b9ef0d40f05e2d75c657b08783b2ff7d9a687af45f9a78a7c414f88c3c9e779b1229a113ae01c2c344907b7e0e1f83b6fa91c8ec23a1810ceff29358351eae3437a6b0daab12f153c2a426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb28d25b6c4c7949b3cfaa3843dfc5718618a7a330e0d9e67d9be05bd0d7f5526b41e4fbb006e8fcf98ba440f2529f5775f9687a45aacc5ec5c2925a208e5ea2861a48d4949f3eac8a0d1508976419e3e6b6718b595c2797e23d55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1179f853a42fa7246ce89d7a43535a7c455727c651c2bcda622a3f90b26c47207668dc053f3e94b0987308851a97d6661a8df74c1683e7b1e289a9547d0fbb45ef7ec900c0d75003af344ec24ffe49ee601d2706b814245ed2093f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11356d52f70e579d93e87ace49b77f6b39955d675e58c69edf31eef516e4e2e914a74aff4eb3af977b30d0bb440e53ed48933a5b7bd9a79e4d033c46c278cffa996e499cff738bc39cf5fe42eb10140015129d8bb492f624ade7255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f6b66cfbe72f6bba4756b47499861fea55b2bbae4a0ae5d4d1a2a9ebe4d2ea21e9477077695415ab1e7a952d3debd0c7957e0ffa5ff1d88dbe042d4ebbf4e70f4f57951aa57393fe547fe6d55d7d43bc3431ddfa9dc478c04008d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a8e78d0f6db18b98b7a13e6d8ada775ed10905fb592005692b5d7198f749094f3258ec360d7fcd789e36333431d860f7a39095ba8078560c6b8cb3dc888018e28ad4f9a430313121063ceed6e1169f415234437138a55cd8ee979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86f9268994a1df71576c3084bb077cae6776da11cb5ed9fee7dffab8ce2d38298b0c4f52ab7cd30604f7d8d10f297e4700dca6b4ee5d632d15bb617decfb8e56a48580518a9cef0a8b4f74c88680adc2b5cc28cad171d37ab7534e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fbb929946b3a9adb2f89e74a160a3beb6e3f8a40de102a55670227041089e6ede6f5f81fa41a7db336349bed3fbb8323be3adb0b19280f00a71d622579fc6b8414174b770a1db67cc113851b211a3e31d627386a9178454543541;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha44c86b15e287ad7303a2910f55d0de0a4bf19c3b5fb9ecd8cfced8eb51a1a200f43e7cd7c29131079cdce17b628b3c0c1a98a00081522ecafe538a4bbb54f43f92993008db63861a8c748fefb0c9b576778ac6c0708a0547dd8b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c6b666a2bad9ed0896e4d639482f2536ee9514166bd5591c99bf6916da08e4ac586681f0804da0ead0c7785f7e67dd8def3d287eb726eb155232198f395b03a3adf3b7f39eaa502fc7062953bc42de1356efe53b374ee31b6eb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156ef02a76a22a6e2c741ed5ae9b74a47966f197497a81dfdb1036c496acdd666cb78c4756b7d59dc149961a314448a6ef5b3a6615faff33645510b7a1bdd94854a5bc8019241dd3cc88be2f0d2e48f4c997862ae48e25cb5d78e3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47cd0b037521c7fc77a1c756e243faac5ae5c3c814cb1b7de5bc1cbe1f7c357a9037b65e4ccc7d5bd26b2e9c60f4d14e53f73732706530bb5b7ae40f3075fc19952fce2f964c532b9e7f2371b52ce5ac6d485c51cdc55b3e764616;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6282db1514675a64e8805257f399216915e866f937eb471c450c3d4a2931d72ecfd427a3de32caf2d328af160843ef54a1b277029c78bd1adcb710243a78ce482c3586ae16130d77c0e29d2c32842f030bf4f98ea54108f1a44e12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f5cb2665bb143ab39a54b50e39d5d1ed0f19d90f9794898e0baa21ae61c91d0a4519f8abfe4e54dbd2ac86e8cd4ce667b673d5a2ac11c6d7fd38b8340c94e8ae60858b6fbba0493d0261c39fbc8a5bffe285b0d086266d3906096;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17be640b71f2ea1e60a8e1d09a33ad3beadac804bfc99fd8d6aeaa88937b9da657640d7cfffb65dff3fcbdee921d14ae9de5bb91642d68900f48fc34df69ebeb31466f925e721df2ab491a68ef7c26a5ad3c12a06b3ff6da4b2ddcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18985ab4e48df0ca490da8c1e918f2f97d79bd24724ec2206c050054bef2324d900903fc1f792f868330e0dc6945d7461cd9e8a929185f7bb0116257739058e2557fb4b5d5caefb7cf9d953b7ac4d1b0b7287e6ad6f149f1dfd965b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1077a4d7e334ce4b4f73730e6a236bea576cc36d458aff6bba9adac287d34c201aa7058201b4faa8799cd8fbf3d6726243eda7cbe484151eef9eb1fc88c3f0183bff6a6b40f1a654a291decd517285c482624ea2058a5e529f07e9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h624d1e01871ebf0501d05a0ca9d6a34a3588b1d6e76b7ce635b7d9fc37ec751d8f0d10cc54638cc17e32f36dece5f103864b291cf59b7b62b67b2f322165f9cba83b0c76d4e9690544c38ee1257a133c9bc9c96237252d96a541b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c33f874fccf0a1ca8ac0f029f3fd4e6ab28bac4e161b41605ad384278c7e12b547956fcb6b8647e339f5a5b54fd3a29a55b2abfcd1cbf4daba0f55658589be464e20235b14e669fe4821f954a4c7a5d1c4554d8da3167485be0f88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1523e63f7861e3695ca72c580978967b9989f0de1584c455ee2cfa8c17d2e6dc8cb39f16fa91600d07847479c24007e41b8f3d48d26064a0f01e8d1246434d3695ba51bf815e31c576c18fbe714a005b9964f417a387e2dceeac4b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd29e64399e00aa46533f69329cdecbdf3c4e38d1cca43c29495857fb5d2f70dc4544624c5204b8ae528479bdf6025d26db2a9ddf0c9b5d6fb73083e36670009ecca83e5d7b3c13246a023138f12e739058d0c00b92305103d17c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1980a924a3c5fe4bc86545f46d8092bcc8f0bf44189628afc8c3edb2dea8ff6bee951784eec7f4665e54d6305c451ff42af706527a2a4816ff2a66fda56ab02827390677b0cbeb3e0aec573c983f979f7c02a417a491fa4225bf426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1038c2dd0f6e4f75239821d493d36bfcc6a78c035d5441fad480b9995a5d108097864ba10c8e115cfef9288d36c17964e86efc4d89c3182e385655f3fbe7023235e520acdd5ff2c048b92b4606c4e6b4ffbefd152d90fb459292005;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3eef2a1cd09a4920ba259bb0e426490cc3a5963ef0fad5332396deed23f724899b7da8e7b50dc2df403014c85ac78b5f9e465392ee41b763de9be0124f56338cac533b9cbe77b0b00f21474c062ddae2c315b0ace8d24ce03c05ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb58a0fb558e10dea8ecfd3953bea2ccfab30401ef9bb57ec693312ea87848a9509efcd90ffc92d1a0fbc05c278159eee474f17e12ff96f0b7ebfbfa3f32fa1bc107928e9d95de32d1d1a798ebca7ccb7e99e2843370409b6cca19b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba99ab825eec600c215545b577756de1b0226e65f774ccda5485135ada041b6e797cb788b1418ec96095cd13f6888cd8278329bc65eeb7f5570c57940bd84e31d5d5cf1d97e32d067e1d388461f58c2c5c816deb12182816ee12fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128b6cf31fc0e6f2723a032af2df8f34633b5b2997981605a8be95a076ae69a44b6b171a8f35d4e874fd76f4576945d81a707ed5d4b7e5c2e2cfa640153306f52d0b8869950fe0685b810545428c17fe82de70e3d5e4bc5449bb4a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c28e831a2f32b136df27d20fa0ebd7639e98ffe2bcac019703cd78e8f575ffe1c25799dcf8107277d3154be9df0f11684e7e92bef4253fc01bc57939ad56e838703be476f816b25002c118e9301377e0a3843438e3719a79254f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaf7fa41dd2667d2f676204a80a3fc69d70629ecaf9c1f96425ee3f685836cd960d1ff81d2cf8026178ec229f7815d8c78026387c51d2bcd53429f063fc1aebdc8fb68966657765d406b08ab34c90019d41a9824ff336c57c3ba41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0fb5be5e3e0d8808c06ff42100d55cc6a0754f3f3d9558d579b01a3b5978b55094e60177ff3029aebe9a633021b2f5e4523bdaccdb3ec7aee4daa39b7cb0bb1cd8dd3e02d69f116f48965c0d7850c2263778ba64ae94df8fb759a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d6acb9757f60574c0b2c6b107ed34b5eb71ae5f38cbad297e66f6ae832e3d7211bf41f267e6620bb6d07062275801d342622bf7f30131741e9f5b65e96e698eade97fbe4af45ca5f0d78186b7f22e590ef1f820d52d609b5ec90b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124c7fe942c4fd99a5e15be8b8d21f9fffc31cfa71d0c497e161c6548037f0984d9731312781849e43ef87c483daa0c28f7568bacfef24f0aab776fcbcfea0b79b1bee381a45d5387e8d23807b59d2b51e0d4b655a3011f56a13069;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7fa1bff9a1dfde6d6a56fa331c74cb8520733901d4e2c1aed083edd05b02d308d817e97a973ddab7299121fccf3f666ad3c0953b94f3ac978a58322ea6f24e165185239483b9252788ec949fe50e82e952ab84482393a6b0371762;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f77fbd80f63a9b237523d5b6eb76543c0adeee0fbf29c3c68c8ee68c80223403ccedf9023ae7587ef0973aa090be4fa0b46fbc90260912d07992bda084424b84c343e378df8c1d768d51cf7a9028b31eb829276a4b09468d946857;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87251e7499e6b1f26103e5374b56074788afc03aba30c68995b11aa1e39a6e29ec1e4b38cf87a7e3b956bc3676f6ab59398b358195821cae3ba7fd97a6ca62452aaa00c8bb934c6a83de8a37c9f824f29886efbbcb9486afbe655f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c42f713d37b01ed582702f8e60d85585717c4db3ead7a14cdd1924a9f319d92a809c49e051d556ec5731887ef5baf24d7de47d6b90d5177a21390f3025c3da9799398b5dc0b696838215368e94c0c32081d59d0ab2c9c31b7e62f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16497c82780640f5ba396997561e0dcf515b786d99d36d27863f11598bcf5f4560f6dbcb65e27632e296073633a35a65466e9a6e2894597a2b17dedd8add8b38cfd2302e10bd8f947e6d94054df92dcb5a098001b970b277ebe68a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c5e780702be294d39679ead3dd511d8e3ea613360072ffffcf1492fa5d30cd67272093010c24504bb76d9ddfddec5878b4a91fe803688493630fc7ef8d5509c89ed5cf8310eba83066696be24bcdb6fe038508d240e1ceae76794;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haae0171c9e686132edad5e2ee253873804083d15adbda4e192f36395ee62fc0f3373d632d100fbd96374b76f76f28a24c2109435c2910bac3753abc41160da3dfc4ab033a36cc5f2684917568312756918be26c4c000089eebaa4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d82bab3449d16352fdd549992e9229f9ab96cd2f403853b3412317271628a7535a83a0cac789f6f633881c0765462343640d2c816d0101a38497cacc2565402fe471eb8e59eb329eb49b9ef4192296cd77196ca590f603b50ee960;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c54e3ed26f5321920c6f95566e689177e5e60851e9fffb8ea621db3cdebcef4aea75ccf5666e31625da06ed386b01d2d10372040a18e6fccf66b7fd691c1156472e4fc871380040aaacf3e69cccd9efb9856ecd4e250d695c30d67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e469ef44cdd899ac7de38f60fb3f9a1d68652b29ba1bda1f518eb030dd87713fb3177b6f28356f7495d94f9f15423b4059820408fef8ed3d87903316e63a35a09086a2fbe1fe68ce0d42e47aabd5378e9c3be2f1272f138820e6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c84b4726eb9f959aa81d32db0887f0e0e16ed14758ee055e8ec3381fa2d1e5f2e6e2311d8aa6d2ce87a925d4f841708f8cb4648f90c90f6b62e324085f1cd1764100abf1d4f8d6b1d516d83a84e4409ce76f54a51ed36f5646888;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f83f7eaf43a229ddb42eadf7c1532fda67ad132a7524b99d8af3651a1b2f21a2c056753185a55907ec7d63196bff1c9a591416f668b5a2a9aef62ccbe09143461f6b5ffd61525aa4df35ee1065baea3aad87cf219104e0a60d8615;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cdb63a772fbeac96bebe4c5b6fd74de2481122d1e19f8b154ebb71466384d8db511941859543c44ab98c45cad2de92a801c922506bcf6f8807f08e16e0b1adfa7c6617cd0fc86a77067c396e6ea595d8f73baf049d48db784ac650;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h145173bb75419f9e19814cfc9805501c04b458470653aad00b014c8ee5f428e62fc19d4caa8c0b5f948bfd3d4b70579a1954cd1f719f8e821cfcc8e744b1149074ec08bdae0d7e81ae792b1640a996e7ecc47a527d1c0579462286;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bfc7dba10340b9aae4400a63ef11762ce0217ace2b5c42e344656089a259821cf437aa1af6fda6cd2a38f928bc9b37394ee38eaa6c0f2379d6ef2444c59312c7ac155347a41de33e44ec4cb830d679ee0459a321fce67e5e56826;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2131883f11f27bdbb3fe696200326957034715155bd8c2d57e47d1604d10fb1b5df422a4ce3075b28757dee1dcef8c415c72a4ee4eb5bdf4f2e29efec4004281ff2901fdd846b2375e39b3705317bcab055d246ed9aff0366fd17c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he230983ce6ea035d35f6dcff0c167da729e57672dbdd24e18772b7fb3288f44465075777c8b83d1b90f04fee9baecad6ad7434d5a1a575f137d0ca180e66f77efdd1597e651e760dbfdc8c8ba2493fdedef737bebe822ed7086bff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h599b28406f875c8f19b4cb43fc1c83868bd7f0ce7562866c4a707ee839885b93a1a4c84bde26f1da4bdc5b8988b783d165908ea09feb33c1de6bf1745d6ee56ead072c8e297047924d946043135689072becf8df8f5ec0d5c80f78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9588100e6baeabd5d01e98b610af2c40623752f57e5c1687d800bfbfa4044c8fdd033eca8d61af30ebc69455600d33c128d8dcba0b8717a0bc09bb17e38d6d80834a3690ffc3fc3cb1e694f70f74821102ff621fdf71549ec6e205;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7020e75d3e0139b9ea713b601e5d6cfa5f5596998837e2a6d5af4e23a8d91d8ed90c23bfc0ce9c47a076e21caf588952521e666e668fa7e753e0bfa2d616e161eb2ee797f02f1917e0c70d77875421239b44c1ec99da4017558b3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168b97ecad891bcd3e19283819cc7c57a8b97823e7d014eab2799ca7e6f750aab98ffa31f93463eec1ed93da2e6c4c7e70c1cdd2a5c728f03a4da9166e70e37b8ed5c3036441c2e99e9746a46bfd7118034e8850268e64f5dce1bea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a23141e0c7053653d5cc943c7cc88a6ad80fa051c9710911dab894b2af1e9fbc7783c242c8f3817a8093040d43e17b0bb854f71d847b70829445a626edd371436e4345bf23056bac28a2f1261ee51d0c53d32ef4e81fad263809a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fcc5f51a16c3fae4145beebd55739dde01df48a9874f11d3e04fee1b774830d1726b4686224d2e194eda9e6e2da479d0568fd0fcd778ffabe1c3afcb564f7740d35558212f45783b50994c2a37df5652eae2842701d87d0c0ad20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcab6b7f7a0e0d411612b574ae738d08a8f588fcd7e24f0e67bd217195ae384ebd0c235c1362989d1d41963b513a97f8a81668874e3c60be968b674abd0307dda0fc912bf9b5d50bbc0c667960cf337e24b2d3e9ecd7974429bfde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bfc0601a759008e58fcf56841e63ce29ed7696649a10c260ee4b9f3c847b0661ecc749a350bd3fe1dbe522d6449898b299bd4458902754946c5a2f2b0b1031b88f4bd13d6809523dbaead283a4256b1ad4cc27062062618316eebe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169d476ab96da7ef636a188b5ea9d7fd3913a81345e918210a74f57beec0ee592d7c75e317cb15507055154a0a211dd29d05425ed76fe47b79a3215f93505711374f7ca15d0914c8b93309139212bf2ebf8c7e990afcb04c1ee9e82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd73b1bafe7844d24bee8334fd4d59739d987da1655967dad3198f7fd0a8a144789129a2f7d34300e81d2a12be94348e27a879c6405b5160bef633a4c8b7c4d670d835cddcbb21e90c158fdf08808b7ae0e92b0753736746a077c60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ce89658fad65063e853ee495b6447f98988d50039a9e83d54717e3fcb17c804708cfbbe8c03d30842dc636e084de3c047440ebb69649a1d11b3ab47a0fa839eb136411e2ba802710ae13273b0db2cf14e5e17d592812640882668;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3286734cd756bd65ecf85b450b64676267515f509b7fbfa3776a4d61330cbc2ede823ee290482ddfcd690cbc94b5daf3ea4c61a76c14cb1277903e09fcfbd7077b90ae6dcbf2fadf421eaee4ea70bc95cac9117bd02406d04a5e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e36cbe44681774b2f2971980871cc8b4fe560239966d34298fb6c4271cc3fddc2e8748d51cd0d2f23c111ff21f763b9da649b56fa9903c7524cd778d480e81792705ffb2e4cf00adad8a233e83c619c477ac8113ea30b78343654d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d69e302d11a0256851084c1afb2a6307233c3e604947f75290f49920adb1d2479825d10bc213fa9d72c66b5b3adeb62c59f2713abab51027e582dc3bfe91587ba11cb6bf3f2af767ccdbc87d2d0f09aaf4fbb665a5803402236d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e22d249ee279a71a7fd35071be27529d9c95652b5676b053e6682d6612ebef133adc780ed5c7b898289b698f8469b35f918e9bf76886a31a3d2e57263bdb38453c0550e776d14fae6554a5b624ee2b12615233e520a742d3daaf9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa9bdd23c2338ee9ba0cad1a8c20dc49c92098e901590adb7a998ecbe615fd0860cc8784abdcb2df27e8c71e71f2dcbc86e2a62b0a043560c32dda974c3d54d81519c4688d87dc3170644337ff41e5f2f7701629a3de0fd12dfe75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c3b3d39a7fdcca07d8ca83ba55917c8e3d26a5b698d894286614e91a5f20d3a231c6cd6065fdcae76679c2e9a588a22003ff541978af56e132924be0c5ffb80c654a87acb48419addf070d51a7e4dba7b0b6917bf26fad0eae541;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e4f6a459e3dee087528be3bda8e2af431295cf1d7776fa72a7c33ac9c429f1dfaf05aaebb083849d040345cddf7a38e5ab8ebc87639b5dff7d79768e60566aa0195106e225554e58f8abd1fc911868d95a7f1bea875f27b40e4f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac7e05073032b43423e87d0b93ce04dd12a1361f6c6d43dc094170e4de58f20aeec8e364bd95eb31049dd01b2b77ef89fd585ac2b5365fa8e03353cbea5aed6031a11ae1ca2f757568d87fadff3c0e1e6f110493f775aa8e30e67a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5608fe9dd5f8098fda31a1788dee0e62c22f29874da096632f73518c5ea1b1e24c42c5f91d5152c3d95a5e04e453aa56da868cc88fa3ab3b5cc732d9e46853b58c0e44ce5f38e4cb5ca0db3f3181157f7afb82bd9ff877c0af452c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he64f5b1457853a9b956e566731f1e9e7faf40bf9795eab7999d2e63141e5063dbb1778ecb7f5cb557a611a94d1b65f067e191a7c9374f33182345d311d71fa1b9042aa0bd07020d5e2fb4ac236df256189e9fe5f7ed3e1846b3d3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4726eb139c843ec7516ca0f323e1bdd6b16f54798e415035307814180288bd217345d43fb277e92370f8d15bc657a6618babfd9806f4dac11c3990540b8ea9d3639a1dd70fad49dc9bb33e8c9c0178d4f023c760a88cf8ad1b4746;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144e71c112ea2aa7b9946e1583fc9fb09e35c22e9a9f10ebe33865925991a98b2afe93cb04bc5262a20e8f256f42bbeec0b8f059af65145a1bcc0ddd5081f51daa2c216d765ec465e05982f05920461803d46f9cb0e239709da5f61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dd2b4141cd3beebfbced060e9ee5e40e66393cdb710829f13c83d5b6547d78436f03f348e98dcfd553ba844a29fc8469ceff9c3f8e59f9a1f4c92bed683dd897aee3b22dda6d4ea51c603c011e0a67da753935a4524bfb07321f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b6a6efbdb90a4227cc3ea2876b84b85112ca2e7458151f28d7339de4c64bd2f4f54bec84bb8dc64b5335c91918d1952b262151ba6664bf88b4de2eeea4f7094353c9c172736abd8a0e7c9bd395188bd2344686d782f8048aababd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1957c71f39a5785ad057d27f2b8b78ef401776157ba0892b0450180d61fc42988b2fee03b22784200819d87de39be1375cd478f1157a08adeba78fb3b09d30796dc1b191935d0a2e21d56f42681d35b7ce4bf7a2fa2a0fa6226eadd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a8fdb92120c92f7d638301e48e2aca3ae34cfdcc72eef59e58e5d0356688d0c8d6ebb6e6ab8acbf0ec2d49b3ddd45f607ba3acf2c2c1c869bf8a8e900c20586baa3fc06a5bd5e8d1a25aa8bb42cab436039eaf46a0f08220ef33eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c31db964785b3784b5f9ada0267a6b9baecf797c1e9add68a66f56a58a537438a0e5430e15a5cbd1afdd172e6a14f2ba06b409485fe14e274863f057af1ea5b8c83af77ff2296dc5142c505cd06a49897a36bdb462379678c99a48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d8d86641bfb0e0cad44ef936cdcca9175fe34a6d49ef4cfe68c25ecb933fcee965708b42b455cf3a6895cff2bb4095f0d2b6766396b89612fc2536083b98726a83e83b27328e55a5e1945e3a57c949e160dbc89945186c470fbe7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf74a0d7675c3aaf46abab1190ff232493a16a808507799b9bd3e7cf23d81c1616f1dd131df8d3067b5d10e33a80bc15b551fc0f048fb76316efa45391ff9b76dfdcf6f56aba804c1af71d03a81508b6ed6b37ba6d19d1927b62963;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bc313879d053caf4b1df02ff35515d47f1884a60b1230c5c641b52c61e12794de8417d3b33ba34dc9f85c15d35d1068549bfbbf3eb1fd3f91d55125ea8be5fa61148206a0e5a3dfe02eb3d708924b83380bf613c00cece9b2f8ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48da7077240755477b8bfbdbfb0311604545069fef2844d24d61b661b2dae21728c26840c404ffab9e5fc58ac54fd1eb26f76302e66b766663fcbe99033ad69128966e79b5355f7515275af6c7a1979f7266e0aade683f7e812cc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7c51bbe0aea8ebbf04e6b75dbe258566671f2fd573630556667f7524950c7005260123c5405d2b1c87be0eb5a42b5453b350480015028e35967ee05ab6e8f8475eec5c6e7a8c8f42b0743aff7726bf5eec04412a97749f3e6af85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa39745ca251f1affeaf51e45a0b81ae724beb18fc6ddee7173fb2fe35be3b08de1d5e9bfa2484880bee1b082228fbb2709b69eb0051c40130eb2cf43d67c03f8f84e9504f879244b8f38f3d04ad0a9b797dc32444b44fbc4c17d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171e31d31dacf731acb294737f4ce7e3c623c5d4b5b3dc1e015e8bfd1fc3cdce18dc73f267f4e8348afcaadc0de2117d19e61835e0e85a3b6230b51f8632e8ce929d5029a26faf4e0142bc54fdb8b57d1723e2f218e2e1f0487a45d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e3f6915f69e9b4ccc40dcc11286c3fc9396f3b58e84beed2e25c237642b8a385e1dcc661017e8ee88975eb4fc3a84bb72e877478e5443d12a30e0e9d37984c1d6ca295153fd567db8ac27014b923024e95411117ca4c1a1a11264;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ab135b2b718842fec3e03468923c0ac0bbaedaade6b160d595b7365f4c48c3d3b6b969ed9bf90162a6f55bf8d081966cc4badd21252df3359f6235bd69bb01850d86bbb9ec754bc4f1b444e7f81ed9b5221a7ab93b445b7c0048b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fa9a8a896a00020d761a1cd6bb53d2fa1b1e3edd8d4fb0b0f8a060e4d6cfe27c756904e9b2afc7cff6ccaf42b355f2f3dcd1bee7265a7819df055c455a28bb214a7553579e8d8401dd6e2a4d336bc40ab643910e883dc2f9e6cef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153d34bdec7882f3d74555279a165e2448294b4181e37f722e939923a1b4f5f6eb8d9370be0ad7158d0a09ef472efedb98030b32e96cd598c891410982350ccab4071641ec76232efa949fc0a4ea676d74a22910a09ec85f31ef990;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157221e270d199ec754c486a1bd7efbc3d621786592728ff92ea2ae5084e9e884c75c7c45919519c8aa7fbed57cd8e574ad08dd02afb2c6be54dd2bd55d92043d46168895a22745936154ad6b8131e87a88aef5319e1fa8a7d072fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d329579981821846f85a85e17d701043934e0f5204d63b386c29ba627a64abfa17cf933b3656fa1a739a45ed4ab7f3be591e69133af687b34127fb9c378763e617df3afb6879ee86364d79c16b49ae1abf5c3f724d55408741b58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ceec6764bffb6237f70672ec15066d9aab69d08af5bbe3d83db0a9ec3ca132d570580858ed878627d3920bd26c99452b437b73ea49c1be1e9e278e9c5a27ccdddc3f29d8525cc5524c73da9e2474af6f4858df3d5dce7498a11db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1100504a3e98719e4bc457149b74f8f0cda0c13a4af800e1747088c4533d2c53fbfc3d3b0f477753854b8a1da4ff35295fb79ae08088209bda2022fdf4a2f41be0e0d8b2bb815d8eccee1e025867a045db3de96f7b83907d1e6edd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e53c5f37d96446269b66585443a161c25c25967c40ad24b74ec0e95d485ef39e1040e1567bf16efc13ab40a35e20cf375055ab7bcc9411e9ecf829cb0564c2571be53d7727fa05952186f3291ee9ad8ee8cf48f738814208ea931;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea69a459a1158d8f2d071473b2189fba05125a96c5cfa355231147d8f9b813d0cd72c5fe0a2da136136756fb82882363b2d7ce83d8de941d787bf0c5beece152e929ff296518aa4c30b7904bc163e6aaeff687377456f47353f6d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f992c67c34ff5a47120503705576fa65eb8355116196a156cef7312ec681bc0710d5840fcb7354a75fee121e3b9e51a4dd2d6cb93259fb922a214f18302705655e521957b18f9f594cafe199de464c32a6992964b36c4781684c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a67d86e1507a459547e40df8e8cf0f02820f281aa4f52f79de2239c0afc7302b825b5d183ed4e3bcffe4343ae92d36eac9f3ff768e320a8f9a10156e36a3108065e1b6e388ed943286a4265062e6d6b443f5f5fea2c02c5567fe1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fcedcd49f04c1662f795745bd46137ec4b9b09319b4b02fd4085f8464986f342a38a3c3a65af9bf39ea2928734a241d9c3c1049db13d87ea9d70a56a095ae5957d61f841ad400126fa88e5a67bacd8c5eee2ee096e6fe08c7a55a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h714c71afc8b1955f9691b6a8c2c3d9c617aaf62cd850c74f1fccefa9a46cb8d65c0548fdf311a6b785b2438cfc68b8286a5293d03f84c0216ee67cd75cf1934556c7ada66996b216b007aef11601230ad3f859adc33d62fd39ad11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1722fedfa4e0d48aac96aeb130893eb6b56115de6999e143ef3bc50497e433c60e1b8cad76f97506bc482eac3c0dedec7edc9009eb2b719c7279dadb482f830c33d7da4f9aab2eb0934b829e5048e2dcb21dfa3b3c83f0389ae65fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1721951bae694f0ac92f4a7d5a6d04218fb0020689d21d3d6a33c23be517ba52063f0d18241f08c9940b336802bcfea48475521a5b227bb99331067d3c30de54261a808396682f504f640546c81f9cdc452b1879dd24cf3aedf5890;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haaa5fb7ed309b4ec0efa0a026ec3bd0b8e1ea941e663d3de788e344b3c135334ff53f4841f4fa9f80ee6510dd0f0fb80311dbbf9b06293a4ba9afe4e5904419e7f035726b5b81fd2ed00b2682b7c63c767d70a5bd3cd910e5253a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f80b14f5c08b6d4e805eae77330042b9a3b40140178832ad944a334543c517dff3711a4f7fbe73ec5d5ca19237ba5e8f12307bb7dea003322434fc8fb5040a3786a4db39d7795147d4aa0cd21340aa8cb02c13eeb1c888335818e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ebcb963baf2ddf210950976c1d2edbc76413f0694e8eddc9d39e61c0dc4af37a156367550536c59fcd398eb5f9372c6fbbc476d05431f8ef5451ef9643895f7adbeee66a73b51ba37530f00ad4cd4adbaac9fb97f4cbd750f27ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d4a4ac64551a641e1ef2b84fcf1a2f97fff311a72f8d48f0426c2d67726580355af31e2fded7d8a6826f432785c7ca6e966b07282bcb486a8e3cf5f0e672e6b15fe4abe08f9ff51d6917d8f3c4f642acbcbafedf7481afaac6174;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151e116da182cc683f80666beaef0928cc14b9c17e9a2e4ba96fa9c744c0d65a7e93fce2e64b01c7bd878a526413ab5703b92bdaf2525cd56e1962bdda0b69973f669d32d70f59135c63aa96808e83f82ee702b90bd47b78b4dd257;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ed7fa6e20d9b9a2aca9942f556e6f01a52e370c98cf638a3115332f2cb0b31bcb8097b395e5470e12bd44b12c092da713c0abcf0e4814dee984a796805f38f4a7cdb2732524c5fccd9ae88a65f39f742815b57a995696608fe946;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he85515c20ea3bf63ba0a6b3d5d049cef7a6624b4e75063a0ef3b1e0e408439c6c2bdec8c427be7c8338784a6f74d85de946ead919b87cefe5593e7c8b0ce7fa1af86a3292c1501df79e4ea31703a99e08929bea23e2d5aad7099aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165499c46aa42cca24233921438c1bed19f7d23119044fc03ec1058f1e304151ab8b78f0b55505b3c1a07dce42ddc28e520acf35bfc001bed09715c8f72896c5bc10981320f7d03f73916d9559bc67bb86280cab143adc9d0ec317;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e6326938ba913392fb67d26a362ef326ac3d47b677cd662f3751b74b45b1c9b9b9df1d5fc414302f9657edbd6d288ba0a628e6c4d791bc56f62c841a0eb844b7735e5de4c0d3d3dc8077903aa7d22241b13ea1a8e6fc000fdd227;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7eb671e61c9608d18cdbb95649d430e7de14fb20306dd95cc08d4f81eeadeaef5dc08da6b6a7808b4940692c86e333299505af14505b0e29697817030ebf96fafe2d13b2d66be957da8c2eff871206295c90ee21548c41f1853ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1460ea4044433508a7aa93ddb940777b39b91b0dda9af787c05bf1b9bc9575eadb5ee3a32610d3b58849aa94d2afbd2298aa3dfcd52135a1d24f4dd4959f10b592d0c3cbdcdca0ca27490bb2cd4042b095f33a3c034bc7ac313c97c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f792a8d49ffa9fe350a2771ae003d16b43bcb65dc106dfd1274a5d40ef8e4d5796f34d78549a99e40bc647039f3ad38f430e407a7b359661e892276c9929a233053090d4849a00d495665fd59b7cb361311d72c8b187f4953797a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dfe22f19e671f32d71c2c37fa14f241722f8c6fae393d299ac8dde43ffe44d39fbb101b090496e873c43d13b63edb952856c80a49c996d1ddeb0fd92edaed5e9c015270305f8fab0fb3d664c48e1a790def99a54ab1f8e4ce859f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e65fb53cf8809ad97b83714489e563123ae272d377cd0bd47aa764a2b9c1fdd027e23a748ede5e659cbd0d610744abf3b5ee9231357a3a72f3ab714dccdc5612d1b140e07aba0c1415e1d721ad0541267b5bdbbed5e487910ceab8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172b44cbc4ca208298295e106c7c477aa7591508453536be00ba2349e64479bea2479c215459b86da3a81ec9621e96ef6218d36bd7d85fb53bf9fdbacf0e2f82ec54a1f4630e0978fe7b431a5e1d5931d0793ea51426ac36e97f3b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ab2a334f5a3db55f67f8b0e6e95906eb87eecd9c62139b0a0900d79247ef2f33aa0686ab8884b27704d6496c9c203b09c9ece85b3d412367d15c7768d906eb413e71597fc054adad25d508c0b2925a7b0b9bbcc6b918ca255c7ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11460a21f83f182ee078874db9a43f43ce7b9c778e9e719e865f8e77ebc7df736238dec20c1400bd3f40b5cd8f57295c6b443b29fe2274a5d8ed75a67e31e8983d5890f91279e80aa8dc0fb69d091d2690f782de7a7611bd762e49c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa03f73a1bfe92f617175cfd255ab601c78187b0744201b04f05f99416ac5546da214ebb5cc1b94a684d5f8790014c65072b6327d8e71da05f91cb1a84211012c8f64438fa15ccc5aa972f2a9350c77b4a407f1bb49c54d864c774;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d81a95c7a4d4e05b5a66074b6ea9aa9151e8b47fd6db3d9e22c410ed0cd046998f211b7ded94a048b68c14088c0769cf90c022f51c09cac5761a33e94cdce4bcc92140e3c21e99a4914086f838a4c8cead1e19b7052fbbdecae065;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eea64c5711936e4c2f9ad977f8fc5a12e82c4c90764b636fb755ad124fff90f9a26581db176756efb35e921be089b57d9302f0a41b161069e246a706185e52306edbddaf87e695db418ceb74ed447fa4d3800499500b1e9447a7b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baedfa5424dde7b3d8aa12f6baa8548a588c499e0d25f0ba188c7678f449234ebee4365f5f5bdd00cb5b3dcb003b75ff3fd25d8eb46346ae281eaf820d00c52a0b06a625ca078e0c08fc211e2a1512c13081b2f5f154131ee6bbd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23583ebbb4cda36283945e5692fb9443db72e809377fc60515267d1ed5e91717fdc585735f08d97e8c3714f4b153ef13f7c848a8d52dd5b5e04ec1ce51d39cc041d6f5a41a46da32d4d16f8537900088ef1acd6298fc87fc4a5be8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b1223f9a749da97994dabbbe2d01127b5587c0f990edaa62874046de1c43c17d1f1dee1a56f1c4de109c49ea8b2df8ea64b3be548c1927f7d98f0639148b8035022d557fad76d24e079c764493852fad847808877bde021e72038;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1305f245d431751229f74511248144d3fa30e2382fc7820754506bf812d942c9a414ace0d25d27459b27c1e6d9fe7c46a36879551ec5528d9e3bf9b8f74593385e78f35745e35debd100572fc148a04da41c996d73d765309a90cd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116fb0aaafe80a8a0e93a34d7114d1c9fb44b12115bede36f89b843b0ee8c33b3c119a423cd117fb497cf7c127d8591f4ccbeba91d2791fda1772f77bddb403e359492e35381131039ba901ff502866c457a7f6578ff543be76b040;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18108c51197c27cad0ccab3dffa404634990221a3d6d83d5f1fca7399b345cdc7289d36dd0151d4611f6358807b74abd488e20ccabb699de4381373fbcded4fd1f12b1b0120f7701232974b2f4db554842702be7048182b66491372;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e0aef32638b7d88ef0d19e22a383755848227bdd5c970bf0c4c7f6937c155f2883d597e0b55354a7adacfa7bfcd5ed07cd69f58cea34a5c59c6886f0cf9c795c7c008740c978768fb0b74e26d8030b2c4800f57eff46af0ece90c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae76c0b24972ca3cd6744df6fea754d2bfd2246007a55edd83770ef7b09e6b4b9c8eaf6abb5fadd91a441688cf12fbe85e590f6afd7dc6eeebb1bcb702a919bf7505ed0daddf95641bd4d6a91eac8a65a47d8a39ef7dc0d40dad2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ef3439fb2aa923c27d24a4564c901d203ebcaebd2b8c39b046d9de1fa1282d531ddc3c9f105aaf4bde947b509f979452b072d46af84835e9c2b392dfbaf5c83a11f7381d66654b14ec6e6c41f3aa15d8829e6190a71bb4bb0ee3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c1f19bcf1821a45ee300750a23f8eca525f0894f71fe7bbd771587a228b6905f85bf848cecc0f1d463f3ef85ef6cbc8fd50bef9ee0bda9bfccc66325ef08ee6dcd12e5bf9bc486b213902af073411333d861905a3a07022ee4f07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bdadfc0c6ca88ee6dadf78a7f3e4a4fd0bb503baf874b381383afbacd0c313c48d6d558136e535cb810de073d19aca1112c1e21d119261a3a8b48c82ae1e5ff4def4afc75aba69ba37d29450a12d9086db297c0014c02759afdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5eeabff6fd4c6d323b19dbd1a0b05b88122a524e83fa1dc4c2a9f714dd9ec29d36e65d2d3b8dc2c16c9db325e5b2da554f5ca034f7c3c27dc3ee39913b405c65d85f85d140cf40e32fa99f0b4ba289893b2fa486f25c578f823277;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87e4c75a5cb50b3dda15771d7b73624f7b0f32d325730d84a8eb3b11b525541dea8af7ee77cdf4f611c365cefd230ada46bf43591e27163dcbd7b44faf836ed987ef82db1093f1d8b9ca0bf44866a59531252ecb325063fdfb9b60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114c15070ae0d04515587fa836270269d7fc92071486fedf67c7b8d92e66fff723edc853d6b493fda9ab8b0e2d29ca9914c2a3f25c032b3d62c05938d6d0c0f9ba759b57a348a14c58b4a5f4bd2f309b0722997611e82a4ae48bf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3eb3be2ed4de362674b1cd6ca5419d1f3fa5477f5e7506d4c2c6660add7cbfa4fcdda985f0bec8a68d4c3ebdbbb03aef928673d43ebde4338873ebc2d8fcc1fc5066b2080bb54fbe903852576a2be1f05eed0534744ea73ca972d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a331effb8709fb5a74410668e4b5a105701d7a3667da5591899649319b3372a1d27d9b762974674176c4e27d9bfa834ab8d2864487d8d374ea34e05bf417c14e5df8d4d7f36aee69d5f4582530e9b7c632bfbe7a677ad54c5e16d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12edd5538992fbf08aec984ed745bd65633eef107db77452745bb0ff6f17a7343a920f5dfe4f2076e47589c15281c1a46cb37469be09f49d40c849925a4cb1f264e822b373e583850a0d3f4b68372c5082a9582eec8fba372c847;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f0798929337decd6810d7206514bbdc54719588e914aebb57382e9ec0bb90ca717004349e9a0aac10ce4535a50e7c705907ba586ccc6eb122f3c2a923022f42d75e8c8aec4a96fb6847eb9d5e3d9d594146700b57948bedc6b759;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bf1779015b72df534e40eb41115516c9a3f84443768b28e98122e83782378d338a6c799175756db0f154a493e9e616aeb52c7ae5c7113e17df8901c0bfefc138238cb3754233494762aa4da3bbd7485939cf5f137efd44fbd0a72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d718877e1e1027ecfd90f2c7cc384379330fbacfd540cf81bc0d70698046ca0ac776736e4612999746ade79b62bc9f754689235b9227e13ca99bf9ff774e229eb3680cfbfe03c1e34e9b25c3e04ab0330000ac41c01dfb21858b2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha901d2b49c694f01d9e140ae9a22841ff44df6be4ed54c6ba5245da080144844ae5ac76e35fcaba57e43b4d1b99e9a0ee30c83661f818c73bb5fd4d7d8153def7dfab1d0ad65dc98d8c6a94ff8f32e1d797e50801d5574efe7690d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c12c8f287aac8f0b1a4f8204e243b6bfeeee861d627327c34a6663bb639bf762d960813a8ad71c44f136f15159a5c2fae6ada5f501a04a335ea70c2f64c96191ddf3062ffd573b87df5f2f23b860f0246e60847958a2d20a2d3a8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6398d97a2c395faa99826fc6a1fa21236a6b46f19d2fe80492ae193026970855290a47fea4dc5225270ed6d78639e48cb3d87cf4f7031473ee0d8fde573368768edcb619c3cbad9f2377f1f7b216bfc0ba16d2f3e1aa1429d7958f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1396562a025c66ab3c9445f73fea5102b8e23f12b3b22822c3c9d964c87d6dca47e91713500abd673d43085731be3341e028f6f7f625b2ae9320e253e0c40b5ea24e658202cc0fd6e5b576c5bc759e76e90c6d191b8cad30b7a2897;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec71c1354ec950df1dcd294fe80e5bfdd2945c08841a017199e0ea1ce916101feb571ad23d35d01aac9a11272481c425f81d371dc6f7a8f9bbf3fe0f0c70c0d0a9a5038949881927f4d5dbd1bd205df58f63b415d3ce42619b1778;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7803e38b5dea79319cabeb50551052bd9920966e606b9aa56c2431f40cd575cf6768f4ebb188305600312e476a9fcf3d7036901f9a396705f8c919222a25e4e09eafadea788c62cb970b6dd8136629734feb1b902479bf92deb460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61ed49d55a248e606ecf0f8c9c45d2a407e31e835036731908dfd8787586230884763a5f1c720c42673685378e56a318135cbb708e791364f5730d016a850cb43325853d1c72c1857c1c6daacf02c1b9d24e65cf898c9aa25b4cab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d8e11961255ed3e2c97e211f9a17ed559b75b02c74236576df12b5a5eef155193d2cd191efb440b0fdff8e854da5b5a9e7a3da39997fc2e82ea1c34c17525345f9b02649ade40370c51ab16e8a4a418acdc8557adcc4a8e45706a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3cc8dc641f8d4b88d3b979990a806edc45f158c24260a599c7b162916c45bdf4dd294ed867790f5517c4ff55f63cf5468e5d98672128be1d76015c085547be99442efc84a4989b923a7d7314ba967ad3147555b28039c62bdecf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17934f99e27a7750bbe4579bb3f22b7a93660cd85d6e4be8620532ad7827233ca1e4194d70f54cc8a86d9e17d0f1135a3d6a9ec73d8be45d737de14cb4cd8023d99a293602bf70fed38d48b938a9555676a7725dbcfd0eff8610f7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bf0a6c487cc80c3e24498acee0f76cbc9cc939f21293601a0fde4dc33593203263564bd68206a25f2e27208e04539cca23027d76b3ccee31d71b6b5ddae0ba1a91bd99deed04ce848624421f12d1e331bf8023283ab647cf8cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdeff990b33f61006fc7ef0c86f68c871a575e7bed8bd0b1ddba6dab20a8eaa1fabce4e6e727dce598c4b7ee279b175824d0522746e00dea23f96577c7004653653b6d1aa705e71ced40f7748a62e8c6327ae451d62f094c6712c36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70cdf1300a4e42525d4d736d29c458e2dc835685368014c2d6be13bf3064b8b52c14d2c9b196ac6bd47173f6a0ca0e6fa1779d65d90daeaf916a2179487481c9e02082a21acdc50f36e4dc201cd98896d2026df1708071b031fdb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h52f8717691df4dc39dd763db1812f986d09eef21d109a8dd5a3af6f7c6a77e103818d46620e7b2f4b17980e9c5ec70d8ad754cd7b99945f26465a830a6172bb4f50776e64b2c1e54bbe1816778b1198fbae9309ccc6a111e6d4d22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cdd995d2b9d34bb98adb2549c357626d2fecbffed59081ab7dee18f1ed0ddf4a4d34395bc142fe51513ec557b6c0d0d9887419e7b2d8f62fe7dd336a3b0acfb45a23dba81f174a999401fc8717fc4cba1a9ff1610aa73e6fd3ac08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h249810838d49c69e29266bf45b8c79670282344d2512a6affa7abda57e28d73086159c4116dc85d80c3efcf6646339ddfca4780dc226bd9bde221b0c5ac498dee281719deb7568b8a5ebeb69f92131417395610fd271e0c841cf74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b726d25151263450b5157207071d33edcd7282a404babe06982543b6932c4511ce93acc62e7df890543c4d251075da9be1e762a5fbc7e42b76bd5768baa6a2188c7291ef6b9072fcc3f4f40a678d478a82d795b845892a7d70959;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea4c747692a21f9a898ca099ca38d7791f2effa7dd7d2459ac76c67b5aa0d2dc1721361be3b692c08f736b764d5a055a49e98577071431480753f8a9e72335fd67cdd70570bcab1b6e6cd63bdd8eb795c079b53056fc421a363421;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4a959b41f8fef9bd61b06e13fb7f53dd7b0ad95c5767aa0c78088c8f9e34f298d56fb0903d08f102acd70ede45f63fb1bf7c995bdaef24a0df39393ef590dc906c5f29498cdf8000e7aa1a1f5d54a2f0e1f5d8f272f9247b248c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83896835cefb72d78a3d25024e95ef2692155a070dc66c898e5f86960a018235abae1af26b31d3c1360f2b79f33e2023a1d791ef2e12fab1cbd4fa0227078d9e91ef0d38469fa34b7360a78fe3f7ca1ea52d68891d907b0d3f068c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f624d2d57cf9d6717d958630eb7cfea53ec111d65e80e1559ece8ac3467060cf78e30d2d88a8346ecf3c6d093116612e2882e8789c8a917bf7fdd2e62fe23b355af6eff472e5dda7d5b7f3630696f8d42d4816d20d49eaad45ad6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c667b1e62235f02a46a0abbe487dc2e23624d105236bee0d254220788fae2985e1d081917d28273f3afb747d3056172c3723f7a2481bad189bba82006863e3c41c4e0e9fcc7150272be1af21ed9805a2932c38bf56ff066af6e39b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d24c1a1c5dca14f44a81ebd8e8139c5f0570c5eeb5d60416b17e0520eaf551cabacc8ee10dccfefaece5624b2dd64ff9199cee59291367eb8254730a553e47ead67ddff05cbcab6a57ae016c3d144a67ed53b7876198aabe6626c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db9d0985c2e8e935ba4efcdc27b708fd9516ba0b3db679669b8dd71b3427068514da352b58c3dfaf30dcb1222bcda7785963f849f708dd95e74a782599d855d8811ab0cf49fa10422857e823705c20e6226ff36e1acf2fb72946cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18343bd525da50179b86bbdfa581beff3d07afe9a35502a47da055d76708089636db96f913f194a74d6faa4ab0427011f0bdd7fe69a2db26ba70192d79257e7b0a4fed2b6b8a0cf41f4e385ed6911757df445a3fbb01df39efa55ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15528c535a2ab8863f860916019e73ccd27ed8b7cd9d8a23fa818251ec36d0f0464f7b6a299c847272213c147109be1d584fbc6833e45a9b321a7d54aea3dcf0106ac81d6ab54f62efb09906d6ac6b980c83de420413ecb653c6523;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1886a8f02da608152d6169f942d407f97bc514eb8e1c4b0d3596806fbb8dfe368dfc2ef8039618bfe29923a235ca8cb1547da2a993bd3a83d16105d87ab71e8ffc10cc090289e4898a14287b7a737bc4c394a7fbdfa6f9e6b0e13e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h252776f12c081f8bdb5b12017bbd11b50080978aaff26672d8ecc3b4ec2af03803bb82e565765cffe7912c9185630c61e092886988e62bbda6fe27d42a4cb44ce9ade3f213c74d7aa1eaba2bc35344bd4f9b2f73e8880781c865a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bba0631e8055fe435099596925f31ce5189a8cb31ff21bb2580d3e6b85a3fdfb8e93bcb918db74969211d6a30460bdbcc4998295100908212aa88ad369db9140cb687381c2524e94da6c5471bae18c1e50e6a59f17cdba1c992b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha22647eef9dac66b02375b29da2a469490e49e27552f2d8684498b017d16a0216546bea437d383135f50e1965882e9c61cef447b0c96734d5be4d6a7bf060e14bd8c98cb39be12f0d74df89a55ab7afdc988af4c0967e4538b88b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69ff8775a1bff566c7d4bb0b0cf007702d4a035c09396e8fdc42f66f59b9fb971ab1a5c907739f0bd333435728d49bff92d3a8e99213feaf559e8c1a1012be38f19c5595eddd828ac903298ffb1c6b9ebeb428c87b0463f86346f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185e20c421faabe6c081687d823fede292bd293f9db73e70696f3e5ba32d32e35edb7c3dd885c1e11c05af6683140531f569fd1f9d7a948dd159bbdb87a0e4e9f7f8f2312106a3722a31d73f71c50a6bc9d509d1b550ac36ac38c71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbae79de1af0209fc4b8e7952ac06a83d6aa247fd772e36f47dea0ba90d0831c7d1890f52f3a582cadd1b74d80f37fdc97e11b1cf6959c79e0fb2c78f9a9b75d97616c510f1d3d4999f9aa42e76398d918fa989c6acd18db5ac6f35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67087a616a80e3852e54d7f9a2756c041be5b4a5a487cb7928d8f9a8c2c777d26c477666afe83c8cfea1d30b9e0d94b96b18d835dbf7dd86b1ca9d28b3e8687b651f775f0c345e09b57bbe4c2dd222132200660739ea9b0468493f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f25495b244eaed7da608520d4b33c3b89afc49b425c2c38be74dd2458cc80f85f87cf46433d8d04c7ee6058c032c772a55988a90a8211aa1316bbfe1097405efcb405fe409b967839364411d686faac2c470498863464bc123e60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1007bb6824b78133a4480b531c6a3957450de073c8a724eebb766fc84a4c74d662c3055437de20badc77a49522abc6bc89d340b59b1db8bc77602fdf3aa81d75a435e8abc9ccb97928cd3a32328da6a38947ac8c843ec53edd64cdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9e31c7c44d795a687020f20d0620c431270812fd50201b2509949ac366e20ac741732d4ce8e757b0b876ab79ffe2f69540ba522a89edac816559b13b6c2adf3420b13976886af5a1e0036f6ad47d7cbe3176f8607d68fdb35f6e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0fe7fac389120fbdfabd7e05d7fac27264d91bc9a548f4606c5122790c98c6066e34b35876055655adf3e62e744c05a35c3b46f0c45afc6a97e221c82563a354bf548e0123286c72bd10d2d8314263aca41e8b7482e9241aedf59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha07861af9f862e5ad04208c9d036fcbb02333b74c51579ed80fb8cdc7ee78705febe3967eb4a5403dd4aa2c6ca56082357c326af352baab6504e59299174a538953d4b9faf0058c33f9f85542ddf667ed259e717d532931697596f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7aef4b6122743f97517aa4e942e89cf83feb77d80f8d4ac9e44ce952bb7b3f775f607a3ec3a9170209790550fb589918a6428704142de25bfe6f9567b1f6560bd8f0fb32d62078f85488e111ffa91d73778c1c65f04976b8551327;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf855d97bb0c03f16266bf9cab0792eeeffa31c6a11e2c1d83fffb67bc7ae2bc41904a45126e8713dc76375ead83ddd86e715e63eafc46c410e106cfc2573b9b952209504812e143532a71dee7e22de9e9ff272563e68d49e43df42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142958eb961980c2819ac1bb6a57623eccb01d8e63a1ff2e0447c482c626e0d4a2b9976e3b82dd3c6b58552a9ab0ce904357e61ce440a7c5bddfdf9fa401eea23c7ec03286ad8e455ac78383726e8c3b20819871e41b60c351ca2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b933ae03b96280dd2144342627d139100a481529eb574ce148ab7f12dc80fbb0560f39270197fec9d3899289535a3f500b30e15f7898c6795eb1742a51e91d007975ae830a5cad6ed9694a37dd8ac75bc92ebdaa67dd52d367a0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166da57c3f9a528afee4a3ac455fd6b912734dd020237f99fb8d9628f31948e953ddf37453767397156a85dd456d06903dc2947808158d0724ba42c5bc97b8be2a7ed5b56cc7271ce4c2dcb8deb77e67f23a00b8ee021b8c97241a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1ec641d35190c9feb5ed092cb1603f00676a36ea642827fc0c7d783f3d544be7884f49706477855b7fa71ae23abb76f63552f5c0ffc7a36e0afa1d0e602986124c09904bee96c6e0b1bd47dfd9a2edbf9cc5cac6694df9ba72a5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e45c2f9549cd55b5d8f9975343f1424ac3bb9d97eae5a9bd0b37954c7f60dbc48b8290e804ef3da681a5e76db6fda88e9f3e2d29016ed101651abcfb9ec6002c9a7738e8b6408483df25c67760413fbc8cdc5b3d129d8f006bf173;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb225fb10c1bc80fb341405bca7a93a3c3b12ca92440aed367f4d9df843d8cdcd30c0b35f8acbd95b3d5ef95c511882fe507c283ab20db84e2b67f591460249dfca6d736dafba2d22d3ba440b0eb4d4233e431c17d5fd448d27c08e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166cf621347a9feaa59e5696c337ed2b2a608261385b4fe6bc402023bf141fd957fd5e15c992d525362904f5ef49138f5d5e6117c5b0456536fb83b0ed243e02095f68cfd704619608c63261d4e71613d7ff0d742510660584d3274;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f6a290a17cc3ce21c995d4dbfd828aaaee14ab481a1107dcb55e28120acbca4f3d87ffd24b41eaf240ddeb428c24023ff2c8b16c7287cab12a1945616a6f1ea641162a3f32e5dfd9b3cc6d3b05ac591debc922ed06b5616d527ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132a8fd678c712b2f2e4f3aedd85619a28799728086e6145ca1f762df93f57bd015d19c3999d856da33f6f90f9ef67cc8f7c399f4ecf394b00e5fa725262b407aafe84a80f47a0df6aae88b33ea0cc7f9622914b21bf0e58c16076a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6f0bacc085f08cd8446715a779714d61751bd09639af5a55fc2e68adf4bcd649c9c57258a4ee82102c2bd26dfd6bf7c827ff3cfe4c5d7d5b5139f3ea4cd3a55e32385f258fa054e33fc822cae604f281fee4bb19e5bc9188277ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9b6105a609654256b993ec3cd830fbcf1ced8ae5e1a00572931503bd02b35f69a9e4993a586bc5c17f28a9341cf0c3dabc2a7ad8ab4b0473f718512429306cce6f93050975b491741b668f2a285020437b65cfe4a5b4356a4fe16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77242d2d7145ce1cee95e0a53cf158128a7213c1483c5bf8b34fa9930436df40a4161fcff9dc6fc86e0a5823ce21f611a7bc6744abc241549c42f7a2986c3c4185750f723ee6c15dea3c0b14fda2728fcb50ad2d5295bd3e13074d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h896c54939bcbce868b65c38971d76fcbc564f42cccd528455dad8aeeef92eafb586b222dd8106a007fa2053cff8eafe53c0f1f62d89013aa248bd1b67baa2abaee53781231a20cf046ffbc5ae1bdae86638be7f1f6e787f5c2cd03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54fadbfcfbd2aba139c7f6e81fa91129211b95619bd9acf3b79b96b3d0c4956fe6488549d8e188c3d4e7f9f0ea330e750137a2007422c5e9df51c192ff83c69c3b5b74134ca4005f49cdea27e941324844eb165c565fdc12b94c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7021cf7a81feb2d14e8c6f21b8ef96989183533b13982c01d52f5e42a87eb943b2142a8d45ee49c320806c625494fdf5a0ca06016bf537acddd72eaedb351eed7b415e7829b078a4c76ec0e7b8cc4c48b818d48bcc87a31381cc07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98e6d8f2871195cdfdccf400b3de62e3942c113c9fff21ec7357bbadff3da49406b42ae1df19539c090fde7bd6051a0bf2e3277bff36a6605468ec5b069a785fc01cc486cc9962326606b42a211482b8e8b2edab0c3b697e56e110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c641d1662748a4ef9d7f25ef08b00ea0fed13b2719f8994cd70bddcca50e99f69d5a0e56b596d0d8ad22710dca0698888f892fd89a53c3a5f25c98c3e4febd78a35bc83a9fbc2e0f21f47fddf97253962fb9ad944f32b5b9d1db84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1effc2fb091c4c86a9b424f26ee9604299b4ffa4cc468773086c10d94ab82ffd4fa3dbf3d10d59db3ac8ac4f0e745ee9dbc958ac6d48a6fe321a33036e8fe14be8d0826d3ed90481e87b6f5a2b54f53b1dc0b3a1134d052a9b57fb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha65fd2749af827ed60fe6e07caaeaf7bdb1cb54466353ec5d7dd7151a53c687de2d0a3a7405b31417bbc63cf57cb1e94d1cb471771aef5e79ae57d37e563b6dbcfe97599577206150efbac23bc5c02981156d0e12958762ddf0890;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa1edb737739fb1e7f0d8dbe1c9a0e10f75cc1d8defadb8176da2c1cbf5106f9c1b2a41fbb5c4be7f263f96bdacf57699869f470b1f6b54581278f1ac466492802c721d4b1ee5798f00ee58a34d9a1e1862093b5c26259fd3ffbb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7abe6b7a57d8ace80f7c508eb863289da366fc2df05d37f97a604df52a913df6f25e21583399af5a7c9f9d7132a6454107a805abc6dec86a053d36efa3084f14df3c105c1680311e4e835a93b6d77707e81880bd193ec824106938;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1691ebb8bd6ad39aecbc4aa14e50a17fa8895662b71da0d9ed6f51bf9f2e15c93178542c5151f3a2e71814f02e53cf67f6498b8cdd245b49c656248dacc2ed67a93dd7385dece9ec0d954addb6249ae06bcd67b26e45d2ba3a60f04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11685c5f94a112e2bf79caf83d624d392b59297d2a558ab867b1f2d0ec6394d2051d5bdb36b04b6661bbfc6b034ead8b7a61a506c1bfed98acdc30a963bce6463de7be7c802e9553068f80fffa1a343552c57e51568ee3ea51f9225;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c3465b039c7d9554e585ebffa3693a1acddcedfcd1c3c72df0c8e9b21f123cde0fc2808651585b08987e711b0b463bacb555755515d2f03976b418a9a91f03c49ee71c490c45252189f21f8cb7f7b19b8884b04bbecb056b1500e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7127f39e8563fa1e97f5e72a656e62597d5c117b803739b0b9dd04e15f8f1d6ac00efd0956edfe51867a19ae3ee502046d915494d9bd27d4121c67febd586574d43fb39ce9a7abae4822e3621979d298590777b064b1aaa1da0cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11aa5c6077a555a3d7a5e5522b4c34df1d77d37765252ef30bcf477bc45d8f7fd2cf9ea4fc141dd82e7b9665525a04242a78666546aa186853bffe3f7959a8d61bad1b0d15a1c342376d9108c76b1a418bf2af683a42e38acf78e27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183ab66e05ba21e7ec903a640569aa91f85dcc3d9c2e46fabb0244e5939538d8f5ccfa537eb000de30f244ea2ff7799d24d28d018bf9eb88da92ebf48781bb71fc475ca65c2d9b4d79c4789b3762e723770c92780ed7d7a7ac8a7e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178578a87e05303884dc17302acf884d88f046c1713416f18ad28f351b23d151d6072cba94c692e3dcd5ba83ff434309e65f037f7aaef3cabbfbda6b87b76c0a86b0f667c854d5d268adf10ea09dcefcbe5070f48270843843dc839;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b2d007860c86b19a748a5d94623fbe08a90e47118232c4b867136084d6086d28cb448781571deac1fae5378d5da5e7a96617e30e6676077f9525945cca680a018755cd8ab5e5d6a358b06ffc2bc703d877b7c3d0fbfa4a987da27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2affd4f9323f033d38109748160d289361d41b7b6b5e04329ca8fe783ee53535e2971d77400302c6df28416bd8a821150ec9b75ade0d2562c75c6217f1e2808069fd0fd8d06dcbb043ca53e0eb0b8af0b0546f8d0182c1f22f9418;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4261452646b5fde0a6185e18d62cfa92de0ff7315ea905a0e86be31f43067ea347028eaebbfb3cb8d487125bc3cb9761c8e5f608cf36bc0f99c9cff8f51b3792f3a0be52de0d27a078d1bf2d60611eb3e4c2044509b02da21bd02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f47f0d43a2b92bbdb1f923c1fb47ea49d746ce17370a81d49152e470e51dbd42aa6c5d7d6312b3e94e154c7d934a9e79771a73a80e083b664ac3e009aa4c1d62bd0d05deb4a2a71431fabc3f111a8685eac1586f422c0001a795f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13bf7beed9db95199c7b6240e0fade10c78aab5b03f06b0dc693ad262ebc612dde13ec57ad30d8a29ec85ee33f9dca5476d9d751ad71f7bf933eb102a0f47b5687c028a968d58dd7fe9e035cd42c8934a27c9a2f943a89027a6bd50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c7c5c01dff9d0abc04a8f806b92e26bf4c5265df7f399c6fb40b1f717ad9452a976e6c8f8bfa45336ae74dbd96dd0db4428d0e4b44777c5483dfd327fa16e1e14e566cc1e420664b7ee2e53b674a901db148af7af934c6cbceabf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5539c7769cd7bc15156010a1b7fa352a0dbd82ba837a02e2c85cdb68dc1899534b3645c2bd52440bd64d84aae85e9cf4b7b4bde0595baf9217809eb636af9b68f47b31599b2c5851874dbcf267846017599122d33d9494b71246;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143b74579615a59d0769b753984d0986298593e607b2057f854b03bf0bc6613a715b8b21e22d97f78bcdee501a3916d9276eca70b3dfb02bc4429ed227bebde19517e026ca13dc0413d3c90c677e241bfaa3ea31014e28b4f6c82c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db71e1ddc3dfae4c012efdb49d70620a18be3e66eca4b449b55c1a62fb6dd1f9d5b4bf8f76b095a60f6f829ce7b0a7bb74f3921455056a5b5b643ce3f7a3e1d770acc14e2a066f134308cfb3154bdff59479fd5ca58fa25c7d92a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134e414018fc7723deb155c9212463decb17e10f94d2506e20001bdfc466e5a52708689c3ff1a40bd7106b82eebd10a91a81dd81254fff881571a80d59c72f9d947a055b5ce9f6054595320fb111458f2bd04830aeaca33b73f2427;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1808dd64e29a0d39d65cbec2e242c9b9878bf36606043f6eea02687f4752ea26075f8608dc35567137bcfa97fd73166174d984eee3f73b34392cc79c1e9a13f44f93dd1aae40928d6d487f2be4745701418af330d1512afc40cc7d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bfae86589123a93c06d4adcc42d86317ceebf60bee808f014203a75ede2c777d96f9f270adf7e06619655113294c14d97c8c471a08df004aeb4430dcdc358bfc4e88eb0bb5c112b72e6787d29566218ba39253e6e5f09fe4ef7a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174262752469586ec10fa3da85a7ba0c73bb5ec30764422ca93ed28d9248fe40099f1e9c34373ed0904f658ee1515ff9c5871a129ffdbaa51975db80de27bf83b68ca8afcf2f2abe9b998e8dd148ad86090796d881f218ec02bd426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd04d0f17ce9d2fdc0aa12d10335528025cf126b86ea7348d279c0a6eb1cdf83e470754bbd71628c0b1ac83ec111e115761d930be71e379daa97cb278031b22d4acf05a893be78e0bfe444487694615f9cf810aeb9a375f304948b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130c15a974fbb66089f80e89577f2506556f0415557ad9f9286844cf9947a84a023e715d38b2d1e81a6e725b8e1feaa0bd75d9d5481b6982c128ffeeac16d78e48d9cd40ac89e2598b1f956309f166b2f798c6d69c05aa680abc4ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d71a05b16d352aae55d3ac5d5a9240f1f67eb17f19f03677055fa8e281496f0061787bc408cc913511365716f03d4df2125f9631883da1e4de97ea6af8545c006385712d1026ca452a9a0111fd9a819c5bcfc52d053b4fa27a0390;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ce7c36b107763ffa8ac8da47b7cfe98f27e6c24b0e1349217d515fd864c47b8f4e257c02c0b941c0b44a61902096be18c74c9b2bd520e624f5f58b940f56ededba86beddd5388c0baffd0a2e3e7321f3703dbb8778a886cbf6a29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1569ad37c78aec4cacac0f70d9d4f24798141d3ee4786551efc86e5d727597ab34a663f1bbae596954ce95a6eb593b600635f08a8646a96e0312afa1d385296255c05ff5fa91e986f069c36c90cda8973fac5f09247729aec627f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baff5a57b51eb5a6f95b78194f1942fa30bcf07e0f7694b95a187d70bb27d986b092c04936ed278fce3e0b8acc490ee2f57f6ad884bc5ad5bcf5152e3757730cffe0952e849cc9efbf52ab7eb63ea7c5da8410fb1b07fd6caab364;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc54502c56a1d37e3100bbb6a0e24ca03bc8c6c19ef13054ec851dc07fcc16fbfe62fad1bfb49a8e9c1922c9f9d3ac9294cd4e2fe15104c124af28c081beb53d33645cdadd6344e1b938b3f64079801658aee9198c1e9db2e4fc4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5e2246fd0a09e9b4559d9d30ebcb891306cc6b5d1f0fd11818d5d90a3e26d94b23f6d3e82d234bf99cd3fffe15740e2491d1a195c71a88636f6e3ea9247b75d78c94f08323b27af56637e300a07ca8c33975eea02a5faa9010b3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b6bb360f341d2bd79b0d9ee0b7664a3c6dd335228f651b3dfaa1f95a4d8b7d54dcd3346d4b06cb5f2f6bab54b20e60d5fbb564bf0675886cb6925acb855b15a57d3aa0d2348b5788ab521ca28447529ef268ff28766eeb3e9f836;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haaa573e926559c568e2491bbc9bd2e722d95f78d2e69a2f849be0c6ecb4da6171ead358f78f05b7fcc8262367abb5b40763d55edda12e382eb106e08c903de3267a474eb1935ef60bfe79694f7daf1a13ca888def57988ebc5f8de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a50bf21d936f3061e111af3c28257b26f9d5c1be7afeeac9b2953ca67310e0bd8cb52a0abc77db2766647b0de674250e5941b9ed73b6027b365b816750886ec35b2a787cec21d0554aeff160429851970b9bf9ca650aea55d920d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f63e006f61b15af3dc42e285fae8b197c687fcd26f0ec7ab39d411169d94fcc3b9632d14d64459f16847fede823de3b1e22a8a905204b2f44482cbbedccdf3417917137824430c4c589aa9dd7c8eb1a1c9ea18855f9c000b207dd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f54165d256838cf2f75e1c7b4b0cc4b65d228431429ced58e939701400b262ca3c970857a7b79c12977ddca7f81292f76590570bb1d8ecdbdf3ce634fe9be49fdbbf9c254a43ab040e65cc9af5b00b97fba78722dabeb54a5ed9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fcb912a17c670996758033011dfdf6938a38b3914dd283bd8b123aae34f0fabcff225019a0f31d7fa5ce4ec2c74ea3287ec3ffc3267cf2b89e33a0ab45bb325063d0fa537a1fc79209e574c71bb0732e74d2b3bc06f504ccff0f8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h346042dd24b008efec2e8b1224f1ade5a24cf166ad4ff3b7654fb1604dbdc00d69251d7f11846a9e622f056767ef924ceb7665b63fb9889a6104ec167d2e6f81256d18989810a1d36aee700481f4f6fd1674ed34a247264a2e045e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ff9fa30b4f16cfd49b5827d4f70bf72e43a5aa17c235d197f174de75f41553144741eb47d61c886b2800cfaddfed03a3276bd718c5a163371352286554756e56b76bb69b863d583ae7b57d8ea8b3c1d570b7d8ab6ebb566c718b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199695d351ae828cf24676b90394ba7b0ba0504072c7330b036c926089b444c10ab586bbc68d7dc11b170f49641c7d829437f538649e3b4c34cb7b812f4f23e51f1cf7651530997f91811d705cecf156e5b2c3f7abb2e185924f857;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e99206230686c0625b7ec815ae3e9809b2cb51e97b3c0ec2278dd117120943061e5cd8aeac7e9147aed0e4e6735c6dec5f2efc967fd483a61ef2c236cb04593e2fbd93209ff673437bd3c8992b49595d955ede96412621942c43fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c86ad01f50c68c6c23838ccbc5f064a2223de0ed54b993013aff30aa4056ca1e6bf06a726d572d47ac129158371cc4fc806f7b6d57595f98b8fce9af820c403991df4b22f29c69a1628965213548eb99229958a5d84b1f86b3572;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10524d70bf673dd3c8e7fa24e8441da8b8c06d1b18d4e0fe63ec1753aac84025381b4d6f3e5eed72bdc50269021c8b1d3aee7c00154bbafb3064076d825169e27fd8d7cb1c283986b85b3d4a9b9cc6010b9c141a6c72f4332ffedf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d2d3f845bbbf76f20d990c2145016d87576390c69bf748821e92d7517ae12a7a3dcc0197f1611dfc017cff3eb5a615e6daa568d01b7edacd4b423c1444f0bb30a7f85a8c3a5616b5cb4c83465a1e64e3eb018251a79af0fbe696e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a031b52ef298be41103cba59ab6e9366fdb2038094fd2f648528d1f4cdc8513ead1b48e67be2c3c036a08319f29dbcccab749094de5342cf670205221723ffd9acdabd0d7e35b78673ee000a22b7fdf72baf1336b12c66890728c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8777b77e0ea757d1612a1dd9d1697c208612faf1515107924dc56b3ee81bbd4889dd39d6970c94439de51cf556253d26046b4bca7ee4d3fde37e4842d2262f3b8e6ad165b53169f50fc99eaf9ea80062a0b307bf009609a368432c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6813c6568589f9ffe8783a3bb0fe18b90594232891e686e46a5cce4869d808db81c8938203bc5c8f3f6d3bfb267ccbdc033b70d86e793f2901e300bad1f9a9ae1033b61550b4ac4a6891f31513aeab10212aa1be6bc1bfa74cf3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9cdafa1ce3dc19e9a5e2d11de5339df8f9ecd568f51a0b3c0c67aafe3cdda7b71b82cf6dd2f0ac31e245f37f7ee1a181be512b2feb7eb5f6f8c79eff60100c124c49769c9db367017c240c33feed276d0fe2c6c52e25570c6a0bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3247be50b265ab075056f16fac2a4c6775336ee0599ff9ccb2d031aadec1c8c031f67de5a53b1c74a323338ebb3d2bf08910ebf92fc969fd3d4c7bd2f5b25dda9f6cdc33e31ea2aa5e83f17a9ebbce12574eae6d67a4a93aff1690;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198a6b4f332db049d4e5180a6bf06fae04f665cb908865f08cbf2d70b033477a035ded24cea28cdc7d6ed880e31fd17bcf3e0068ec50a9dfb7d9d8f9d6f110fafb58f1d5f8100f0a9c769ca6bb2e49d56d4d8a07d0f92e7abebfe12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4281465983ec126771a02eb1f3e966ed0f9e447485b65d0bb89b5c0218ec5d316931afaabad46a251a85e8a57be5a5389ce04d39089b16ec4eaf6e107cf6104d6a8ee8dfae58c3264f5a35fdcd1216efd31b623c8f744d6da22995;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c9578217aac97163bd3ced73e425d4bf051a6c4f443e54589bbf2bb9efdeece8f6056f6d97745ef1b84f97a031d81f6efd3cc1df34413d042d07f21478d21ad1e9f084624b7a589239903b0f23fba5acf59d729607a20549c18fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141a6464de9ce497c2fd4c3fa77145fb8da8907fc14313bc4ea440ca0e4e051afdae7b63ff8558f28c2d78ebcdceaf1c4ac925041e0a0fbc7aff37281b8f62113a89a9468ebd69074930ea8372e25bb8f6598c73a706b332080f1fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc429f07c4fc28e0bd4bc45eb9dc7855d46c74d9f31096d8b0b7fca34214acbf94770102a8771faf5ae8e79edfea92e67303addeb9a78b65adde12a24387bc79f8cb0216e2b4aa27d0bbca86749b3a9f0ef50e3763d6671be021734;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9350d07bd4f16c0d04558e52d87b4fbe72544b39458ad642ab5e9bbfe3b426d77391c2d78aae18408253fba29ab10d6ae3802279a82f6f89a999074a6027a16875f4892f93d934abee301a875f6b494e3d450f455cbac1253266af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1defbab2236593e27a2b2491c768c398954cb335442984eb82aeb437e627c3bd63b0455d8528ac6d38c3a5c120693b1c8b2b49620c403cb6d3e8f2ce5d2df3f1d7e3c1bb147ca62392ef144c6e2aebef049b193ca6e03c4191d430b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1471ebaf780e361ef809d535ce3044dbe3b9dee40bf7239384fa3692afec4662c3c887c76f3922c6bb3d155ffe29a4f1a3daa03b47526e61e25c63ff6c7259626452fa89b6ecc012ada828bce9966c29b4b3ec1738c0225cb7db4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1626a5479e9bb616e02fcc55e69b3fbc63a6a336e3bffe2a986362328365214bf3bfafbb2ffa737bc3c97f996482143021e0a1747c996f91faa13e1c98172a4a199d2bf7e66c8a702b7f984a7fe9f7ab5b1b01e499120b41b19777a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162df4af7676e30e228f2eb370f89d91d059da6c71f9c21021e864d4f4234b0c605ba717aa8f4c4a45c6e2b7895dbc9b1d30455da0ada4a4efab7455b492b3a6fc230ac29526d68c59e94bc7d5dd8c438f9873dc6c5207fa5d2a4dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9db0873bd912b5754f2c77ba787d10dee2efbbace4e5ecf4f169f655826105e74e89f12e48698cf1d6b4187586d2a69d9cef1d756242eadfa68aeda269e863f7d9d4a622c33e3aca6de5770240fb8853712155a27c7b45aa60ae9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131c02baccf60f027c53d77bd09d9ed0fcad54742739316c6ed54f1e8e050c433db732ca0cfc7ed47f30ca2f3fc87575931271976e1ad9c6d52e442f6b7dc6962c44a3e4ab8e6a646470d455244a5db8b25d8aee30a2174a675fedc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e9c090f89503816f1bd9eb1d907d492ec4c4fafcf04375224803066744cd2861eec822a1a80c7e7f82e48883df21256588e04f65a1cf5e86f51b04550b339ae8f94165ace1f77b17f340815ca38894551cb52552beebd8d0874b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc3cfc53539d5ae5613be31aaf95afc85ae17385b6c5d44aa379cad8d1fd84cab3644f14a3fe983bf29d1665dd8a2d8952b82254085200e6dd66fd959969ac38a23c8278ca70879b2d0eef44d6e3c0e074f4ad10fd15bc6b8d95da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fb71a0b77cb2aba2651ab0803dcbb2f6f0b97bce54bccf523460dade5ff08d032b7a013ecafbfeb86e4e54ccb8d1b9e91d970001da22ae05ef753cd44a92c9fd6fc6909066cf4ce0296bb0acaf2424305dce00dcdfded51b58f86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12062b73379e64aa557bacd6d096fb268a3c9ea60dedbef52e084dce2124522dfc9aaefc4fcf6679a456f0cb220cd55b9997467d3f6b6065d66527a7944f6a7c3d76f39ecf587d62d22d87ece32e62543fd6ee2965127998604d247;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bd5b395ff8d1f64215e8696ce7e5bd43af6150280c3ffdbaa0ded5eb24028f62c79d73b11f6b366624a751e5e26fd6403f22be56d47637b4fa09c7433e2fbd5c3e9ba66e196281f74dc53951e72873c407bbc2a6e2357da3493f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4017b63ee3865c989d06d9464fa933e53b6e0d52f9dd20d183a6f9c310a252ebb4b94b4d20ae42338850b3951a8a6f6a76622f18970dd3d0e9f5bdd5d0c7b65b8f1cb09232c7246b7585db8ed89c6f7a849063ee5a8ce3498cc3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17200599deeb4cdd64e42b651323139440bfc09e2bfd506308aab163ef06e06b39e506d17f765be968d4e74c67659c8c1801989664eda0f1d67763074af8f479701d717e52eec0ca79517ae1eea1f9f0b34b3a2e60081e607e8ce12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17af02abea260f303f9e56f203917f794e6fc9d88691869180d119e64dbf86b770b624166ccadd863f346354aa12c336b11fecf969753f935476f479b1ee61dfc528056ed95df2534fccca3adf1a17693306b62fb714b63fbee18dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2d9bd094c6b9b4dcbc65c347f54bf79737bfb3515c3452326cffcd26f05f7b6f9e0cee05c1b595300bf10201e787898638975b7dbb3f53fd76c25673c45077b8695993a7f15759ad639b7322a22399526a8ddc62384725895912b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd70b3099cb12ad9c8729f3a8ca359576c18edf0c656737e94ddbc1cd31e9d4a243af23ab8c043a82921ce63c5bbccc65ba9e9cadd32665edeafccd1ff4f2fbd83447c94947dda6716c1899c57304bc5cb9a1bcce70b28bebdf737;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c391d8d0b4af36cca80df8499e8a1f9ac7cc4f79f2fe382c8fccf387c3f2e37501c0c6833b01522dde042fe6010bff50b32f0b5a285b0d861af323f4bf9271b48b1cfcc81a9e211e5c00dabb0147282f2f4717a9d63bfc3726ba2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e391281748b847c4421e61eb00ee77ff5ea73796d3b9de078b36d08e8ea16a127dcdf0d0f496e665f2e633eb50a28ad8284c4e50fd7115671c3063818145c1637bd605cf0cb33af9e60c2e0917e25bc6182037074b85768ccec516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d92b7467dba7a9241c8beb2335bc64cdd7cfadf77dc0bca37a548075a7d6d42b60c24310530ded1a8d97a31a7e401fce960f555630550646274d0354439a34011707b6bddaabbeb1d43b00229b12f1476792bba4f7b318dd3f4f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e0daf1f14881a0fc70d2f61f863c8684bf012938dd548b7ebaf87e3eba27670483d1e1773d513a769931f943433a2ac6a7539286fe4e9fc1b9bc926ba6ffbae59b56eb60744627b445571635f21af632a466e30b70ca7fe2280e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4efb4dc9fbf3b2c90c67cf7c18e9271e34833ec664dc44b19e610d109cad0e46204a00e192ec98316acc4f2397d423165e4e7071850683a2ec2a458848354fae6ec91391a6c934d037b3a73631caef33a3e83fb887032ae76d717e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4633e1948752530cb8ac6ae6045350b92947d2f317812156173c5ac06637787155e0485523269c765f4051879b9a82d2517676dc885b4975f25b44efad72416d99b83867c043419e1f77e4826f7823b82b6ae722d22e633d9ab50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9d2a7e7366466941aa6f69bf2f6dfb074495b155dbbc4c43ce77ac5a695201532c7eb38f36a15659b904fcc219cef7b58e055d76bab1dce1a309964ac309032b601da27467858b3772a4b19c7a6794b253511c89b3b2b8fb629a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5a6a90c4fab774871355c385b841aaf70d59b95889c1a1743c4fb7d0a039e696bcb2b73b2665cdf3b92478b8fcf896c2cee5ba5ee1353d4c484de6b01199b773be90fef5038e7c6c08f000e9e20cdecf89c59484784c2fc86a5fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e7ea405025f8a6a0326d9024be63457897560cd1dd933e9e491c1df3179df13f661803aec0a16c61ecccd855b8983d3c5406147ff62ebb8c4711b02c77b14ec864b053baac7aaa7bee92758aaaddca56ae14f4973dd6531683d06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9e2be02bb4cfbfe29c544cd6ddb2f7c3b338a5ab052d3df8b25d8345a1e5efe8cd0b3211ef049cf35bdaaacb6d74cc6c1f55c2898f10b5dec87aa905c164ee54042b8f9c3c50789809dea1664ea17d9861ec2481cf66f13da69b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139d10f1c38ad7de3a05bfc8ba4ffd2ea24abc049c447f93ee52205cba9530e8cba26f64e74f7f54fe97dd9239ae75ea26f7a10669135ba88d250540df312ace7094c11dbfb7199130ce328d5803791cc4902e7551099632e2adb8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47ac0c21526eb9de06da02d7269ae241f8541184666755b998d7e0a89dbf9354a2e4939a54f92d595fbe2d16c2cfc40daa61a5f23923885671b7fc099ba6a41e1b3da1d60be50b6764992f6f53d36de0628e5b4a0c7f3ef6a4911;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cdf9370e45d552a551bae38efbd7820d1d484a873f3883cda29a793adbd4485885af1cbbf1c3ddb3c125fe94f95f4ab991c5a0a9673bacadf7786dae48d3dea13d8541420ef10696bcf3edd346df7bea6fc1d10b331ee94c3ca6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d85f6edb11dada4e765718995315520fa0b41fdc32d27a0ac10f7fc639889153bc96666fb9cf2b3c5cc2a8cbe13b4853f35e31557fa5eaa60994c5efab18441dd69a817f3cd11d9cd03cc073e66e94f63c94d4432577c312baa33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17739007cf99bbcbea4d378c3955d5bcb9b54354f3062fcf3f140db07f53e105383685048ce48bb2c4bbf395db17e394f6b9112c04655034e04580c688882a333c961c67801b0187707925d124140a410b4d384a7e61b2046153d01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f19dfefb9e91e6f270f92d2c1b43e554ac90214e23b626d21dbc113e38303b5979df892548a7135173abba8598467a51864fc015c6798367fd439f9631e423e375ccf15959ed2f89474c1e1322ea561932b5f1080600adb7748fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcbaf047759c9d60c0cbc241d6bc20f65a184758fd1333b7d7a0e0d5b92e04d7a3340e510b8f05a948135f138ddf9c84d9af1c29ae4dfd963d691138b7b499b98ac9ad848a20b54ea8b12abebb71f0ff5fe5d1493b70d60b181b6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7d4cdbe7af179c59e389b66f5fcf69887aaed46bb69eb211cb1f89f6de55b33338b696e6fb97e0886255d72ec62ed85a9f33c4c43fb6e9eb667bcdf829da31ee24333fa7a952a0075b9caeb265b3a6d4129190d40618612561f94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a5bcd8209f4e484ee4184809c27fab9da3f621453fcd8793f862a382d8657e320045bcd4277612d7a64b65ec802816a4b02a6d01d451a58a0748df8c2c2bd1015684f4ee2fb6eaa2cc6c0ea2054363373f6e81ec8245da01e088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae77051d91239f588bde6b66e59ccddbba402cb3f1d8ce27f0fcc6c85a2d1b995da2259dc520150b87888c35f518422ff6c1f56883a2d816fa2130c52f5dc3a2e46d5c41757130b2ae4aa2fe88e671b42f7d1ff4d9e1622a3d4de4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13507d33a85dd4d4f5afc85c373934265e7e06b6a2607719fc0381472e382c4066c718aa7748e0659968888ef9f2631c5d72bb8c7b4089fcb735a30b883ee5b85499e3bf8fcbe83b48189a66d440f80465ab0156b1186cdc9cc97c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e72569a7338ce4c7a1283a87ce47eb335a74af23ec6c752411261159816531a02ee6723b06c8a4ae5cd17291aae6c8c980ddc9b324119fe876454339bf3b0b1c66423709600563f34bbe235d6649a292279f891c03fbe9fe7ced74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2af21ba5bb81aed5be5c5993cf6ed88441fbd280859b49d81a1f54a39166ec774bff6f3056a147ac3af69dd81c0d647e74ca7ead3bb2f828fc32953cfb3f1a94a9c8774912bf1efdc82209ac01fb7bf67c456b16be46830c430ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1365f191dad993fe8797206f957af1b114b0e3ee7e1ed0aa79b0f374027d9b667d8a75c9cbbc9c8770a7e03dac5f405a3a3dbf5a5ca5ff76005e3176eca0bc901559398601e21b1fdb943158f1f09f1c691394ab806368eb460a085;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aec12c87ebf8830cb79c5ac548187581e609c42dc3c8413a35ed6902979a7d9df5653187616b23f3511136bbe09b268b6f515b2d33ffb3727fc682eb5f7d5db618b65d7ba7b16b54727328e0ecb9ea5f59106f354801e87dc614b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ad10939c61d1c95f5be4e00e92bdf437b63a788fda5a110ed4dcc52552cc0c439871212fb71c5e8c4a7faa87d6664fd2a60f72f5200ae0f885d1ebda32ddcb24b1a2f4a2c58d35dea432b39cf0407715b37c313182be76776e523;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83d74972b9639c589e2057c0cddabdcb97daaf4fea4e9f54724570615c0cb56138ed67f685c98e4156501ee6dc8f8bbac9c2778932c58ac7a6285ca0789474e5e2f85dce7240d7314c7f32454e9e718236ad47d275222026ecd27d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ef041ae16a80e69acec37c4fee6a928e1aa008eabbaa74203e7b52f1f76099bff142b88e8d90d8a260559b59bec5026f5866c054ed70c5a3162c01df52d708758da3e5020083de93d5be10e58b7f1cc165a54077f93fd8b4b03f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1035f51df4cd7d4c5d34b7e89f458dbd574ae2204220d1bc0575382bf891a14420b8c6ed8c8cf39012a11c29665e19bccc768ec49d6fe81eb30420e52664a1372d4ad66ed35e8d0848cfef403c6b5ccc18e383925e7a3b77f7a8295;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce590276f611308c36880c821126c9dd67be314e96eeda71f506fc134481a62ce8359c6d617f4146266b8ec38531cd14df1d71b9090dad47b049893138c572a118104b926b86a8106f2997e2067d35ec345e408dac9444ec7789c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14beead1b904b9824fd2f051338f84534c2b93ef12f1b82427f25cb236f9e258cd27ca82e6208860710b1ab13728f6280246d9546e15fe67ca1ae26f320c3cbab2b7515f4f535ae912ff7f48037d33cb74e7e63a94bd305e340dbae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166a3189e2edb4fdf824a846e1befb931c9943dd4a4db15d7f40dbef36eaf7844624cdfe84cdce956b235cc7d89e98d001ecbdfb626d388985f3ac03f7859ee7b0e790705146a98abb2c7f4de5d836d59611720c464dd12c271d088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf3e5e880dd32b47cb3876c9e6cbcfb4a2b14e76bf9050ad90ca1a04e3e689c59a907578dda904731d6d2183e735acf601fa68286bdc15f20024473c7a2a2db47a0cd5a92bde9fadf23a1c90b11e2359bb6b195ecdd30cb897d732;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c83df500b5c899cce6f4dec2b3059970154818bf7cc00cf47bf3b905c0b148b96dfda7489768f1b5291c7d8bd9a991d0c965b7170f83ee3ee4793d319d44accf8ed106f7c5c2e80db42f23354c4404bd1aa3d8d5628abc18cc1bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17796fc01d10941cf80a37f5f31a3b86b072a5619be892e3243a5df9397f9d0e1ad2f395a9e16fd848167006fa8074e18ced128bd461dd8b291486d89a0470a4d5a3657bfdab5c6e52b09566a722b44e0569e5b250568ee28b0b4ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d304add4ebc90b4937a7da33c7b7e00e60511d903d309955fd886fb7481a4a28b8c7c1053645b677698695c83ffa5007ed886e5ccb079782bd39827a295d673a74d08a36b2ac26f48808037fe32f034c97c5572de52c446fe590c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc7d3ad9602ad2bbc6a30b7dd2be9ee2e421f146c3dde07b30d63c17870f0c8033501b9940856fa881e4837e3a7f43dbfc4950f619931af2c2b968aae8642896ce79f2e45385d01b5b912c7a9c0ecfa46d8b6bee40a3889c8b3e55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5adeaa87876439c2e9de96ef3662becf2074ffb9a1b9309d2f61ffefc2f549cfec10cec9de8e7cf760d96bce18b0380bbe3232123a929fbd285bdd694eccd71639ecb16a93a67144694c3e15b8333662968225dedfcab022e25351;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c2319d74f9a8b58a440fb1a7b4a060b6c74dbf8906bf64ecf48993f345d586b8af6bdd5f718595600bbb6f151720c0e37d9fc5da4527297db7d4cbef9990dc6f1654e81df7562014198944105e944911cd31c7faea62e3b2efdb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a4ae5d037775865f2dca1890b21eefbd10b1ac3b2bb7d9489f2a6c687491fe08f6d2cddfbcc525b05ca489a43a1bb523fb31ba227d5b31c3220c0acb5f5b0a6af7d4908de257ffb7a4c170c3f9711129a31fed49c930a0e8151d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb800377c9f478b8b55974453c0d652e42ecdc2164d1beb667a9969fb9760623529230b3384668db618b0dcc30308d6dedda139f47f3ec231b23f3dde884e4e6cc973fa436b56052eae3de9a024266a03cb69e2856fb4837ad075db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133c81c4065d9ac05ece636137ca7e498f9fde53d2c07dfcda0e97dda7e083bb7d7620de9ba91b35c516c972f328d76824c2b29fcdb3ad6aabfd5220fc17b09fe2dad3cf010ab28563f5feeb620a4eaeebfdbfd7d1711be1bc0e7e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7625b5a69735f202cc9c80df1dbb5c77a6c5c4e962da8cdfdc6fd76af9578e691fef59828731ac1e1d07e821d969412883809ba33e02d5a0cb6430f3105105cfc97ee9a43ed93a200eacb2ebff364fb661a3450601b9befbb64a80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19748fdfec73a3698b2506a10ea940822ea0db0ce95fa115af673a2a6d9bd4e0b150876341adfa293fda4b043d784278add74328792c3b82220838041727dac3cb201e180dda1202f2398af5aeab77dac511c28de556750e4f21c89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde4019add9dfb1b9aceb93133ce8c4a2bceba3355cdc1ebb51905dcf40cdf4ac94c8389ee60c4cc030fdc6e3774ef6252b7d87bcbac7f9c8a4ff0c98f3e1b81954a330994a60afdd777f8da9e6ff151fcddce8c35a539fc009063a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db5b017697d53e47036f52bc63c26be470f9d875b1c0b8663336294f66138ea253433626973be9020d79021c5e035ae3566b90b68765e2124d80b0eda71fd152325b64a420ca427c8a07773f1e54b906a1c8d960805b19f6651066;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1105b124b997b32cad14f187aac1baa024fd53f3f82850ab4580c2e5d9a75e3ab9d285c65b1500de93bf96ad8ccd0450d5f7c49a22c49065f9c12b7339b92b8a9640b0bdf8b9e20260ce6c0baf1a16af18497533dbbbc648ff544fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4961ac292dfdc21be051ff6a292fe49ee1bc07cc0c9886fa4683bd1a08620d38c76f53c4ff0e1674ae447d61b47f3c4d3bcc18a7ba0c9393ba235c68e2021c9d4065719aca3adefc9af0eb8698192f1aecf58a8afc8ea9c8f0bc58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha413c763f9bfa5e92c8e8977a1f6d6084fb6ba925f66dd547ace9c442f2ee22b606df2b551627b4e42b666be5d3a48d41e0bda1b1c6ed014ff872a83b7b6128b5c4ba53b3c26227664fd23fb6622da0dc9fcb2860d2d09a26826c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d7511eb0c7ac78b1efdbdb389a58aa29dbe1d9909e1feaf665fec55cb020ff18514131880ad622b5cd29931e12766d3adcdf54941fe69b501e261750818eaee48b9c89d0edf7334221a0e6f14c1aded58b9901031af79fb7ea043;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cd2c5ec0a46f39f721da02b325fcd322e99b2349c7b96827841196bb0b6507999ed7c7ff4c564c164c884d0740fad330563a5982ed73a9f59847b3c192517f71c3d871e057137be06b2f9a7af6210f1c8400ad1e75dca1bdc396f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f95263da13f579bda756276239248d5929615f11ade42b1f5cd76bf671532722b4c9e6fe829c0bb4811aef2179aa11ed0946ef741e5aef942b2c81c93b505f8969676576a4bbfab1238876c72dd15c279cd767f3bc78b5679f649;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed875faf91c940c9f1c6c4fa79ae78502cb669511e663cda17321ee6b886aead300e79e73b3ab06283f8fb7b4b11fc5b5e518ca4f2f482438b821ddceb644fdb989cab97a00169113fc104dfb36b26b20350beb15398ffcfa13b0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca466b2344c1fa5be1e0eba13d8b983df25f5c71f10c6cdec962aa3c9f8b1dc5a7a09f9d58c857bbe3e6450727b3c9916b8a2cc3c88c0131fabc95cfc2238bbb0663690db50af17c22df7b3c67de82d5050bb1471685c97ee400dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had0170f3e1c49b07fea92b80ffc5df128093787d1e9a148a99d166315a7a11adced8f4540b049462e08ce252a69343c605119bd1e348c645a384e7f2e73545bce971928e258e1742f38979426bbae5fd5de1209ce3d28998174262;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha35367633923bb5e4f41d829635cdc6a03f5bb754938d420db46713a46e55a3940fa31488e60fd28439bdd9736c13b3991338c43b8ad508d8caeb5775f657afdcba22dfb9f54800a8cec86bebbc619fa62f7e18b65323e40c72a3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f5412dfd325640f07facb660f2d7953ca56cdd8da1e60b6774dc15411101b6875e28a30f2b3f55304a1b42424fa50cfad39e4f5cbb2a84237d286a02e97d3b5a5e540f0f057a349e9c9d8c13a579edb55157a1cdcecd5d35b45af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3430ea87c87b992a13869217d70ae30a8b4c7022341dba8ac113efbfa76356411224187db5c2c3d89c9cbe1d68dc1f408baa5950bbdc006c468643ec0b1a42d49f5e6a68e82bfb40c1127bc8a69e1bd58b56b5dc1d1f6fed5f65c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7193833013e79f219051e5fe6f07811cfb5cfdf9ecb2dda601e454635bae4b88f136f9de117b70539a9c55efb296d34e1a8476138ffacc5b32cf7c22ebc04bbe0353c62b36f18c47099fe70844b4edce51f0c3c08a404cd3400491;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1faf1ac954b726953db8b8cdde489fef4ad554dc2c0ef1dacd07a8bff891531ec12ab07d21a21fa7ba532d6428490ab960a51332cfea544abf8f12c8935f5f6d4c3aead3a4b285a2ad6e4e5a7c50b33c4bf6944aafb10bf33590192;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdf95295974f3fa9bef540b213fb990e5be83d145a40308450c536e6a505a552084312e2bfbd561667e3d0e5ed233a1f246ba37778f5fc60a80c0517134e640aceed4f55b8e34813725dc33a7099d81fe534b6a23822f669c7adca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1670479e7ac1062c7574d769d22705b25c7bd3e5868db3acf9a87f6f0af3af17d514ba91c9c092cb2470998f34f9f73d4b3cbbf100a8884ef4e5c239244a75c32c45b76e36428517d6bb9ce4457e83469599220f84d5f281b32039c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70bb809073c2bbdfc4b1edf3ca6f7e8d32cc4104af94042f711f2563e7643e774d100ef3c8ddabefdf9a8a31ae80bfc099bfe10144f9ad5eb6fc08d6aabff8c69d1b3b23c61ba4590257bb0852a03b40d31a2ef199be443004ca6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13315121d96e2757fcceffa363a7e4bb3de31895c70e195c67418fc132d753de7ab5b01f0815758a8a4a2ea5ef21aaeb99a2930c222b795e739534e08efc04e6bf872da3e3b955aa79578ca45227d032a7a63637f716fde4beed01a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffadd66fce4c3ef8d610506bc10695d20c0b761d2730a5555e06f4119c243c62ab20f2a6228043ccd538f02e94d630aefc77f2e220a9dc74e60daf6c962299c3bf7ab855bc3fed20fc0896ac608f812af5e5e879ea94f5c2aa75a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb174a77ed13ab0c82735839a1c7b3b28747f501b738b8703041d266b156eb2c43339f3345722b342e18ece2569d250f9d7dff4a13c710ac7ebc7c4e3a0bacfe7f32e525c899af9dfef29c2f5093669dc760c28faca274e05c5ad4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f304182e388e7dfbeff496fd129e444c2a7df40d66a150b4bafbc57ff3c7bc0eb56c964c3632d201c8c6dab7577ffe3ddd52bc502b669c4ee97410e4ac660c1fe170afb636c8acd12174f729d09f9195f238018e5db6c81e86f051;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156b127cd895b0c72192dcd54dc8196221ea8ef47e46aad33133c1b7f096ab5398adad975cdc7a24538f38568688b874e504de08ef7a0c15ff091719afb299ed9d5c848ebb103ebd417fd663e67a38b0897dd77d1bf53d92e4ba084;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf24a3c54701d187b3e424502417b2afad2b3716e232132500d2c0058f01d0868225d8038be77ef9cc3cccee8efab8e89141fb0be13360619cbc93d33d9ae0c4a0de19a94b30fc959567d7f52f70403d44c7e676c0407fdd6ff9fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19cb6e1a1992243a9d4fb1b1cf1be88751fa2f21d3a0bd2218cbf181366976acdd7bfae48d5618e2e3ce3895632da088354c2ada7435daebd3c7b5ca57471aa20bac5e3af7288e0b6f84474d8bb868112bb7c3b2ad0d1fb62027f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ad28baf3bf0248cbcd8887f429e02f69672615787a286e18adeab87d4b9fd1d9b914b6321bf137535c15fe1c966edf2f6a7397ca098d84ef13f4ab8c5242c9462d27ceb2c9cd201372ae43ea8d822446d08e0e96a2f71f7b0a969;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87e088f45881e854d98d0b97873100b6b4675ad50d155dc1663e70e9a663b9cbcda50ce89729b62720fb3d5cd3d7f15b1e9792758e34813059e5e0d554ae8f5f497b8f4984fc0b902e9625b306ce5f40af7d1344bddec5e82e88e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b402a8c941031426d4b232724d3dbc21cac9749a3b0bcd28c95b69f1cb272a8eb29fe0095daec4a461a37809802bd2e32c0ff359d15566c51f1f50f43483823e0dc9f3955dfb6d084f8f727ca13d4c0710123b3afa29bb1ba4bf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1775d12185f2acd3216cdc84cc2f0f09519fde018f8304524573f6348204ef6d2ed4b8ae55394d3269d9df3388f6a7c0a9159a1295af0d1bb6241ca9e0e8ab2693806560f2a8caa276c42e94a30641f17484e4c7a0907280bbd527a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de80763aa120f3810853707834930fc1b0dfd2892238ac2ca030b66676d263a3f0205e6db81908dfd2c956379138b4c5d11a036f9aaacd3282de29627b6e9641a3d9876591296fe969920ac89c258ccb1e744465972bbfb002b90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a4a3a710ad630de52f5e8cafa70e29f96e174a24d8516ea642813f209b1eac6a721ce10dec9fadc139ff00402476852bf94e814b9aacc14340b46e45a443982f8ebbfe5086a07a157b34fcda2e1ee3bed05f2bb4d76d60d96e383;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b284ec8c663becd58eab949ce489647817cb44387dec791c133c8349761e807351e17e242711ab7051cd9269bf1c7f8a00ed28081d806f62ed633b31b9cafcc91a2b812f62c927f0a15015de132c6982dc27ff6c81ea765e9e0539;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1133efed1efb62031383d964fb620b367162f831bce49055a87d78d2e4040f08392b82f1e2bd44f7bfa00af7a2b14c33d08258dad9951390e6d4eeff5fd098725129715f17d2535b1571e3e3f6ff7f99d3c04fdf0e1ff3c49aa0a49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cd62b5502768069fce92219907af93ac5d41d26a4499dce3014bc99c5fbca0255629bd93e08f07b8d7560ea383a1b9868532a4848f2e5dc9fe1c5c09ce4dd7584499f0b89829a0cb29354454a311b968d25095c9233e3c69d4306;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36dbc1b6160f166953cfe2e100bb27816de4e2e75672a0beb2630b4731c122b3da5ba74ebbd8b7b9de4080b4150ae51f93e00bc15c683de81e3775efb849203743243170d23bd31d5e2b3343328814527eeed4a35e192b068f5135;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53cf361be8e7fe7ac2bf9d525eccc2dbac3b894a5db1059b0244414039cdb126a21d09561a1815d0ce644e1a4c3cb2d4f85452b610d936164e9add1f078286cdd50806bb82fd6206745b90cef60d038b3f5191c97e37442d10aa32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c6994747d565e11ffe14196e08ae8186e867406ef10c415feb31ff93244a80f081375d5ac656910afae7fc6507024f287d90b4289ab799e28aeaf18f188393684809b2fa6f798f74b0b6afc1f917c3f3f8fc79d6e3f964592405e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184e33b8eaf6df6a553c5d710212263c385000451b0215dbd2ca6c6458c4c4a1f6ebd5894c143a54d2e238c722a51e93b83fd815d0ca52ea8c1ef8ab145cf66e6796ae0450772afaa3b773e9ed6eb4301ef84b71baf64862b4813c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10dddf316ba1e831774dee739fbfef32c5b5f7d2ba8216c8c1225ed2045fc2f573a701cd12f7e557b02df15a8c7df8273a9fc9fca0249a898ae1f9f483b0d7bba5730191534b8ecc9ea63e3197649a283fe5787e9505d1a0bd1678a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47e054fc0799f0832e04f43f9b85e976fcc1171bcf2cac9002db651f699bf4480fbc50b0dc6e8ef36674b3c496af2c3be3a948b065656a307adfe808846d394158987bd84ffa21fa960ce503fbe9e97013ffeae03ca9d045fff88e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3906cb62b281f516f122fd790d0d1665f1973bd3c90166e7b501c7c11428576d76241a8aba795b8b20a1c7a8e961cc5ae71664a6f0c1ffe2fc8e55f5dc0e22de6a3d35c5c1f78cfcc373436e13b13a658e2ecb2f22854e4892ef3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h316b84169f77c79ae6574e254a432250d65fcacc240a69241911f5aad73a20cf91c59de9954f251762bc36f1f2c958174f8311b2522872614a503358ba4dada0789b9cf23ef68f5fc2db09dfe77357a01d3ce39fd9e20adee45e65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9fe89351628d0dabded9ae9b0fb3d09df0f6c2cc7d0a15d9be94ffc49818b578ce7e5c7cf1eb8d06ea6cd630b9e55520c3bd49921814bab19605bda4ca71e462f9fe7c7a6cf7debe7c758098ee7574db5965775d194e545796084;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffe846768fcb955f59444f004d2fe91480b33c544241e021ec8a7cc6d0c855b6e6d2c73eb1a26e0fd50e655de4459d90413c44f0f7a6dd11aacea6f151d7748c87a1bee5421ed7feb58fcd8d0f6021dd620f37db8f73afc02e3ba0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123c531d3580e451709facae9aa4eaceedb9597cff9557bc9a135edc7e4a2310dd81c3548b2aba620baa0956397cfe57491d5b040c45ef0d8d0faaf5aa06c70b8685e5e4af56c0ccaf2cfc90de39510fa91221f9160d04ceecf8a75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8cf359289fc03238c851ca9301d9cd583955f1e59f85844428c41571ad22752bec5345dd2300c1fce4efad93f66637c2555c17f9d4dbbb8e19b61bd9d66ee032940ba9ca603836e22608c9e9811d27e6ae9aa46891878b6aeaf2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h577d9314265e4b87d56c2e16db6502246ccdc2aad575ce14926532e4c276bd29455825a021babf7289d9d0bfad7c27c0b22be9dc253d9c35eac91f4bef4f29f55dd69dcc457d5fd7e8fdef08dcee9fc32c1135ab43d80210bc88ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haebabf1676bda6de8d8cc6f665bcf1ed7d44ffa76b07f3e1d99e60b70c237d4cbea9fe166b32f9f4a81525766d6a0a9398729eb11787a906db283a97bde98e7c84243400e73e643a2c4dbbaa51ddc0024d03c5c4e91d42c59b633e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f125b1a1bfb89d7a7894ce6414b0d97b0cc4ddd58ccff6ec12e70f1ff0b007abbf41e2de1763062e063a6f96d6c506b1e2398872b0ee9771c79dbbdb3b9ac8133ab1f6ef249730ed7a613134a22ef6a4b3303924166109a770560;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37e5b797a1a3a280f7f70d612ee7842c3dfbfe34a8d316cf5f3ac119d5afc3c5335d5b634debe3645dbbb8e6a3535d359de8eac6eb9ea5917286b95a0c6dfee0953e535a16b128b82efde2fb84f1edce029a7af2b499726d461176;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64e0920c82e04a5446ab3cc66815036a6d515481faf4541be4e4d94be9b868a26fc77728fe00bd3ef48e5d70f52364caa7f9eafc7ff0eed699c5d1b56bc7be794f9a5c0a1fd5b7823faaa0cb077287b82ff87aab39be9f2f6b801;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2367773dcea4997013d8c414be91ce0affeccd3ff0c81cd4daa3a20a32ffa75c9a31fc81c133d4609e832fb8cffedcb4890de4d2637b4e4a2ed4973656a93cfe64ddb310e4b9bb2631eeab768c0a47c86542a22fd8b03d83321112;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1646b69fd2d594ab2e845d6c4452f13dea4c3fdc37778dd1f451a86338a2f90cbf3ca560f412cfa2ccddc6a920831938e49c97c2e18633c849715ffc2ef3b14fe58d5f3e3f322698b36088d2bf6cf43ad175bcbb41ea7161db8d085;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb13cb4f84cd84dcc1f3115ad12b44ff4d9c6a5e0883feaa2417f23c883dd90e88eba4c5c372549fa72673e237144e8c8d17016b2e96c36b7a5565dadc445e18562491cac70f029c36400f5076461773ae194b0f8226564466dcb10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2cd459ee9e494a7e69788b3a7747557d03b5e7268b5b2e73c8a3553c0991c1b338efc88bc8d2475d8cefe55abc73d2fade476499ab56241828db938f492d9a344888319f04411b9a6ed4726c03fc076a165120ccc3cebc1de081b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c29469c3d7b7753db15ef738870e8e9faf1c80a9812161f9ed5ab080411b4dbc686c174a599f482ffdb6073dc132b6e57699e513d0b2376688178f9e48701e2037e5e80128532047233c5d1ff02775a5851a368dde1ea3cebe8280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1802e641fde6402fde3a52e5626dfcd5aa4fee0afe8a42f8f161424598a7e6043b8460a9ba571616a5a4d6ff03f39ded60135777fb0d154628dc5b262b8d0372f10a35d5a719f5feec6756f2bc0953e45d5e9468047c59dd7b4ad9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h739a97e1ed5d23010884c72d9fd1003eaa0968209245f8bcc1130db4ae7f1e1c34788cec963600e6a583f1c18de8f00d1778093f57651c868ef03dee9e560390628c927bc8d319421aeb97e90e2380c891b0edb1c2c1878ed8b182;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126bcf25fc31cd0b8a2846f03c995b7561a3abfdbc9edcbb6a7ae2eeda4d15feb2186edc3bcdbf7a6a7392d664e0ea4edcb536017f16c42a370a713f98394a46cca64fde7e7d1bda79d6b6394dc07d37664c7046e82778e91ef1c80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9ac82e4f520e10bbe40711709e352876c48a1c15f0f19e1d5741f9a6c5d2e065939be705cf9498a14843358c45a00ad1b3a87a0ce010845af29803673b87f85752e3a7d855f3af71ffdaf3fac939825571491c6285fbc2f311a1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1d381f8b4a6afd5b97a0193cf09e2e85c88a33ed92b98f551e50e5c69b004dcbc06aa7112dff9523d6080220a82ba19b3e36f08ffe3c9d195221d2c3740b68dfaf933963cae6fa0f61636a874dc4f1316320b527469ca66776a3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca17dcca76a837f2b20d0abcfae3ae944adfc34471e7f3fb5bad05ecfdb8a6a90892eeda17e2b2112f6341e866f5e30ebc37f4cf85410b9c393b96dddc6a02995ec8b785fc474f79091912d62d0cfa8effcc6e29bac4b6e6953aae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1deef2d5bd278885fd593596d5ed38773f37a668df98d2423d14ef2c74fd460909d5c3c46540769a47e4c16372cdebcbbd7035fb551497c57d0b5ad66641df2915d2306c904983c6c6277de20102ab2c291406305e760e6b148f464;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6744873b4907407785775fbb356c107d0ffd4451eac580ff5e99fc6d9c3f3cf2ccbb09b12806f172f21d3a00407e4b7983d0414bc09e5e56f6e785c5a88a1c8685a3cdaa452fb4b9d5a596276c23dc0e35db8f014f2e18912a43d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe0ea7dd666de21f30d322de97bacf739dc430559c3bebae5f5ecce56130f381af12fba9ac1b72aabbe29de34467ff84f35919921dc2cf61c3cafafe9934f116411d1f37c9c6d625ac94f50e620bd0a362911906c4ea1f0a4a01a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb51c0e2f72c8efaa30c5511286e8dfbfc273f3bd07fed01de7a6f2648cf076312abf7def70f790be5a8d9374e9558b988a76f1e525119f3ff5cfac5ab887b2c07a6f78ddd2c520a6ff211641d5d29f25d687daa6e9b23d831a50b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113a7e77c6583f1211ce0f5558cf3e91444f3d96842432a16e1da0d0885504751a3e88b0d78fffa2ac3d90430fd3a9804b0a49f3d01f4126dd73d9101040e4a1f11a928ab759b1ea8ee00543a5cd9ff9cc714f7e5d6c7f91cc23ab0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc79d89dd3390494a2f9f84b6ade79b268f97eb62b976bddffee27edcd766eac21d9719a97e65fbc711b3b01ef96d27e48ce03a4e88d4900f7d4148782e2bd7df737be3ec2b4922d35aa060ce9a8a52fe6090d3d4a45d0f7928d563;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b44d66b7e34ad866fde32280bc8722f5875a83d255850020802994ee397999995802a3c529315d7b36deb07fb18ac427714708cf7687d0c5f07b74647ae85a961a0356eb12cd9cca8b17e984a1addd97cd764f34f6b47b3fe7ba6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126ea49f9015a086b7e5445464204378e7cd5c63b1e03d46f3697ddc1545693c2c191015b290a5f7ceaf1253be3dd759b4de250264e181b48a82f6d5ceb1ddff19103027556f04e6fc8f6ba5e8e6514811f256f373f8ba647cb5c58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196d60d0235aa3a0faa2b4071ef631da7d4f0f8c08bcb98b5423c296e4ec26fdfaab057e18451bf41730841461b8057267e6648b7a921bd36cf07d06c9ce50b1db63aeab7b95afdf5a288da9fc0724b572b7990a140a85d22d8f56b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5d250940203471c5508697c97394b5c24ed4a2468fe104d13f63353cccfa9855841aca351d818662705a2f622f1af35c1fd245ee9d24f4e16127833899d44cb1080111a0cd92a87a24c9d993daff750d996a2fc3c9697cb68a1e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h702a367d31e1ac7443e4dfb626e04e2ab658a9992a4750a6dfe9f4f7c30d123b568dd6dd8f7ad17057436a092c72948d8f98557d9b84d0e83d028cf45aaf8997da6fe4705f1c0a24368d80a7bdf11dc36d6cf2971b50cad64f3b22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b5a33580067bc4b4564aab7bddefcd4c6a5f6f766b2eab52d7b2f899cae7f5fedeb7054fbc834a0ce74b28cb3287733f0c10192dd2bc8818d120bd8667350afc098841bf770a404c0948fefb55e527f8a0136efc72f7568819815;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0530914241205fb63aa2d18b5bd920aaf5a188ca4a48f4fe7c234eb3c315624f7cf1e789f9a42196d3ba57aa7c66c37c6044e6e7a093d5cc3f4c5ddb166ec71e6b6a71f5d3d44f7687276585d64950d6a0ef2b5c6018b80e3c7b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1cb2cc7a9a39d8b1be3eb73a1e823c8e063e7b9b686f78dcbb8b4145747619067b33b4fa29826fa120e060cfcc4f938d2ce71533a63a02a51889958d5f345f5ff1555ad7f2392294720af2fc56adc3d45e552e1af158601bee548;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62f32222e56864a52892181d43f9279c5299b28eeeb3333bb4cb66659402eccb53dc3b5193ca1f63e0eeaf49f1a56333d1059259ce8c291046fd2a352eb6b39536a074d9ee6531c9a6bc6ee012b7295aa787e9d383bf01438e4d0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba7af3c7a5c1c4345a946ae7e6621cbb2c7f463eb96b822f97b546f13bf07358d7b3fb917f001a1b42f696ee7f34381f8d93434b45340f07983a29947cbd3507a416b678fcf65054b02d29098190f3c7df8fc5097bfa46c814fd4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50d1be44ad1af1c99a644e893bbc8c9a6ea3ae384e0478ed1cd9ddd6d3ab6444aa1173dc2e29ec9ca0d89a6672200106dfec50097b88530047a8f86bb44a094b3b14495f47ced8dbad9dbc3a303632143e721ba3f5bb6bcac3c07c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afd95e3e67976567d8f3642b077b87d2b75332690b7c8b65a069afeea2713aaeb05f379a36b3d3fc0ac9ad0b6b9e3d6b0b53cdfddac3e20bbcbac718b46cfdad297abf75026588eb8dd5f93c048567ef4d7caf4105b9d4a2f91d7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e8942afd7818358c9bade560d10348a935dc3cb045ee5a694d4992cff15c1615491537cbd14d0697cde81e5b706903750b7e38a22248328e0c884f582eba18aa3095d42abacf545d30064c087402afc3d13213b1b819260dc1faa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11552656b127d76a0b362067aa5b82f4a3c220543193298d96a59a48d8b7b782c5d6862a16a95eff07671c4469567488bc748fd0d3d81909c622e5c72a4cd358c8ae5bc003999668d8c3921b401a5a350ac6a173d855df815ea54c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1090b18aa044ae20d49962ecd270045951c519ab8ce6873362c4e715b13f837665bbb50f33307c0a3662d393f0a37387c13546c0bdef5029cc2222b848e91d603613f4709541ebb8753798128f6a30492d478db5257e4ab84801b27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b6b53d0029bc7eab9c20f02842417a35527319c53960e842a19e9a5a7e37f551cad51bcdd2098b05be8e74def99ac39235bcf2f77413c7f9e4ed6f60018342235498891423e6565a1736e4d3aeccb3442e8ab77a8a974d77c3909;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1084857efc8a38276a49c97443561263e62f4c67c53a36c7b1fb7ab296234648054a7bdd5270ffa43d6c05aaa43df699fb1935b832445f11266143b690dc417e70ae7e58881856e696656e00139c803ec3cbdea7107f986468f4e96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12018ac2327946ad5fdb51d29d0ffe4e873858a68bcbc3ac3e003a4e2b089d7e29a6362344c83280bae8784ca4c4f669cb0dcde1f5ddfaa9fcfb0875323a6b9e1c5c07df10c862fbab5747b9bf797b917c164d5cec4f25eb275c01f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc276314662f48dc963bea59d9e295dbeab6e9d54d204c9a50e2ebe1ca5fd317b5f18b23c18b4dc7ff011541b534bcbe0b1f4df91dd00f8eb6803c75812934a1ec477b76a0fbd9051ee88665fd8838003cb62c0f640ebd84eef975;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6365169b67fec7832a2d22b70b8f77f6838d223658381be5742b10dd3d89cb91b5651bb0c742648ba48948294908cf61d06ab0641985207139053d10a1ea0ecd4c87a0035ad5345cadf4c3757dd946a0ddbfc180c3244118b158bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a48dc44b4536b86a306b3d814aa5e23de5fc61425fc299657a080a2544fa5a7314a9ae01f10b2567e09ea622837fa0430da54ead7ce64d92792e302f2567e9536b3d427307e3ca654eded880617930f0cb14394ff84a5c62ef1aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105150d2eb30e0633b0fe1f774d4b5da12b6f31bd609782ee48c4622035acc3052a17c2bc8f9693790c1575a81494ed36b6be304c4bacbebf2b52c04a72b4bf7f77874b96b05550680048327b4d67f6a6b845e0be559d0ea1874f06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d109b3ebb46a35838bad9adf07f8d4d00677622c39e469440b40098d40c91433d5bcafd4a7689ce8860217bac976a695f0de00fc2fb685880cf5f8ca4c894d56099b4bf33037a2f0d87b137c6541a8e25dc0011e7303044362a61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f695b298b8307c469874cf8951532739b5a58e6b9a1a44c422c2294838b08021323add307d8d55bc6384fd8ff1681c3a2caa671983105c006a1767fc3b6b6881d57d0fbf004aced19b48f446e81af0f5976637e83ac348190829d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76d0e48efe38d540d7c58a2017683334960d6813a3b289603192740058d8718e81e00d4e687e2151da63e4bdfe57867c381327faa36de09b067d243a006640802b084c7c2fd070585b559178a31b53ce1ef6e1afc797ac00a37a1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f51dcc5720e75663aa756832cee33c13a9b14b5f1f3862def5c73cd9ef6cbeb745e7df5ee414e65da4b8cdb7a309850a90e2b2b3559d43975681a79811a9ced83e3e11177ae16f4a2f781e9968e0986f5363b1e02731e9a50abd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1663e89b07c17f8a4d1d223b3a3c95f3a4f54db4a151be6557a05b8e05d40974603053aea4579ea892b153d247f30776ebfba09c06dea1e35879393460f9869b02621325e243be123a8e4fde327c0b5b230e8958035bef411fd02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a425af8e2de58ae175c17654636dfa86f475a43709faeb1f34b79bba7ca7ecc677cfe99d57ce6b7c4c7c2759a5c7b577002b825eb1443b9216fcd83907f9c98bc25e6015042bf910f163410e73a3fcf3fd9335c5b332fb79bddfda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fad521610a99cd2e396d0b4d4f519c113a31a5617fecad1e3b4ad5d1b1ec4a9a8e6fb2f42a1553a5cfe0d4064204737d506034218222e5421b7fecf7edd488e1a3cedc85c8467fa3161fbd96a3ecaf13ccff7ae9a2da21b5989bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6ec81e3e0a5cb68e0f6e810de579faf032d44729ae143c181b09115d0193ed0e7a32efe770ff86975bebeeec063f83221679a3ea7317d1d4a31f8124724d76ccd5eb5848a745abc515e6fb0eab3542196e213e6a2f5ed9abeed7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149fde1bbc6ad4d9d2f223257ba013ee216c738716d0e0c6cacedafc0714d405855452a5a0e71157141497ef4b0089556b1b6c44dc88c94c98e7dcaed1b72b1d1e22b14df65922fae5fadba8d245ad52cbd6619992a1b0b10c7f57d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f61fb9f75aa9a42bf3d947826ce2292fc99f85e58b277f7503af9076d2a2a3c27ca9f326bcafb825198e5a5d7520c3aac47780a2bb3c3104cddf776b9eaeb938cae667db44ec7dcb862dd836cc2cfeabf456e56a2c6b12c24e8d19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110c2fc5f2fd97c6822947103d04d1717e98ba628ea9cc9b95b8fbce4699643c69484a79575f0999d3b4b24dacb842b46628064494668bc06c87f3f5ee2d2c9df4726a0ab3d426d2c863588388b5a27dc14e7c3d9bae82bd74029de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha762d2870f702c0a4546cd4f71c862fab3aad2a06e743105532443a568ed2717502642befdfe2dfbd23f142250d6df3e80555c97e8feba1d19a4e888b83ba9f6d153a1aebb4f14f64d657fd6e794aafbe5f64946d5b9aa773ea85b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha360e7c51e3763c96a54ac6442695a22596e66c882f8dd7b1f75f880822dd7ebfe5d5040cf3aced0b8c6d468e199c1c7b0213605f45da6e22c788f3ce743c52abffc0d1c1af9f4716f92b22ad7378e98087ffd7a98f040d74fd1ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4be82a81d66388226a0f649c388403f5555a8e5e1d51a402fc019604d9783b25157c25def3036eba454e7fda5e153882954e3649ba1df668c962510df1c84eabfaab9ab9711793f842cdbcb8987ea66622d91576d36f8fbe320c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128a785252730e91135ec7ff2c2c39ba9c70d8952b83eb577dbf06a8460b7cf15438af8bb67b96de7f26e04bf68eb2200870eb6751bef18183edeede3286341e863eb5c061f87b3df9fdde6cc7a300f6eabc33acec1fff7c1b86546;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b6b7e4ba73ce753f75365702ef4f7eeb5fcc6d587ec87526afab5a66a9bae3b00ff4b53891bed7b6f18221feaf0e7d3d572d0af1b29f97a06c634023a549790a2725a6767a2c76a908c29458990b4ca88a532aebfe8a6bf64e297;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8cd4d41379efed382c33dbcc5b643682bd564c70ecf08ab29e09d1ab55b8bd57a1f33b735d4eb25a8259b234b35d512a7ca8bf07f085043d8187efd8d4477eb940e966bbba272c785a84c26111f8e77a3c7d04ceac2d6846417155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1836194f8c984f71c1613f94f1162b81c215dcfd863880318b31783d14b0e14114c1ce17fb3088fcb805d0b31201849c81640b9ebf5896dea4827da395b021cab989a8bfa07f33f3d2ae32384e1e744395c8f1aeb5e19f4b44103d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f5f7e006ea600bb2ca6dae1aad4a137cc204863bae79ef3d63e5efbdf3046d26e06bcea3a99f8473360b6f0bb425492b735b404da15efd9e0f23500753aab99966280055bcdc9400ddc9bdc87fa6ac2cb8e0df72436b24a909245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5de83b0e51b55cd7cbac446818e79294e8413be1443cab2f7b8ed7d7be4403d36522c3b4a10b70879a6bb536c4921bc0278599ab781df952dbe5abde30bd2ec82bfa56ac492c0a476db04e185f2744e891d3c8dffb0a333d49bf9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195f92538eb50eeb3f7be52ac095c08fc14acdd09c53189d85f552bfd5c597fd3de99728953aab76fa2f7a19cf0dab3c6dfc78ebaa23d5b3b6f4b6ccf00a7ea55f358d0564b14e0913e43e8f944a7cf472b578237af9ddf8fd02190;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182d439559177930de65ab41fd25284bc36a1012a9ef8b240c4945da9ab1f3fc2dbdbe7fa1dff7784e5e426aaab19f1f207fb76ad1ad2a1124e6242cc5351b544186436b205cb9bae2024996285a09c7e50d84699c8db192ecb346e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93bae544690b6abf3ba2ad833be12f7d092a8c1c31f85ec57e847ca65cf0523b05868499cf61405933a5bee264c311c4599ca82c6d4882a15a6ae146f1cc7be86b63dc41fd54f9ebc518e9c697ef282e4abac334a3a29b7cf02e50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0ae120d817374f2d07b83fb8549c450ec8a01432577daffb7c69053789ae710137dfaf119c0a2322495a9d4de889fe06f654f741923d313e6eea054819526c28747a4f497988e1c91079e06bc39c673313b5fb06c076b4ba1ecc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee10cf0d3ded4a5c03c74af15cb59fb32c3276ab56c5c66432fe99e553c6b745946e63b705a08d5b1a52d4e27d0ab36bf602a3004754ba22fb63ec1ddb2e371a0ef3f96480b636c1e436713d55996b55aa1df5c61224894589b3c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1775a5d1d7d3f185a8d5fe628144d86407b0cd2252c663a640d89193dcbf65460c5668be5d90a9332500ac3e8de128cdac7a55a5a670fcbeae74447fabc1b7d3aad703660c06986f1d668499a9e4e378d51cfdf0472dc4c5d3c7696;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be1d933c4b1628ec1c8b5eed976206ed89b7fc52bcb73b595f727a6f76d0a7252ffc14fd4e9a9f52cb920c785671bb24235985cc01723930b0668810eef7cbfb958d5c790591db9224dfd645cc8f848e8bde530542436178c5c904;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ea73d846a35c460b97985b3dd9b193f270f0e21aeedb5b0a15532f3e5953f2b0d18f89228c65bca428d08ddfc588de038dd80b9d866fa8cffc88f11d3cabdbd386cdd4cb94ad425d9319568dc7385e5328d5a5f76691603ea936e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d920ac5bf5bb8bc26de978de2f443eb2f2b3fe7ae010db547515eba2e5a35aa9928d7eaa1e474067d08f34bf52b829c76235b4507dd9823c3e463c373cccea2b87bf061d15898403d98093041327bca9c4c4d3375c0a2915b1faa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b01306545d45ec570337247c9f35b2324fb8255769dab94478c5c2a86fd48434d443e0ace89635cbfbdac2a7d9373c4ab30750b3ea38a10c1f0a71d43c9e842ca4e56a0fe1ffc82bbf369bf93d8a44f2213aa50d3a29d4abd2ff04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8de63afe50d41d1f12c5ac72b595b2207a95b7eb11435cebd7bd5765d2dcd5d3f2a0f30a352dcc86b6be8d3528f320d030ee9d020a57fc195017f64b202379c8451bb90991ee618a2e37e34b888ea0c8ab650e2d4133d11eda5017;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc8aac95cfca2dfe44aa333d986bf0402ba60143676a5f3b0ce92b3cd712fab7e3f123635b122d6d7656661dc7ce658f70ae6632a76057c88f306e0a04e548e4073794346277eeeed9153b3074263eda992e7a81f6721b549624c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e59171bd46b582de6540f0453668b733b8e5585bb59cc160501af6ade6b62cf9fd9ec3fe3d42e067fbd36a1c246bf508d0a1ad932216ce56c800c416d63ee259e7acfad25f923ba6ef61dd4bde40d320b3dd7bcce8b8c664ecec9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197ce78f58866ea501c301bbf94c05a6755d96e33d7f37b4c67b70f794aba440f524d89d140321e5ddfe87eeadfb703274bcde59ac17d71264997f11ff821940003c6d2f66091770a8ff19f9ad2c73b21633e924c2af21be0153623;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7e9be08b53be7627570cfe1e0a7b51ba5baee79f3d6ccdd236a2d8549892fe9ee97848cbb72199ae276efac3f5ac7bd292e199b7299c93f6dc0f068a117252c5348387a877d41bbdfe11e183616b61ae3c4a53302e550e23667d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9131a553bdacf784719b93c3995e352dd19fa0c69c456c5c984e95fb7530f5cae7d5897f0f0b159495b0581bee379a7cab3f2fafb376c815b8af4f534f428dbc480bd51f68ce0c876854ea6e7483faec5774c6e941ffc2c973e9c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dadd39391a1c43ecf77cf68dd784c06fe02a4b580412a82b8c759eac20bb5c9399b025026cedf5b8fe89883235d51c0ed9aab25676e1e2d6bdee871b17f7dc7904a9e9a6a892c47afbc7bd9893bdce80844ee847d5641ac6670654;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a038be6919f0f2781a081b0b2598efc35b750f04cd7ed3d1efb67a5ca4c8300d70a7c334f66340f399b52fccedc98732b05cbdfa2207dd3edc7af690bc89d340befceedc43a5f532177230821860e82a23105148c9cb9f469366;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8c50c490f554f9857e76628c515d7f302d9ebe75854c963b8ae9e70164eb6748842989ecb6ff23cbd4287aee00db2907851b9e310d59025c0eaaceaa94361c636345fbb4ebe49e2d90d514f0db0eb440a15fb7b2ef2c0873bb224;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90d648d36ab57cd2abd89cb0e1d69890ad6b51ea41d7f3fa42bd9fce5cd3c176a1fb4c6517481e52068cd66e72b944a4d3894292790d5e1fab6663de3846feba575bab8e5c4455da45de6be0b76839b8816707730bdd3fb3cc0e45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9554b089fd4554e16c65b2f1a9cc8e7b04a1e005ce823bb63a0a4c42545efd50624c1810ea06e751b3f7ebb91230b83b2048ba791ca85e088095b662c02e4080ea7fd7839c586bdfb6291d348a2c4c3944f522e611908ba4fd964e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a52a6e5057838a5fe003113daa5b7c68a48d9bf028d8c6d220272c6bd72fe0302eab63aa52795c2b403691a5886cf6b57e5e84f33412a3c5bc27490fd28e49e7d0e5925ed9da60f883f2064179275d650dd311bcf6fef2f3b81d2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba1385ef5317366a1cda3e469a9d2ab3a95bb29a7166d88a764cd1541e7d987f08d1b78acbf133b6549bb1f73611d726e4054b3a552107465efa1f98e334b0edf6cde8264a2b8d1b1d0df06dbfcb09b5c80c41ee2b0985f27acf6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c1c1a2e1234bab8d57d7af9e25037cab45744bfbbf0c502103747b47255d3bc1ce6c21b555f84531c9574a2388d2ea22b08eff198011d09481e0e865b2853c4ee33bc46af627375818075e4cca75f4f4a30840231eca6865b7f6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7df8f82222ff90e0ee28f5417799683b1d88360a107b66fa5f055b9c78856827dde4ad5fc01277434ee464941d6a614d41845df73d8ea1d7fde6fb4454e3e32d47f99265e50f018777577f46e7c40bdedf3fcbacb133b361ad167;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b241dbe0b2a1bc94789428180e8bcd33fc24ffaa0285b0096682899ccd707305b484a15b077da5a36a9e718bfdae70e386a20421c8869b79fe1bfb607b026845a9a4ec93b075923e7b70ce60adbe045b02c474dafb6cd4f624ce38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6ef8b340649eeec8737bfce8ba2cacfa328ba2dd8a54df6fb908a64798f6e7ad02f0738a84f8ce55e1f0a96f40614f2ae793a5039472c9bdad049f80dcf69269bbdebdb71d4cda8896bac318846a18a97beb5e0fcd9eb4835ae1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36015f7733e87a4b21d32992079dfa66cb8c710751b83e5053aaeaae585cd54b7ee12797a2b32cc73089c7e0bfe261885618f07615de17d631fb54baa85fc49e43c44ca5e5e912fed1c8e5774be1549147c85973f9e72f71d8c155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fa45a40feac8c2cd4665ef63c8ee2e899e6a435f390f3816ca5506ea11907f1d1652e92f03660949ab4e29a50fe8c371acc21d778932e81df50c07916a9b3d1c6f777ac5fa39e233c103b0c8b00cdc78ae66db16aac1bcbb62df6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7f6f32574a1e47c27d0eb824964394a6b6bf9a81fadc14b2ecf973a640d19c94d4e3b31e2b836cdcb31959c064fbf7d2e221aa7f4fa8adbb60a6f344a2022a582bf9dd2219d9ec7106c73b83637ea69afe5e76de0f9e55f82f09a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37c7e6eb324c96551948f7dd2d333d8ad35f7462e816dfe86e8ef56af15062b69639dc01834a62c835df40d5c2bb4a79ae37e7dca4ff1f983d65326d8bea7953907097f9d3975dbdbcd4c7adea1f83fdaa535dc12bf3a89be6c082;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1040fafabcdd56be59aaec055bd421640b8a27edec86b18023afb4fdafd514ea05ab30ccca07240345d52b11c815640c1c41cf396da2a6232ca8452e9e41f8057b2370c0bb6c1fd9809d869ac6e72bb9caffc9eb5135a9316e5b9e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7cfc1be8e1fccdffd6f7a15d27c3fbe3eb09d7ed44f8d1c99232561b8961a6a5e9a864f6c2af164b6a231be7c4a8b3cf4ab35838cabd6ddee36fbc10568070eec21df3f75f2f55a3a95548534c76b37ed06f7bb8e9e50df2d64e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1203accb120b8329e060f4af9fa9a699517633a1a4ef75d27c81d7fe970ebcbfdf6b72c5a1b533dc22668780a481bce4133792d184c84127b02b2fbc0106005cefc04ed0dac1507e84ed241b4eadd3229ae68122dda411b3998fa39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177df9a3f947802bc38c32edf14e8f18704ffefe6763fc7df91064c117d499788db31ac8b8fd883318adebe56723b6fffb5d054079091954db4eae16da235e2416e511f04985043ab041dc839f6bd4f6f647794c08eca37e43de1b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127b33afd684a4703f4785ec0815da64c73591fa9ec42172d0a578f2e31e03866e5be3aca445bd38c29fc9fe01c78e3ad3768b6573341f4a6120f57e97850fec7f704f3aa2e592a3d830e79cd8ffdedfacc4908bfd56809a3282fc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h262d3994975403635af7c5121d9ce29143c2f1ea3668ecc61ccc9e60dad8ddc9618d57acbd7f18e14d971df8c185ebb2811da16fbf5b4efefd7131ac3a5c8e3906c15940753948e34bd0b24b811120d8d0fe497376625d43a880b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26d209ed450284614e8617c60f6e8462f74456c5521cd55883503619e80ebd68d6cc5aa3aa2f8ddc9c61302bcf1a8ead5d1f378916258581f59f2adaf97c3b5e86dc513f6dc3c08b5b8fcbf5df3cf59f2c74d02866c2003544004a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9d0b7b147ca0c4a4bd9439ce4cd626166c2d7eef26701fce1c8066e7c6f358d089556c50d6d5d8cc2e335997325fc9db584712d951b4c0d092d3b05c245d34c00b06a77f56560564a52d5fa6507bd890ae8d3a1048da1557865a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c7e04c0ef64db05382d0519d81dee6549f66b7f22093b0c353613856924115093ce52a37cc68ca51136348e958a24658e439bc5e13bf39d96ac49f8c651b215eca176df479a30670fd8caf4a1a2e86a98e8baceda4e47faaf0acf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha540ac927bbd25a906dc3ce15f160b74954a016f07d1c481e6a6f860e57357e800e9d02a676e8fea87ea5cdbe36e023a7a6dcd6cf9744e07815a35fe7b2f25d4fcc06b4377e3b43a17b6935dfacb68181bca622fe3ec6a64c0705c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4293be429378c01076466ea8c2312883450a8c5a6d9c7e2789973fb007ce04aea411913a7496ef1aa8a0f935ca4e86e9f0e047b89d3c806019db0c03695ebec092e792b49cffc17503b00169e8d44ea5b224680f171a6ed8fbf894;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1418140cf9a0b009b483718a389a067a26afbed1fb02f451505f7aa31c474220d7dd56b8d7e094faf4a213f545649efc2fc6cb5d44730fe39d518267cd59131e7e3d3e3feb0af7d60116fefae76a36b59c517dd762d66895e1c5417;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefa3da06b9a0174005a994c24e9cf04789d5fa6a7a59d88c5a3160212beeaa62b9a8b831ff934d99206bd1e0a8e1466280246cbd0b1c752ef6fd574c10741c203c295c32a5fae747d67f51ca0de189b7f03e2cd0a4aadabe32db43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1a7447a1f9dad5e0e569ea307fca5805ef37d49902ea335327f94a089ea711162b9065d0fb43af7dab83b48a416549b95b1def2b185660af3a941f45d55ec9547049354e95f34374ea4d096b07d3851c711e937a15ed00062354a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ed74ceb01d88af6f31271cbbf6dfe30cd467e32dffb1f8a79e7c5a9cc85e0c3f5b277c97f3d3ec9400c4880366108b0d7ceb6b1d5c8dda67f18033c7438155b7c8e58788701c25b4d7ccc357168afdb5083245948676634b549bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a40cf47aef4cc06b025e8cc8662425af7bab4e1ed2ec1fb132c513c09988fadf82e977a6ddb35d366d21ac8d64fe04d14542f8f50a7510d6356e013e17b881b87cb9f879c3b5268990076ab9060c2c41b56cf31a528d550e4a454;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f9913e4c3afe38cf45766d30c40bdd5d6f32e026c00c0ad01860751663d7a51d76622a94cbec962a82fbef5492ff57e38755029397628c92a98d87f874ebb589020f25a4e7dd62b84d3b2f7709550cfa2aadd919730603765d2fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106ea0cfc2b738b27e62998d612066e02c07ebd9e27670094272b18bb67d884aafe5bc225d642c090e7b055f979b3b68725c1b7eb83c171cb4e17b4a7ef36a918fbe7c749e266c37cc7c6443ab117162e0e2a35b6ff2b749dd3df0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e3b5f74a4f41196eb9ac3ed8e7621e7c0df59a132c1c4fd5b12f26893274e8a8aef7a6a26b1cca6d79d161663b2ec78094ecf67ddce13fafbf824ce237db4609e7d611087bf3f04115735031a23e20f8609966e9df2cbf3645365;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1fa93508bb0c92c0c8d8f2c8031be2ed68f914d0ea97b61df5959ee6bcffb87adeb8a228d116cc970ba6915da1451f826bcfdf70b479e551968c1605aa0613c0692bb777e2b65043eb438e453b50401f536ee37b28a5c5df992c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ac162eadcd8174ca0a8bd4abd424e09b4c7ad7ec75895db5bde9072971be94e1241e564420295b0238e50fa7b6bcec2c31373986d3658aa511d2ceb15df725b22fa29725fafad2b2369da894e66514add09eec99af1a783a92a14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1961c5c01b00fe4d0e1f623f37d2a97670f168b78afa2b52c231c23db87fec97a7977e7fca3e18686664b2911f5a788bb88ece544673fc32f73784737bb3b14889a9726e867a966a864f73db8483d92f44864a60894410e96172cec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1466e1ff64780b49b24f0d09d52d30fd46dbeee2f3325591ba4fe41997bbc49ab724910464034cc6a45a5896159dbd1054377a54b8f765fd06270c7a3f9a2f3be10a45036a84b801da323817b90c6be603f6013806cd5732070463e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dad63645748332043c60fbdf61f47fa00b094abf9e09970423c20f7fa740bc370d39e6f3827e5c6e5f4c0a7579a7031e6fb79bb1aff208989f9ea2db3e7a47e184caa7eea9cbd02c65f69ae7fb8cd5632b0db2b852714c99e317cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0b09d446b1c1daa28611958765adeb039da489c96c833550ca663b25e72b45603969746da4004b76feff2b6a8d21bcf568e120c597e579fcb81ea66124046fac6712419006f1d3fe888e3e620ca7c80399a427348978d7b45e273;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9b2136cb25ac38cf2cb5042cbae4023e2142d69300e5b837e954d0e195ec459710cb0303149cb539474301f00b8fbb6bf3300149b7cc28a36c037803f200c9830c5d090ff362bb1b2dc6821ed5ff3fb1a54c769e4de882ed66997;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fe718b80892331c97ef374ec5fb4c9141af32095ea74ee65d8a344f025389a7e0ba48435f2d5c0c86080d1b7d60a35831319b905089917726029730587138f9e27960cc6ce5847efb56b88d1c49bdc2b8d53fca9a3052a4b5ed32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce7ef3ce9118bdcf50675cb6e6dcbd2dfe8bd24e4d5370d32ef6e8e95741cea32b4b7d3450d203719c23f4bfa021172df5d391106500d305d45e8ab1cd4c87b3385e68e88d8aa1c5c14fb5d633baafa27b5cc9e62fa6922c4331e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59c9da5bb36fcfd046017393c38c796c3b806412885c38fdd492735683c95f6038ec149e090029c97248b794e97c79fb5092a8e9c27694df5d85e57568a2e596271d4e8f98be8e6da66453c0e0df7e3aa13475a3e60074bbc75410;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f10dd80cf042f52480480f46634370ef96da0b6513e7f0c8480497b3a3dc5bd314f6c4717d6899194b6fe3772937481515c37e3fe4095c2f942a775c0c0240483ca15af919a5fd70baf3cef2c379766c18b8178fe854250e251d2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4629401e6e35403ed8b5f82d42f3acfe81aa3fc867898bd02c698cff3b4dbfca9d6b77adeda652215537681801692bb98a66f9bfc486ecc33d8bf76e575692d3fc4e6c0f99c0b74a82b3dbaa38e0bec77dee423c2a6a788144b9c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119dbbd6052609d46297aa4ea63ff792c0e14afd54cc038049e6f3957591a6ed4bf315f9e9132140c4e9508ea382c8d8e9d41e336d52071b3c25d4cd003d42d407cd9fc04da798149b05e6815118ebee822218f4c4b285c7dd9faf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ab8df773f6f85382746b4d6d667320d88c00a67dae25ecc32db0873b1471fa1aeebb59c64586613030fa2bc2ac3d889b32bde4799d567d21703ef87721748e23efa8cdf2bfebfa64d39f427aae603bfcf6421d188691c14f49cde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10106aa1cd07ee795ece3f12b1ad0ed7692407f40ada0224ee692d8b13885d021401d61fe1a3c86f61134d7a9e01bddd9f9e360743f54b8ab74e014705f7547adfc7ec07c506c5409e1ac76c56b423d348d983379d50677445a24b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12761f22586ce8e5960cf56f41f71f2b1edb0fb818cc7a712d5680579b1c9848d3dbef9d0e2b2dfe99df2f0715650aee015e87211a5c199847dc325440cfd2bc287894c22b54d575587867b5c721e7b903b019958662d32dd70b854;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5dbfbc14759ec88f1c4614e3c2ee39cdd231fd3ac57b2d30800ddcc098c70a99f8f70c8d254beae3b80497e3718b3446c3221025f6721eac3b02e64ee0dff9599475ded75fcb4f79fa75e2fd865688ee98edf8f899f541cb0cd3e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dee3b801b30ad70e348115430527670a16ca317340958f8760bee9d049380b2abb36088887e1885dd50f670e440c4f40a7d2705e4a66bf4f55a46613e70ff85689f4336e9686edaddf775bc1a47a4dfa0edcde76879c2aebdac1fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1364f222925023c83930e0525f9c167957b54eb304539a798c86fd8c1e9eaa10c693a3576022b76552bfff8aa615bdc33792f985b9c5fee774ee7e0cb73e39d05b7ced9ef07b3aa842df812fd1469ba29671d03794c66da0cd3ded7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbaba2b34d77d092435ed6957a5f133073da1dbd14a3dd172e221c2167f9752a8080c4378691dbbd3ece57f5346c80c748e87b7779190a62b5999900398e7af0e31f0e4935657818544defc63ee4ac6a504bc9810e71d96c2363b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb80351b2763fe598ea31b97df927a5ed167b47907eb11e8d77952d0e58c5db3702113f6904784eb108a21e5ec31cb7f88c68172f52721d2427c1f398d6b045bd3c5c2a61cbddaf7b2802731b5c3c0c45518512ce30681dc10896ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a50a6b3560f79da89ae74f9fd00219c10055736752963fd6b54ae586d2a6433536729c4138d861051e079738ec8e8b467d0adfc56ab0f81610f6a2caa4212de91089ef1cd33b9e25431a3d266ca380629bc686e12073726c62b08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10af13e22f83b8302f2a1b9f6d7baa1945a074c681815b0b67de9a2950af0b7d957aaa99ff76442abd633f10c38bdc8b36be6a1d697b6cdeba59e61e2a46a8865399d091957f0137ccf8b736705ba00c9426d06eeb91bf92cade20c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h308bd6d27d26ab8b749b7a534b435b97fcc66305f4da5f0cd15730ffefccddc9965311332342d296ecba354fda91ef23f321db9626e43baeb24e8890148110b489c561cc88d43aa81aa84e7b6e6729ec97d859c519b9dcff1f1446;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d4e6925a44a079330de068e2ee696fd3c0c8200d4e536d4e0b6edee6e52fe8a91a7d368c8747101ea69eb790c64b47a780b81bd0e99b4265a71d87af51c958d7ef1e5224db56721223a2adb3fc86ae1c4b42ea56deaefd2bc2740;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efc993b9c6ad2851578bbd16ed55f0ff687d0d2c67e6a816dd67b2064a0842249595d4f138628de9efb245b1ba5933bd5f79f2e23910f22c0974d361a3e7cd59fb4e7101e248d01336cbdb3a3b9ab3520d626d93341b22c80f318e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a15c8f79492758cfeff7f2c56fdf7584f62154ad5d6924d62d6281195549afdff34e5b16e03e888ce0d142e79362dd70e21e24a3ac4614e222b5ee67fadf7e1ee476a740945d9fc02776d2fb774c19a29d0c7e818247cade674be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17eacbeaac9952a30a48f73a66cf09165c26fa94d5ff6fa5d4d97b7bca0464abd3aef10731776551b85e0820070cfbd88ac14392c56f607f8d5d6b76693a187ee39afe1db7c8948ac4b1777942727d92a0048a46242a4f709a5fd7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h879f639704d4cbb67db433a70a6d757abf699cb686c0cedf0008bbe42079895180fe4a76cad8a4ef9ef9b9d666ec245f7a67d7f4668bedb48a590798be7be08b3c1a15f25495a5be56ea3f02b1f492564491a7341f841e97e310c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7b78f750d2ef5e2c60ce90368a04941b8e55918cc14c730a11f4f6d1cb47ed47a1a6e6e0ee4a46f07ef562b6a5fe95d6695ea271bedbbb384e19f95e331c1956ad922f5c40c20f63280af784e8b26a32e3915c0a0f9aad1d54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h434d7b5cb9d07bf377a85af66e25e683bce59dd3cacfc5f219e5b6d9d2e377ca44ebac827e3b3cd7f418b9d3141f5ee14feb0a1843815d0f997fe95c57422329eaae320269a8533d8ead280107c14a06da2c4f3a105f44c04e2ec0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da40daeaad7022f1723aba630247b65c1caae644fb9f1897a715fd0e1bb20ea4e16a78294ffe293cce79d6d8ec51052ab3fde2619eb5317979b656a4e15ffe991727ff84ea104164298388dd5ff487350af394ef9e20496ccc7c17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188423a821709532e1fed6a73b79d34b7d8ab69fda68159cda58dde534b0da95484e15effb65b557757666deb072fd63d62948df91378a05b6f8ebf42f0a6eabf75125e571638a1889fa291088b5319264f1151b8bf5470c643dd90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13bd54b7abdaae732f938e98b4b10bfe634302ac90de14c0e968ac1e11155c664b8d1701785b54df7482de99a1fc42a30d33e3a93e39981a5a378370a3ba787a0b08918d2bb865b06228acde9922fd89d0098eeab5c09ac131b7037;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha48b86abdbd425aa89b2ec5494aff5b9f4ef3dbbb04053c34a564dd9edc854221938d57340ec5dbc69a75c0a35f720c5598929370c1311df8c03aaaafc7d8853013f46bc37da75c5486f52c7ebff947388f9fd4bffcd30953fff9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186cbbc75c3c494a11e711e128a3fc2e60452b6f3a2c9dd0be16f725b5ed53a65c7055de91768ee3a0ff65fd6822b6bc64e9ea7a75a4954a697734f619d57eae3851dd69a1a558e5a9df1978a0fc19b5b9af7d3f474e959f13e8b41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h959223b9391db86a49f82dedcdc412b80f02778626afc831cbcb9611442bd77e28b0093efe3f2d800422fb4d35560e0a04e29320e87c8bbd9248fc9fcf95fec495dc0375f952984bc39369d5204ebb517c341abd716dc8108afa25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h965339ecef9849266072af0e131a84e2a554aa8000ca43f1fd3bc93829b8565eb68cf2486f53293544dc800fcb338391ab66a9b33ae67a055d01471496cdccecb2ba1ddd0b4e46770483c8134ac8d1c0a6c82dcc66a7172b68bc83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6b3f90630f9cd28fc4754a86b8bd1ba709f83de27393150c85128b287b5e2f55280d15cef06e14d37f0e04e7f9f233be1b8a34ea53ecfc955546292da0213f610b6e23a5e6387d793f1451f563d4bf1ee5b1e9f315ef1fa0f188f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1362713989a12f4915e47a84438c06853041fb87a6a62973af89b3bbf0cc7958b4b116d67fdc6a50f05a9a10ba49be18691be66fa6c744e6449bc44b876b7e3671f8c63a754b827a4fb7d06593df845b75f774793a5798f1037a8df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136532598239ff5ec113be809ee23c918dfcfd285df2614f63c8b7abaa99f02781fe63cec98235a15549e5ec7b2aa16103a67b801911142941f02e94dc3d8d8b2d5c07b40284227b2ed617776422f230305d4bfa7ff6ae1ae597b57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1fba94199ed76afd11f7cde8e96b02ccc664680718fa0de5ad37c3526552ee8d5f14e65385c5669fa80c3bd903515557a00c64312dbbd704a9b588c02232fd58c7f8d8d1d5b7a93c5ab9428ea7de08999a04e569083558612a11e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3a57eafdf258162ef0214cd2927d11b4efd1871c3fdf94ce20843ef148c78ad8e3afac13362ee39dc4d1bfbf5f7b286f060dbbce83a75588b937cb720c878ee5d67b1d164e9cfa08dbc8afe71a7852b4c795f108d1a8d31673b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8590728fdec2c969630e5cc7bfd233e4154155560d83784811851fc73fb980709a2e45c53dc73724b4f70acfe3f5d7fa46ece59c6bd38f5aa193762367729df128ce77fd787c288b196eb9c6bea8dbf3b263595d29ce137b29503;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h492a09bd22deb53a34956e18790b97a20ba7388ba9d8b34c001cb85477e9199e784185a8254a7e80740480c6c267af10c44ac2dd910c7f7a7eba69765eac0cd12f5eb44ed3d632e0be296b6a509f449d09880cc04babd81b20b541;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bac834a4825ffe7e1e40d076e18a4a8086106a23278f36e39125b2449edf89d57f3df08571a81f2d653646fca7401079cf21593406ee84c9996e710837c006bf0462fa7e1427567f9cb9985dd2960d62fe8cc430ede2aed6daf4e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heaf64e1716c29aa1bbff18458ec360a7b374304e3d68989678c61fdecfc5614ba9d35ec1143258660e71b855347291b9cd4d05fabce973cc801cfc2f3ef4e2441826849cbafe44bfefa77f7ec9e84964e3a63ee7e2601df5c48cc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bb016a071900dc60b32f0cb9b7da21939b7f889709a9351f770248d4880a5227b624da6249351fb7a1db5b9438fd16ab1854578eafed02ed37fa1b77700473de70c17c0385833551381c3c439ec78ad506fdddb4d75d370a69dd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h664738a0a10c2a17c2e6f1fdcb95bf3ab32da9ac2f85bb03be8206d7ea6f63c46e2f81e505f2f6f02ea1db8461fc15f1d20a38dca5b61f348e5ab4b627ef477fe8687bc40e4d3250c537cf2a400be49b9430a2a4311e4290eb4dcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd05f99612bf3259c1c096b8bb8647d44264b536cb62ec3397a402baf2172b26b728ca49fbdbe44041520244f49644363e83903bfae26005880d1931249a43f3a75a04cb005e0b7765a479f13392203e48d7be400bddf34dae73ae2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12406c0cb598df747de69f5f5a11931f33b4402e4473178181e5940defaf93247b853b23cd03bc7de2b975cf0777ae533963ba46ed737dcba024986d3e7971c1f40a6f134792657d929ffc86f472e36a575279950feeb050851cfbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c0891ed3b394948aad1b8891289704f96f50d65e9e56f82220ea11dcac6269a5a8116141f1869f7d89b2583ce7172644185126d5762ec37541e8bf2c9e1baf3cea8685b3f632b9b92ebbc1b7d5dd0b63d27549da3ceda6d867c46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h288ad8afdc78a06f725abdc610156a433f7f762efd6bed01fe5d27e2db4324dcf706a8b9ea2b1a74b760b16b7fe2c1a7d48a8d24edc94b0bf11913ba5da87a04dbdb494be28e64f659b7b1b839822e965288afb8704001ad89ca31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h237326e0056f39ac8f305c2a414802e33d7d101392826c6e60cc27bd678847e12dad0fb847e69d9b303ae2ffbc979e6480520d599d3953ffb9dde32f74b998f018ce4ff4fc41133b50331eb4b5a2f2252b0cc2fa5fce047f6abf14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8512ec9755732f128414341d7135221568cb6d865229c092d36063ade3fbc8593924341fe968e3ba81f9a34272e4ce03155c490d63ef445a4fbf4fba5ef2f6148f4597757435c982fac86f13cc98ab58e9707d67d56f68c75a3952;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he005b988f3eb440db77aa920a7c732917d7470de2dc116588c42b03f8d52dc8d4c6fd7ba3b80d4519ac3062e01835f6ddf2bcb317c4b8fa54ab8f126826015ebc0b0862d23c3e09f78b6318c9a73855b6df10f46ec4056ce1e5fa7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce6ee94b3c9820ce674401c5043f41b33874b27c24c956c75a501c52410b4c714974de163bd7c81c9274f09c6de240ab00fd7772c7f90892bdaec906b22f3da58774fdb8c227dae61628df32eba901f1950c60a57ab129d57f35df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11dcb937ed95c0b0deb89578a08179136367cb0aa28db9b6ff059a3cc727a1a3b981dda539f12916fd9c107463a845cb446d7d04fe5cc7c3b73f32c7c4a9b0eb5da06b89e44edeb892fa77ae2b398081b9c41e6049dc3fdba2475bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a3c877839ec7ff92312b474d3f18eef8cc79c39a10489ebbd701be4cf13739093288fc9fab73a86949fe91dc5acb49f48e1a77165a0ab0f7714652b145183f7aec0aa5d954c0276584328c47c41f88f4ad7e3220887fdd2f0b95f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106d9100ef3e391604a39397fbac272f6feb40caf8ee86f089aa4d5f304c237a63c711296030ca2e4e53425543caebc56ddbfd65d2f863f44ee09f531b2346853c7fce2df3d4a18df218193bccc8dfde3f7073828b1ef0f1d4fa4e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc853a0ad726bf7522896691428bd7a78b43419642e6d2690d5d7b2342e2d4260af20486c490ca81df1eab851b1993425343349c54a1a2deb7739e9a01a02c2a3196e3990b797824b731e2efb7a582acca996cb0863277ab255cebb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb932d1049320598b92dbd99d05baa7dea27f18bfa9c9d8468123978ff2934da7d948a67524a4372c75c9a9a61ee40c7005b5b9fcb932abe88aa4ab07c0c24393b979c50c539362c2dde8832bbbefdfd7aba46d044dcc01a9f024a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164a4a932f1cd58ff5ecaff61824dc0821579df4b034768051dce4226602d6f86e089362fbd0f8cba425e9bd6bf90698bc461b6b55425f7d578d772717b8a931ab1922e28ecd4cac2fff407b4792d5d4dfa8e3238e84d8ac9b1980d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7226429cccd2c3cc12d624c1f5496440bceac3945761e677336245df8044438d4a7b864cd32a4d5665b025bff338fec9919c48243bd384cbc41e9c828acdfd13d64496e09c2b0c70677cc702a43f13697691ad3de5ed3a857aa9e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7d065b440df00e883268c172eed63d3e3f44086c91fa722ac08d870b5fcccd6fde6cc03f436f1f226624b663c533e2076cf8a20c932cd6c3060e4abe4669c2ba727f04b1a65e24e6959b6eb3fc6bf2cfa3597a1fbab33586cf47d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b10fe64a0d6da3c6052766f7448f3a10611e3276344f62be7d4b5ed6263ccd5fbd5c3c1c22e654c8ec1b46d78fe234aa021a5b9e1d4776c21533ef457388e7ff5e961f6acc3fe745abd813e131871ab84602623a1f29825c99a1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'head895c078274fa877ae7f3c08530de506eedee0394858061b4e8e8746ff430967e6e79ea440d5836b515fea133f334189a9737b5663b52459cda8b238c6f7ee4b4dbbae1e4c15e70bc58762bd5f109a40deb7a928aa95a2711af8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c8b9f4d17002f174eabe21385e3dc35d5bc73ec67855c1d2c8f8d283328a6f29fdbaaf9b09ee5183f00f80ba3815b188e47160860a7c71ef55d21e403ecb3092b4e92553beb0c4b18914744663597bfaca19bbbe0e5c38a8250b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189c175b25dd8d164b3783b0539534826a287ea38479118b349d9e2d9740ab3e6550d54835765bf4bbe32ec0abf81a4f738d3e02a416a070a3df858743e06621e4f7fc4b0c1d0f0ca92fbd21227107fad6d89338de6c8e39b97142d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f1c4be6a0c9c0e15a5756fb2db207eea22e925ec62cd67532271d011dc93e71ff8ffc35c959995ab0a46af2c78c7594ac4ff8ad60e0ca053fa7b8789446f50d4a584c57b4388c6ed190068273207b1efbdc29214900b57d11bac8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf515b2544c9a0098f576a708f1e0f0c54c5d20b56be1003f924b5dd800b85cf55698a4dc87daaf2078c49bac507c4e8a2ff976ce7954f8b22d4b1f7054dd1bc847ef5ebe31bd76900320e1a1a49eb513fc01738834f8e27d9bbb64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106f22c58215692849e9378f7460e32e6cfc96441db0a14f7b19ea344f38dd108cb61b04bc910aa125c8ad8684b44755798027b3038388cb4b005f72abb8b7acfc1adfc7a9e0849978a7547e31021b86dfe7651d112ef9c5feac95e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104adac2efe49cb548c3bef84da78352c03a8aa811f9e6a3a7aac033202009cf7d7e44eff94612d6c8549be78ee66b70d6ccb25b2519028916555fc42fff897d47042f57c5bc77d24d757fa5315b7781666ddc0ab9c750935f3a626;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2740f49549af7fa62fef2177f0f87175b1fedec6748f8682fd926faf293c881038151c98b55631bbd4719d77cd86072cc4933df763cef403425cabd566f61fa65437d153de47198d43b52f9e4107b0510b54af400d3ac6d87ab282;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb26d3c51eb8c39405d03d6ccec5388cc809e4ad14db5024580ede1a2f849708806e54717fb8eb06549b7714d142acb05a287d8216a269699e5e475d0816e596a8643f9a09f21b058bd6e8051e08d08a7e70e3fc5f0465b99e904e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc51d6f6279cec3bcb7b5ff90052c313ff0aa221f45265aeb641436eb2c630d364c7e176c3c41fe0c74861e678971d6d0e9238b15daca9caa7b653526ae664ae4a7dba0cc0127c956ee3804d7dd2959c0c51f5fe71e06b8bbe620eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5d0d9f9aeee3c936a53b0b750027051d4ba97a6f17434b60ef8882bf594a370be6f8ca365b33db6ed11736e8f8bbcc9b1b6181e8a98812781c709acc5966a3d4273e2549750152152c342e7cd947e60c35aaf1a4035c314cfa073;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb38cf35d39a889bcaaa08fd9d01e69ae4dd2b9303c5bf42792f44dd6cb54d45d575acd8b0bea1fb88f4f27dc4b8f5ee2d8d2730c5d6e47a637bb47457808c0743c36e359cadd96c885d266d248615417b65e4a8bbb7302ff239d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16947b29dc34e4a583b628d5c100d224cd50c63d55bf24ed2ff2496cbdeaf4715990190556de832b5b37a05fc73864918b6f6a1fa00139f3e0b1ddcab8a5b3528fb8861057a1008b943844afbaa169dd97e993761309399b11d0e03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h340b1c6b2b0e21cb8bb27282326a3afd74a3a607b36c7c8ae3091e1d5200396bf2ffb7ad659d2db863c70e80d7c86ab84fa534368e0058f29c2d451f704770460013d35d0560a1771e78102da42f4aae67cd7995887f618f1d7dde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc58c553af67aafacff860338114278c6824e46552debe49c5c3bb5a95f441a5a85649de90d3ffa5a7f6790fefd788379c02b48af51e4e0ecc7c0ac84521d819f2fde2dd81fcd1ae26bcc68a6eec5cbd8fe0ed8f09a4d32b2b14b7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf901c12121cf91702419709ee7f44fa65d05b6ad5ce95a3f2c6527596c2875b71f7168f7c413a3b86672e651b9a13065ab20167edb0b798ef92d176dde37dd662d013e084b8a0279156fb4fa6ae3560306fa08406570253d859607;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13984c51dc46375cb2c84f310f85c5a0057c315c273f983e325b668bd6f56dca6dfdd1d212cd7f51e5d4fd8646d659f375cda9e5b233cb72d8c782ea6e6e37985935d4772d8feccfd47f6c337818769c99480377b0230ed192024da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ebb62dcfb585b3d6ab6086f37d07a27dbf7bd0bdaf2fb52e8e0efd2540d30a1d612ffb3ed539439eaf5d34d4c5f8ae9c1a217d429fd8c1bd0dcc5b76a891a4c23161bd9d943b84302ce5d0a9cdfeb60b28f9d7cd042969e024770;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f69cfd5f3d9cfdcae9279c39eafbb712bc60ebcc527c3c85b4f694a33dddf39857d9d2bcd7d4113bb676e4fe521fb3698a8304265d57e0ab51384b27defab5a805359ac4d36fc5f2ae41f71c4555293c2731b38fcd9164ff84bfa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he10514ccc2003755aab233ac203f51582c5acd384ba1afda42dd203310362e436213c988035c718ae8b9eb98d82a7693c71834d96dc124da9c3236a8ed746c94636b36fdd3e55c71f06030b578f178ca941dbf11dcb4cbd6aa7364;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5752eebcbcdc9b6cd5549db57ca4e74f0e555d9535f67396d2565fd2b507e85f63795ae4679bfa94a562b89ab75c15fcd835bfd4a395c3302e0fa86bf3223cb74387b89f76b5ea95d484fadc8079e2e05c312a882c2448118ad373;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1c483bd179d3039bdb0a0aa1da581e3ee866dc55dd97ed56cb3cf8c7de59f66db9e62f46db579cea7a3beda5db46658b231614dbbd78f092296f27c4b34306b62349820fb2757c7a06a4e1e5e93e58d4f6df0aaa31a16e146724e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1ffbd3ee827a883e29057cb61e5a8751675257053fd7e621ce05ba2a2753c0f91f376a05ddb0925c77850fec942592d52fce887196b50843243178a6818a6f8f1efef0b33c4bb3b044f59139b256f11f32a42dda40e478bf03a19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5603815bbdba80a7314a7e7bd0edfa4edfbf039d785e4c49052260c7e900eeb7ab5d9caf38dc3835092fa7b1bf72cc02755ff8c0e6b7403a4ba520398a2b7146b94b7c989844517ccd8b6435b96c0f2815cbe0c8495d6984cfe26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad230cdead00790ea73b4d95d0e61a46989bf0e1fb123051b2f10248454d13fb5c7dc9faf16639e2d9488e57470e7c92ebf9834e105a9e5c22dc52297c48380c4ef822370d1245f03a29580ab4164ab5327eebabf02a8d04909c37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c767ea53cc401ac087accd47282aab7a5abe334f23d15ff0d59a975d292525b951ccd8b821c1de1f2991ff6fc7baf2546411b017ab43b564e61d60d4cd2d2bb2d7bc680d8d974549fc1f88e5b96f14925d0c1ae8a71e68eb07eb53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98b1906901d68209dfa838eb2dfb6d4c2bc880ee59d816f83e5d61f7b49b11b1ad144601e8c3719fd9f9b7bd0e754bafa16078ee4151bb5795ed7d3af261ce66e895d555f31d5fe0fc07b0ba2182d130172d5b19f7c547fde68c45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2aa5831219ab3ad04ab85a3cbb41e2b0827fd2dc7aeeaf6ebc4066283446458990e8c3cbf9dce2b6253f5d196aeb0e689f9b9760fb8e76d96a79c69512065232e689de5940b68c59f7ef1cd8aba91f062a3ac06184ffdbcd71e8f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b03067bb1b1c474f2ef381036c64442ebd4ad62369a3f1d7bfbdeb231be964165b2519b541c6a65aa997e1a3941db1b2cc1bb55b10dcc3624c97edb93519cad787dd3f94e8d0c5af6865d3c1021360431d98be700368c1b61ec71c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4052e2956eb6bef46d2e5b31628529fb0a5d97692c3139f9d8ab340c8217170d7add8d11259b38f898cc33d8af9315527ba28e93a94eb7703ca3486db3acfde7fcc147964f519fd5209e8d04e3982745a820e421af4c67163bc331;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11277bdbc52a46a784d2d97a494b0e1cb6c63c9d8256798a67114d8b1a368dc8b3c10267840b9ff9b707215e75f905b279a11cb2d2469edf7679a3eec63ef999a0f2f1873b6cb892aaee8843ca83c760d681e83a0f0539666a30bbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h124e5d2028eed7af0110f8073776867011b455802458cb45bc30e05ab4134edf5f60568649c02b0bfa5197c0ee41cb1cdd500b4384af1a6a563340e2f2f599b1e1e2d147c8562c0bd828b540caf41e70925922072d3508bfd85fa41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc1ee294bc03d244bd2ee9954b6723d95f6ee3fb545305fd4ac6d65e41571dff4f4a2ea1e95afb41fe3f82989cb7cd9548ca4302327d858d0e70cb03e7d608d6977e01489d30492fbbe654ed0d8dbaca0f8c79cf6898afd781922a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64f5b8ede954795fa44cb225c0266a0632591314b0c0423954efd80aeb17d1580e0cb15c3471e51330399fccf49711b6763b616c4c5da81ef9146c708b999134d6415f7331ce7a7158c3df10a8bee9d9e32ed9ac3b922310be25d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e4efdd74032365a50d9c4ba141993a3dbeca83ff2ef43990086451d885edd23f9f5acf5f879913310d772949e4541859bd7d6e08350f997dec20ba24457b0884735f0a6ec8b7dd28ca4aa866b2a71c4472fd228afc87510747db3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d943181ada2e4cd813ec65c97ae8298c75b71db7da059d6dfaf3e6ac431897c0c3cda4e97bde8d1266441600e9e43fd0bc1366a75405c5bee3e94359035c69d916263d0b93546008e66c561dad2e6f3e0c627e2dc7a266974bd56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he220189e97060e58466dcf706a10671d8b8228b420367d64335965e39241f9ffdc3950307c3d00026b8f6c759ca096568e327b1662740bdb0f7ef1c5ff6d1e66758b92ce0e387e3a4f6f80f1722e5458cc759cba728a6cf75c114d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e4e78851e4e910999e3866f07f9ad99a6e0873661d11dd413f0f86b58f2ca44aafc5ad5c3e913bc0d66ab9e3faade4ae4ed4a225226f25afacd276228c508ea929a3b7d5811b3154f371097f23317dfbb6046bbe4edec4255097c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34a978b733b986e94b4439b31c477295aed55cf011e563e10c05a012c9390033fd5d4ddd8420e7ae0e4a5c216233e416505b76f7f3c9cf36b6586bf4719bb38160b73ba0b88cfba8b4a080bd4dcfc5e02282af43935a736bffe8bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39c05adf6edcb1b204952de9b416eebfb62e6c01f7fcf207218d3659a8a041a65abf5837972bee565ba4713534eb9ec27314f21bd255d5701a0060756c6f9e062392598390101d96062a2e5b52ef5806f0eaf9c7604073c746a33a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba7f78c702f9e643773e7f60a8bc683ab8b440627d2c5e89ad26d9cdab9ed829e02bc9617e548152b87da196a1f2df87680cf7ee6352be71f070e3bf75f5dc733effd15c70fcb1f8096395561149da8fbd4515b4c780adaf38c87c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91df59b3dd0167fe011900346cf60c13bfac2d448fafec53ce1764d7f3b16c070a355108f8d4e9633f4bb0c6cabbe993922e8aa389429a940380b46a8acf8fd2d447a8b2737da1726ce1dae92b8c0136c58fd8b722319c8c70fb39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5544bb32150401ea4944a600d0de264159d1881b23446ed7b701ed61cc523747b2dc94ed3af3a6e719565e9e918fb70f4b732f5421f1ebdf184926c694bdbb51ed098c1a79be5430ba0cdc6e71f7348d355cb08a1e23ff4e17f87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e0a6381b7061419b9d05590f0fb32478bbaf003145c62e5bdf07cda1e413d059281398d4f8373c4a6b47097698b22bc120ed0df006091b085fd0610643511418abdd0097e48b224a952d6a46a874b5dccfe5ecc3368dc14112f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a2b1a8f72f64e51bb3a7fb606dee9229b19c532d95cc96da3cdf2717135b7f65d4266279da2144955d9a666618fae07f569fb10b7915794235e4c58feaf04774e0523f24526975a625a787401adba99fcfbe8fdbabd669e1d136b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93819433038dec0ee78f8f71df6921e5578e37b0bc59556ea65b06c0abd4efdbed3cbd9f2dc04b1e8e800f3d355e472247f49481ccf47fb23b487c9ff032dd1d4ed33d8c55fbebe4dad5952c0ab829a6e704c69ada063b8d8dfcf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c0a4eb657e9c3e4a46549ed5ff95b16feb6dc89f7f682532d489706805577be3a424015fc82ced80cd60b7b59bff39e6f01273ff05f788968aebf2a95f80c36c9d77d40fcdd2c48a921954ad54c2fc85de5fcae96b753ab9fe271;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e9e435c807d1ee69082f61ff21b6525fd413dd8934242c882e2e7e0b441c5b4002f6f92ee56d3d62c8a7185e24d4e28b2e0daf2ab982957e3112aef6ed8c9c1279567a4cccddcd0763517f36134290a7b8f63268c830af4b9287c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcf0f9917d34b75b186c1f5b8d7198913e62790e347f0376658773328c3e2c92c5356077613b874ca1e6829d64be7dc7334baf8d6b3abbdc63b615e1dd30c9babad384b9137a07825ddd63f112b6986a50d1efb5743c388e3b90a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h653cb9f1a320dc40ae21abd9d7d805fe6d8ca840968faaf29dd89c463f771bc10561ceda1b448febf1cb772f3e076d31207e3f833ab4d1e85117ccaaf15efab385166f83040a19a74ee1be763d54a9b291749d4404ee5c7cbf5e2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1375206854ce9114275e6d1abb9dfd130124b3c2b17082b1b3693c719be377da3893a68eaf23eba464f87e3e7ffbf8ff68faa66ee98c993ec6640e6493493b340e1cc630ced0e1abf9c36464a3d0a54aab5af4dfe886fcb40986389;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6eb78694b0ed24bbb65f4823b050ca28e8af5505b2c8a3e0a3d2846bf8dd2c216a2f78b7bc23e948932ace29cdb25a7833e516d5777ea8fd0c13f1e8afa5a67b31fafa1d936825193a4de28e20ce29da734a58b6ae516aa226071c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2675280facb185795573bbd4ee648bbf8bdd7ee4f9c5e255663ab402ec80d46bbf6ff8cc92fe525070eabfefb6341b7ec75bb8c759b81674f76a9581b70d0100bbd81ccb769afdc68a0ab1a2aeecd4cf90367da6a6c90b9849e4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5cc76ad1bc3e1dd789ba2c501348ed7792829ae6b93a50215f16e88904e27c174293abdef762976336449c52121ef25556a3a86f275dabd202991969955e6af4d94896e0618bd76fc9caea07da6e9923265099855a7f7de143346d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1902befbb726703e60151edd49398a93158cee7f1519da8cef36e0465f9ccde2f0653930d94819ea531fb41f8fb6720a9a77d0e5ae77383c03aca0f941e79f1a3c2eefd2025836f842879ea285877dae876ea555bda6d83be041044;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31fd37319a01c95851ff6ffeb8e5e650bb14ae564664e19f7c54bc3009464c728db0f962d3d1ed5460d21b80e96717d77283e059d419050d3153282af114a0a3c723d22735bdc6cd2314d6f45c7609478febb6d89b2b13fbccfac3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf94b443e73d35817ccefbdb17f27b982347ca172dfb318e07d5601409243f44aa7f126a75898acfa945087c5c22519c5edf7758676e541745986374c8120243d45cc64822df5a52ec353fbb899336ba179df93302fa2b965d34ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf63178d52b279ff2dded30da12e24d5b3e1eb27eaadc1c9d2ff444088f7c666382ac3b0cd4e9e572b7303f4a6bc0c9d5ef34e3f37c1439f6d8b65d296f27348645067c4c6d61ccae8acb17b4a5b79300cfcc6895cad25d5b5298f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fd2de58e86dd3ebd85fffaba9560dbf2c5c1a82f9eb847bd5afa282e24bbbf8f11ebfea791fbad892bee2b4df69cd3bfaed3dc7e28de99860b779adfe237c4d43c07e66942c04422fcf3a8802cffd747170faca9fc4911c6f9acb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3cbf2b763c90475329c37d621e717bb7b54af4c2ce17b065917e6e74209ea187f64de7c765897762fc66661323da6c4a37cd5faad91dc1b003b95db18cbd99fcf268f82065155129d98660f292b44c54a62edcbc57b5e6d6060315;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180740c46f92786bd16d3d1ec73c63bb3854582e72e4921ca4296fc9dbd433184dec7d73462553217a255b9c611bd66521437b8ac3f8594a5cb933055710d93115137dda224a2e6b3c7bc334469a6e5ccd92847c057bd93b39bdfde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c9ff0c7b92b876fe29824d459e6adf85eba45421e42bbac89b49ebbdb046b487255d9394fb729cec12e02bf829e404bd61180804b1106d16dd1c88ffe4436e3aa64b95fee825ecb579f6793fe9c02c89d2536cf54ab736650ab93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa1ba18fd0cf011bd526e11153cdfa976b7c5bd7d5f2ed8b49e82cba7d8e6e1365553652dcf26ce8b2ceb5e17d509f224c2b74d629950f30c4fd5ee41a4214496f0b7d01c511cbce4f3737ada154fe2c958abd518e64b6759ab075;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h654fd583ec95c232c7ed0e06004cffec9c1cee266fbb36a13c907d030cb7cb5739e945dccbcba216cfbe2c9554ca7e6bb9e9c6edf9a5aa2add385594a5e6d04b14fb5113a2d4bea41d498e190f8f4d831f9d82eceb46e0691d90c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b9bc79bb54180bfe71de893f2b67109c57582d9d4f8ec0f0cd41d3e11fceab0a1bffaffc36ee77fa2a9ee6dd81ac9816a7c734681c8cef82ff501b129498d1709a0e9281c51418fcea79a29d5596809babff5e8be2ca9aa2e5958;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90ab7ef8f91fdbaa724924adff876c4806528cf652fff82e6b1e469bccd98e6ea4a1910c3bcf72e2b3b68c641af31f8007a1107f78f75f3fa5c7fcf32696a4fe058226a0d2ba1f467a34cc030181c9cbce28869f2cdf6ce2362dae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0cebfa6780342bd4b66c28bd8c52573c3d7b7b32eecdcd9cb19f481f6da4e7f067201986b1313bcd84a44b4e830042456b6a05fcefe8ff75ebb716b946497882d7b3022f1fe462770b68043f7402f9880012f4638df187558be70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a007a76c7031682a46d5d9c30fccd1a9868cc35e5b57ac5068f12a65f474a3ac0d3c0d518324ae8cc09b5fb26d4977bcc3fed76a6bfbe2539b35e0fa27d61fc6ee65be975500c13889291f79ff65d1f6c68762b2ba8f339f55675;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19db0d6bdd358fea7df9f0ff4926f6c85d11ece52d0fde6bc3aea5a42fa401bdee0431d3666fa30f2504c2a5b1fdfb76df7260d04f7e681378e6a07ab254c143aa38d0f1b680f57ae501062817e2879be18ff04ec2d3461810065be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha60da0f2c4535e20287c50b25f913f16eca42a36f9266ba2adfedc04e94657e9cfbb4e16909b6a9c0cd5f971a8bfd4563d1619fed103cfdea255250b5ecd6fd5621a414242e44027c925fa8a38a70548e7fbff34f57cbfd5be3a11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2e4abc4eb65735a01dd0274979377be318e7fdb2ce5461d071a30ffbdc40d5a85d66d9865e150e3a2dfa86b2dd499e1e867d293e660219d0b69807ee698da87d3eee0651f8e5a9f5fe4b881b8db1d51285b238a4e7997ecbef5d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10079e691cd68672fccde9240f38fdb6876d337529b9073df9c474f7e53fe823aed3e95461954cc6f300b37a6a8e1322a5feba9b8134721361f3a7ea26143b0d2316b51a9d8af9c044fb3fa9bf894d3195315d5c7d429a5ca931096;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfaaa8e91e1f0782736bfc36efa0ef33a62cc4db1fc67502bab48ac0841eed62d719f88240653fe57518e99fb83dcf7db508db82fd1ce4cff210a4121776e2c793f870c957646a248803cf36654c7871be0700f04741868f3226994;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4d25abe8dfc74607dd58273edf0993b701c289127ab32817b30cf370b5f263cb0877ee1b6960b7356478b33028ad95c83b5e3ef3e45230686727a9c0314db70c9f56524e82c41b77d4c744e7b0ca74c184b54a27c12ae7e112c55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d47a5b5d81cfa527f3062000f1560d68e2f6e5ce1de9cedb7f06b8dfda0eb257db2bf60dac7e2a6adfa591038061dd783d13d2d98ca46e3589bdd7ee860df6d21fd2079b73f5233480666bff35f7c04b77c3eeea58e4ddd1272e05;
        #1
        $finish();
    end
endmodule
