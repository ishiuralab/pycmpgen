module testbench();
    reg [20:0] src0;
    reg [20:0] src1;
    reg [20:0] src2;
    reg [20:0] src3;
    reg [20:0] src4;
    reg [20:0] src5;
    reg [20:0] src6;
    reg [20:0] src7;
    reg [20:0] src8;
    reg [20:0] src9;
    reg [20:0] src10;
    reg [20:0] src11;
    reg [20:0] src12;
    reg [20:0] src13;
    reg [20:0] src14;
    reg [20:0] src15;
    reg [20:0] src16;
    reg [20:0] src17;
    reg [20:0] src18;
    reg [20:0] src19;
    reg [20:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d59cac4bf6b1c47b1809f49334f1cd9fdc8403ebbb68801a6ba8a29af030800782d84debd4d94bad254513f836af6ea9361d1fb608aeef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c21866d91a960f7e5a8214464c346237107a62cf4cc4dea2b52d235b7430f6b412b3673283253fe5fc3108d5b0d5c4be1860f04533c0e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h573ba33b399e91d75c285ee721a7d103c8808e9a4dab0a8508b43b6ad2a6be37a213c7fb2b18b09916a540b4936027e0b4aa1018ae452b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86f0d8642736b0e04e67794c0801ad2e98bbef04ca0bd6f88ab97262102d951de89a2df95329124a2e7768f602ec53fe0c8a8f31af9fca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177f89e819c8b11fa0ff8395dfe27fa90191b78607fb62b0c9892c09555cb0e020aea8848b30d313b4737aa86e742a5d2a101ed06506a74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5b7288e9bc7d514aad546083404e284e907ab382b773d5dcfd59e52752541064adf83ead0ac1fb22223b85e32f8bea1e3a2efc49c5df8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159683083dbf1a5cec0192cc6dacf6de4a49717085591bbc3a003ca21680b43dd7f3ff12547d0124f95d21119a301ec5d772c5f95130553;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bc73fe9d5b4dc284a4a2fb80485887102fc54c4a5d429bdd7badd526f2e0fbc7e5e6823c4fc7fa438d7bda17c6efd3a2e66e1e2835b9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h363973fdef47a6379cfbb0c8e37d2e1971adee2a68290f432cb3b67f13111495c9736fb391223fadbe62d6ac8b90f13c98631a9d73016c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92b2e5965c8b1eded690663f5a52890dc224ae8643b9b713a8af9c67ebe81f6d4cf8a488d6c6646c7419404748d57dccc803914205d72a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb75b3a937a939c5c41891f3326a81bca2f223dd1f6cbae78bf82cc448fb71d593c6bed665e3757424e148f1522179103f0dafa6d4e8978;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ad4aaaed3b9e6f3db33b3204c683ec85e3f62597bad23bacd1958ed88d851ff0ce7fa56273d8e363ee35082ab03488ee1dd55a4c9a84b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124df5c4a1d3f039fb34a3820b93ca975c612fcb8db80b58f6768b35d7bfad4a2d5b812e6e8e94eb06c746d2d7c17727b8049e9637cf355;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12aa5cef4767c47d5fb1e67b88df7feddc1a71e74a09926025ef4b917738957c98f7234efaa58b217d414232fd2d9f2421a15b35e5900d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h639acaf51d3d90ab5140c782d7c0ad185de034eefae7e5157cf2fc09c92d6a1971b1c006eea12bed4e07a290e4cc9c3eb7d600e1d94b8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118a2aab139ea0701ebc463e7f3152f2e42d605e18e5e261c2194d2f636baff219ddb25c5f75b4e3aba2ad0d698542dafb3fc1cde2e3441;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122c1d25a3946a1db7aaabf459e56a3f8a442d1378841673159bc98bac383955e6117c218938fcd15055a3294595d25300458b2a3d62314;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3baae1516b8b7eabfa78439465ff54e59857dbfee512fe026c742e6d2cf9becd35be3c3d7a58cce6f3f265dc6128fb5cfa688f5a59aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1a0358d5ab6d3d117e3a22dceab8b1a3ef17b7c357929bb940c24241b73ab55e3877ce273e79bd52560ff798b78e67bdc73e9d75b3e59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b89e8cf08b3ed3d1ddb1c0d228769712464d3209cef835b7cc33a1bd99135bea392e22fddc9add23e4fd7af393d199151d9fb01f3e839e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ead2308328026f7bce518955077b0d1f5fc855cc0ddb5c2d01678a9ee38f2717a8969e3ef7f9ca1ee139ce0a53197c1f300be10494ce9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd6471ba90010b43df6c463dfde44ba9526e1ac93d1f4f079d205d281212c1bea849b2288b364ef224434029b9b0a3c9733de534ff060d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f821291863b7364b26933b7c3d8a01ab57d9bd9d2969ada610a3b9de5a93bb97d06adda60210299eb44a83c1ba6c6c90564ed662f0c14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80d8a82d7f0f39715e19fac501c93dbc3cb5a1ce18eedde650d0ffb3b50824f6adfd4c010d6e68f55fe91981969c760eda4f65a09615c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e6f98ef693d3b3b66aae6c6219a3082ca6b0229a82476fb79a9e8ca98f31146d3ba94ce1362cc34d1f744c91adb1afa42cee852ead9ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5164ea82163ae4afd470ab949814e76ad1eb0d516a22b6c91b0a78dbe5d91fd7712acce3ec9b1318db22496d39da9db943acc4833d42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198476efb6de140e2360e7b4995a2e56897c82afad499670f9925a22839f7ec933f45c0444b679051a579f8df235d77dfcdab0bb77ad838;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188dcf682abb8a7c8aaf6478db197a5420bc4dc7d58278399b476c18c7829f8d981f1870adfde7fb08e08b454850ca33e195eec68e6af00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a172cbfc19a58dcda75d884ccd2be7494f0703cc31c1096ac51a3340d12fa54c3da9a4de8e5c650fdfdbb9df7a06366d7cba9839f3c82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fde8c45c963b856a51febfc10e8a6beff14f40b1a0723bf139ab905321d23c4656180f826c40588fa73ce5ae0504c709ce20ce39e8c91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f3dbd4d080cd1cfb0da6c0b1835b4219469a6f3978db486c8360ae55e99ef3999303e80eb5841a90a66d080eed9fe6aef53355b949cb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1117bb1845ebb713419ac2ecc8e584ff2b6203ecd52b7a890766e1d99c10f6d95f6acfb43e309fb0abbd6f6b707c5647fabaf23980d63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35adcb7dbf773764eeaa759570193e2ea4b803f951a1c28f0cea8d189e6120e9d6d2a0e26f86d79acbd4f51e62b71f3c7fb4abc7be2915;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117d0b0f41d066d7a1a0bab3a3e85ca16dfb7cd6a16d441f33897a833897dd63fd1785c4fc97ed012f7a282bfa4fb4bbe9a5747eca1b94c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e575df2a31b290ae3ddc738ab7b9e55c2d8fc3f5d6eadd99b66a4bf560fcc308cb8d0f63b52f67cb93b946bcf233b77137761a12b4e29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3078e2c7e547506d97ad06f18bd4b35a23ec0b684180cba70bfd88bb96a90276588f9eda8efc0b64ac9a83475cd5d368a1fc27a9e020e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6febd86f80ab4df14c0cbad1e509c4939461666ce0a11fed9f11ea4e7f7242d250e8d7f5c79a598cb6b4cc80db8672fcc6ee5113075dcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc550dbe6f9df5d278e547bf51fa3bfcfdf21c5d80c4f04e3902c3c49d6f926d16ffb2bd52fe10a2b4dd5573d35ae1705626882a9e18c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b29cfc596a5997b1143bdbb2b030de7f78ed1648664559ca201871b91e5dcb23ef745c8d859df1a77edb635553333a56e3d3c4cdf7615;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb8a809ddb8d964638e3cf65b24d0906419a74d869a26be6313a4681bc769cb7e51401b9f7f9cd211a09bd2b292b1dbd92f4ee7de37dcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a2c2935b657011c760dac076a68110a3a2b63473b0ef2d9b730d38373dec88c93dbc12210c48f5177768e6fa04783a72191a888485288;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abe523e7b761ea79bea524015f2353595eeb3be1d5bb473dfaa26683f7f0447e76b244aa6bc0486a4da7d1fabef0394049ca575411db3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1d4d133edf2a1e6a26234775065491ee0aa359281228e4ae80784aca568b13675636b2cef1ab21069863455d7311688f9e1ff86fa44b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131eb5615ee8da16c7535f7233cb7aa74e12d7e6a3bb9d497ce403cd53cfb8f9800e4744283ee7cf9fbef6b56e508ae28bfc97071d20d6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b7d1651ead82971c8dad733fa933a231c703b9c082e1e6fd8ebbf0a77443a72888d722ea59e250134ca57c239c3f780b86653db9546cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d90773c40e30853694f5159bb0a7c9f000b7d0b64da8b43185b9165a4040111f3c9da32325de5a99f8c77e70bf7fd08286ab4725f6fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13430c223763451ff249fccadaba40b4541ac2bc73c575a36f58aab305f40bc9efc6da5aad8f3620b0ceaed6c46d3b479aeb9985d939db0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165e28b3a3adee6f5c5b5ebb9512d0bc86e2ba5f9a7a99130141946a49f3d9140917f5715506ce9370061ab0ae36d5f067154ce9e7f96c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f088b1063f07703d60513e353ac11b07c8127852ebe2bcbc0c70d3da7a529453445398ce841286d7f163d9a110b5759f6c2fa75a92c65d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae82715c32c24fc0a786ba5fed0002666f822d1ac192f13ec2ac11c65ecfc21eb9e96f0d29ac7728e9c8c62b2edf53d5fb477582ce8c18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b237485358c40361f1e23f38a655cfef55c8abd31143d0f64c1d8d4879563ef82350eea05ce9d28ba067db5dcfc8898f9ff0f3a41ab5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1760ea93599266426dfa39dd8b763e9f8fd6f2687632f7104054dfe4aa2f396abe3f79cc1da304843a9eaaf547d1806231ab9d387674a89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1056602233095ca10cc0e17bef1e94600a6ffb677f21eae2400b888fab11424366394ee686684365da9e37ff70313f605ca5fc068f034;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h999dc348c9961fa4726b2cdee60508d6f96e35a27a5b8402c97c62a272efe0ba71ede1c041d81506b6bbd4e0218aed91a11d75d5e43db7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e0f2bab4a796c26d9f8788c9bbf223bb5d2d79a898b4007329d47bce87b1fbd52008e2b064bf3b31478e35b317b067b9979fb1ae717a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h810d518f69ab22b6c45f19759ba2580e6aaa0db143e4bfade410b3bca52c54309007ca08f34305c660fba2cae27e134fdcf8cdf0057886;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5bcba75f53607d6b7324bd74e51b6ef829e05704f179a93a58eb32a18cd35e9a81f897ecd367fc84372e07b0ea1e98a4f3978b35a4d71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179e2f2a3b13dbda5f9afd6faefc733703783159a3a1a5a84c6da57fade5e687054924113a57503a65eb139492af5f4592ea06f032c4898;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8bbfefdccf8b0bdf144095d37bae3852e4d32318008af1a364d24d67eb7e0417a476e888a229ef5f3a5485e1af104fad29256a2fff9f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141f7fd8ceb90bb140e440a8ef36c828784f38eccd604e1b5807ce1ac65335771f820a2bb809c805d3ad5c00edd18cd1d5522e273891f9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103210fb7465713f1363dd9b5e711b3059cf85ac1f8d36e474c0af48d8b4da9b10c030acb65f577761ee7607f0898ec5b199df99643f8f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b9155add9bb261f388b9f78c4e8564be9106255a33dce265f488bb020919739c7136c8dc9ea6527bb7a2391863fc5f5220343637470e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153c2eb1b53715f08ba12df5bd4b8dab5bfa8484b4825dcfce6dc629705f78c290aecbfbdad6163f5f45009f9c36a2ec1fded7da2480b58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7abe0e126493d220aa1fc3a2b4d0b608f3707272d65d9e6bf473cdabcde1a0e8c26c15e4d1f49dd3cce248efc7a6a497df7182c0ef8a0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h679405e9bda74d4306f292c1525ac0c50535646ca73dc78df3c08a63a4e53ce8325071840bba43c69d7c3f5590da41cbb6b41d964c3b16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd33f330401f09a43c1fad7a6e5502e57f6ce85d6dfff5e80c80d76d0b49aae65ea240827d889e829dbb2b72ba54ef5e0727a71c4fc7573;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11340d8a116b2dd813a17668c9cb7277ae3b81ac87ca64d18674576b454b03f01a15215aa48a16e79a2a6ad398fd4b3480b9fe9c7c4edd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4f195a5fc8cc6e943bc41d9046a2fa3647a80e88f0c398c2491ee62d88c10fa3a59d2ebc270af6b5c07a18195fb54e32bb11536e679fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20dc319de6e2da538410a5346f7f9cd11a705d0f1d2ae6a9f9fd5c9f1ccae2913d64fae408101c8b5c65c87625b93585e0b20696f912c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101eb925882e55a49653e32bf5a4676ef8d0a764acfcd08f7ece81f25f9c165f964b8309d25fa2025711997c480e4e3f5cbc01f17114f70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d4f31b6bf960f787f181ea81e02973f0e18e80a49dc706a8b9720b0dfe4db61567e1c35bb620783d615c9eff1fc0e0a3690c275a80b24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14146da0d1ba36956709c395f90a86ec4c3b0830951dfb990135217dffdd27303fa2c1160848f70c1edbb4661f28d46dd45bbad2e5cec41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfba1a73a196d06e2efce55569d650e195ca6cb4225f81f9872260f243ded74d67301d02a22b82d56cb293cee22cd6011622f95a51ea2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdec8e00f7e76bb473341ec4385e3b3f9b28dfecd7e69a21c868db1fa27c5c4702cd34b71d30de124553a32d242d4fb48e7e95dc61b6686;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h68cb46cbd37bb2cd019eb19be0ab0bab4446abe4f08200d2b1450457740138cad5ed0c3f99a5559e8e3cdd28cde8415727a2ac7ff89d82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f57bdec05d2464651b750371319e39ef0620634585f8a417de176c94f6e16a964ec96a79fffb67153c51d3754718668a7f2e3fa19ef051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97586b405cf7886634074384478e076feef7ab1f62ec97b0bf673e11e247607a14b4d11317223dd3097f6989a06b508ceed1174296b375;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b38da1c0ba99c158097afec5f811cdf23bf5789af9cefd56e34662c767b58acb3f6c2f1505f700af26f8aedf1d839d64c0e698c1fd2bac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2223477e6c71271c676f7747a24e4fd737dde03c847695a5b58bedc0aa2449bcb10e125e6ac732387fc698d9cb3f02254775cf0dba006;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafa5e8ab6d31d03a3d0c82c1174a607d9ecf8e2f4e171df2f5c3ad7fb923895a27062adab146b0244e4d39b1650b518acdec762a88eb87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8208319cfb587609e98e9caf56f09eece4f1ccb2050212d9466435d5f2b3bd4d6cfabaa273be56293eb8a519b745e281ce780243440b35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb37c1ad9248da526c9eeaf1ae64ee5e3c4cd6e72fc79cefede20204c5a44d5d67d482383f1834de4cc6424337ea049818bc10c47ddc9a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8dd39849865f6ab502b62a5abc1a250a944726bef8c8f5ec2a7e7a5f12b04908a52a01dd91e9b39e8daa96b2fe27db431588e48cfc9704;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f3e9f9d145a3c94b582dfcf5171c51814f1306f49d5213d9dda13ef2013c40fb25e1ac9bd18eed8bfae3edb4ea721d8fa6f8be32d6a75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4096a01100caec5b22eba7ea6f709fea2dd60f9a462e0cbd41205759a79954461233a9207aeec00de933def764d7bf2b11648f7a047d1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce3a48f67e21db371f24e40bb52e21135c4963892c17cc13d38eb2f36162a921e061d280f69929ec61dc7093eb9cb5cd599e5e27bc2824;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c63f0db305928830abad83b7e7181b5a64eee3283b999476d6bdeee8ddd16c7748a97dfbb4e8edf36a4529d37c31e5bb45aee00e8a865;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64eb14c0eccc8ccce2aaf7b931b3436d205c5dd608dade4abfb42967dd765c56c809b7ffad71963edf67b6fb6a56ce113b31983869e2b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187622337d87174ccb608c5ed3dc17f5d6c3654ae8d3b3c5dc58313b19206cce8ead25c825839f674b4c40e4ffc4c878d71a97c01803ac8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13909c27770ff8421b7a4ec1e437b6bc57316f843ec60a7e5fff9c798fd3580aadbaa9e3756e047ba411035b1613c85e3a71c88f5929aca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9bfd1e9e08105e03e0afbb23c49b1e5c1b701139fd86591a25868f0db0c1047d31139da201480706430dc608ff86b090d55f82afdd9f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc089182c3fff5e011e0140fc6c68b8e0948f503ecfffebfe200fae9ac81c7140f3a4f3918d066a3bb5d5ca2b973986d937d85b35fd85e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee431caf3bc8fdbda7cd55901f5697a02d7462db303ad6c211d0317edbc114d6a96a1c40b6dd26b2bd7f7d6407012e39e571b85222153b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17950fbdc06a4bdd056d786ef7ca132bd19c782a1a4f74b80aa362d0c1c18b462008c51c56a91c0762603076817ef616db36276f5708ab3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1ff7f0bf6852a99f5b854883aa902c898db1bb6fa4a549a2ff070c2bb545729e53a3718ad6ddb31519bea0b853b963b7f4236296a1356;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hace5d6d9ca0fb43713b84705e0305f8dc3fb0b6db8310f8fe41402f5f46048d354dd45d1457620b5032a248f8db86222ea870e61605516;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c788cfa914818d6c96bc2a15e680e0caa9ebdd2180a7b56932dc558dd2602e0f9165ae023bce5328443e1784e9fa9d2f64dbcdbbcdf62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h216f135255e12cf3a48d01a2e56ad70084ad8f61f5f544e2293c31b0bb0170d7fabf731def19666536195b4dcefaa048b3fe05f605a1d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0a61fe9964fa50a7ac93870d4e3fd5f5b0b9ae1d51e1c1c02ab033fe3f9dbfbc14e39185bcce522deb7e4b0a7d8f56220a7dca879bca9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ee77f04c1b3f7604c127ad69ecd4356acbbc15c823257db162bf67c12928c8dc47b662211257e2c687b6f41c4a480a515c0ebdffb13aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39ce414efc0abef4a2fd838547986bdd39c9c53326ce99d4b0ce0dc477749d866b2294e56c5007d63974cbf90b3f7626bd3ad98d664e10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c38c785ec1364127742b0c93215663057fc873e6a755c3ee1e3a5a4bf1071875848026873ab0183fb42549f885ccfbfe8fdef9dc09afad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fcce781e2482d95e147546cc2f2eb123119f2f97d5cac169869a7204baecae4ff1691817b5723171e53ef78c584a2bfc7d2dc1c1d83c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h437025de3cf202281b9609a6ff4bf8ee91bf5a1b13f3bbababe0a174800fe455fe14049eef1e5d556a9804aa0373ce7cc56623c112685f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde3aeaff9f238227afa7d4b8e646b1ccd0577c4e4b43226bee6fafc8962f98de13ee607c92f674b7e5f7a0d8446788bf50033c986db3ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1862e4d5f69f7498493c93ba26761b69b23db93b2e1decc23f56a41b42dea03e8f7fe602a71b3b11f808097e70054d36833c5a2e7407e9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cefb8ea5ca89016a479fc93963d906a1369481d13bd0f615f577c9c16ac174de6536629d52a957168bee5d2ba36ee9fb5a13ff82b4316;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dd347e49b1f1cec906ce080cb6f614c1b84d269d495a453ab1ef955a3fd989cf0639afab610c6e186fe9dd28a98f71e0266aaa8f6f9eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fe91744ab525f9d7244c417d3a99505d3e04f8806fdf34fe0be061fe6591cbc48d91fa08cbbbd3a57af89f5916612c164be202981767c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125bbb54d3464da4bf2c926bb2fab17a3ee55d51aed933140d2394d289b4530b78862807fc72bf03ac2c7fbf0a42755ca458158b1281529;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1102d698440c83160aeac5a10abe1069c5891f6b40bbafb422c8c8ecc067a62abd35cb319068794126f770ece27ee851dc52f6d08d93f4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef755b57a12ec8cbdd0d0cac5a7a585ca2b124b346876491ba90fed76e1045dea42592d17a6ca54d1ffc5059f50690489061a3f0de8698;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21c5b68316e207af9e496be0c5f7bc1762160b3ff4b69a555978f666b2fa4b20b01f908131c59abb7a1cea24d14429898829a200cb2b15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc24c0e5e7bba3806f9c748bff16b7bc4b0de6ee9d41b1bf1798d1e3e19e0698c26aa05694a4f7b03a001f294a0e28374d20f7f412208;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha38f8155df15ad48c525d6c10691ac72d12f15ce21da8bb2fbd10d1801c9c77f592df749d0c5e0ba1cbab886faa42db6f48d784e52dab6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1945ceb00f52c18b8b3092669a3432ef51126c22fd7084c95c7e11e20521fc84e72d903a923b47a0b2d452a4cce2482049af6b2397f1a97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63e03658c4c58a89c4bca46fba16dff35434013c02acbb392e4d4e97a542d2d0912814accc495071296d21d33b27f5372067a8f2df8cbe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77b1e68b2c48b6898178346ebac1024e387b1f5f14ca7949250c48bbfd3038786a01e8a6ed9fd452b129505e3deab16d96f39e0544bddc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ebb55d66bfc51b1e4272cefe8e2095aafacee1ad55be0ecba378c515d5ad49bc6ef6384b6d1f10eced5796c0bd8b5552f78c69696c5e86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178efe8fe8009ad9bfefd8034da50d2836f13f12801d0dfd79e0d9ce0a6b400abd42f818a53c5a1a58ccd21c30cb38d021425a16e7720a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf6035cee210bef184dd2628320db2a929c6ee831042e2daa9d5d5ec48ee38634a4bbe882b6ddd8c1c526590eee075d1eaa0cbb067b29b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aeb3b1aa905a5dfcc18b275be70f9078ed1096eeceb6d6f3570bae6672208761e47671519b50ba1d912ba18f6323c2b8cefc5194976396;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46d9fa72158164946c474aca9efdeef849f1a899deb84239630b4120270c499350d1e36cc18af1be6275ece6012bf5f127016284ace055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6528b638ec9cbce7db457924bb66b76a46a3619d56926cb80b2835f873e8b6ba6ef1cba50668abe362116c077cb00ac4aa249fc14df6af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b766e6948aff220dbb0e823d7bd8da498d6973c88976240fb11ae9466afbbc3548c468272e70c07d28cff9894077a08bb8ab9701e19927;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ff715bd9ffd0fc4d00e16c4c2818e6aaa7f7b4e2526bac221cc19db7b89172b53ec92c5a96412abee8e27bca9b021fe249b1ec2f9f96a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f08743bd3732d7efabf9ffd6a472078da589c8e682e1ab3562fc963e154038ad8525b0a483ab7d1f1bf2bd15b197b3e042ecb389bc3d7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc0cd19d5f00aa76bafa3bff4c8228f1e2c9e320bbcedd68c8f06c3944a6e31ea2c1e969c9888bfb24e39d719352616213aa781af43b29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he62fba8c32e4b62228ac5243bed084d46429baeb9d2b14dc64ab69a5b0f4d1a13df5f0bfeb6b2a748f323426e71ad6d5f66de11615899c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127680907648e370c17e58d1c580f3ba96302f4bf502b0eee2c9104692b817b6900f40a6875f28df15e382a6a100d7e5bb74d1ba5cade75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61cc7884ce0191049f678520ab429d779f2e06ee5f3ded7ab0d7d7198c646579e23660948ca0477dfa03865b0377aaada172e273f99438;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc042069b364b3df53dba206df916461bfe3699f51cc4e1f335000068a3838c452a46f1c59cf13132c69c592943420ef21acbc1037bfb8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bad16e4c4ad8b1f53e8fdaba36cb6e74397436674e225931196a271d1548dfe459fa2c7a7a9d6e650f4ec45eeae1d58f921dbe2492f62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e37e1e2ca47ca13b5d7b464d5daa8d77be7a3cf47649ee72d9d85cf05e038988a0771b7f4c80416c60c0c98c61bd1dcad9e59521aa100;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7576e59de45e89466ea49d8a32a5ba5fcecf86568241b9d2d61765507887c99a740cb90f59cc8e98e4c3bfdbbc76a190bab2ab850773f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f70a63ff006643ac08d2c98aca9cdb40a5acd81f985f608e9a978226c840b4326276069ab062dde5aaaab5d580c13f4d1e2b30809d9d72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8aa913f69ac464755aef1f6652becec707492cc8506a5ee67059e7010be1ebf6f031d2e15c149e2352cab1f539f7397e7ee21a742e3e4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c7c297883d7b5fbd5cf2b991c01b2cd36a5ec7902d229eb2c031d5dfe971b23223564a72d4a3edab0f21ad03e9bb10a753ad7a25f13ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa67172d601adb97905feba88401ffc071c16e1ada904963fcc9d491a3c3e28dadc4b70da53300a0e38ee1057190adc0af2e24012598d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9b5b59d26cad30b3d63cba3e50a5def83f025764543cfd6e5e16a418d2797da13534a321d1e687c2460e774303289836f0e62d71115b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1434d306d03b612ee00efef8993dac129790e5f572aee36201716ed0fde7b2533b048ddae7be60361e1f410919acf5b6fcbebeeb0ad0eb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16888d1d9f82968945a7474b838899534143e0ef0cda249fe7d3c1b1f51bd2eba3862a9279cdb2ef98e44d592ee95ef5e7a86e646e6d35f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b3867e96925aba557402d1ee4bab368e67c8150b9e62ae917dbe6445776f436b0670fc48f5e499601548956e4fdf73bb2bc02e40534cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd2faf77203d261102532773d31dcf0cf82673446152ec2f7d9a0b7a32bf52d4001f395a1b5568831e6f7da4b0dbfd10ee5daf6d046a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bc204b17c12d32f3372a1e68e0aecd29609a3689ea191bd5b9ddf2d226b9334d240318030c3e4dd03050b525b31bdbcb3ba0812667ef2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f961685042240fae484f47b049ea604345ae0a662a9b432ba267b83c0f484ff08462461ae69e1db97ecbe384e5652a933191cb1c22fc26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f69d66c5c20081910c4fa65077a6e1433eaa3b39363d088a7b440d241e73edbfc4cfbfcc6a205afec94b5780b43aabee83c84ed378987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf99f9baddbee2cc33b419c87ea250982ad6ecdebb785598923b8fddd60522dd31203603552d544f518d1c5496bbc1061ecb532f98d12e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1810da378e2cb2fa649b7c767b1504004ad164bdc6214465b488c4209d0ac607a21054f0807411f22d3c1d4934c05155468ec464623fc2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120fe50d3531099eda9f202091e04efe9151815a01ec5d05d216efeb82efb1d097c77f5f4eab65525ffbfbe3bedcfd4bbd6957933512bb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89f5a7c4310e31b4b2bf1cf1c1070c8ef0194a19c7046696c5019a468930956ff50edad8fc4ea1eda6f3e4b18e8d0587d042ebb821ef73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1537ff68c3b41be9d0bd909e8117b9c317bc3dc1b35110515705f4a479f207ca6208d1f69107ccbe0c7ca8ad682758b78eaf67d7f9dee96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1252f788d660a956248c0cab537bdcff7410906ec9abb019b7b162b63fbfe2b1565520b629e84968885311b24149ed49dd2d2f2c15fddf5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4c79070c635811cc005f195bfad33fde706725a43291ba7027397bd51cec4b488c347f5ae8ca208f14a54d102c4104c93558f7f6c94f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14aec71ced9be68593872d50148c2f851a4ee80f106d92d7c9a15ec42b7b0efa3b8ed116ce126750171b0a2c49ac9192369dc8b4a43dbbd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae411ec3b1612f9e716dce482965a6d23807de08190110d7b7e933ea830a82dc406e5b4378cfd3f192670913017f1656d666e298afebc9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182a2a697bcf2e8dd592a5b18ebc613b5558e182cc15e98be27b6b9c22a49b3bdfce99224accf10308c7e6a72ad6d1ea94b4b67d5997881;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heef1cf99c70d66dac5c72aef2eb643b5ec0bdb7444d479f74f5dd4a21237908a3b8a1bbca2dc850b2cdfd6930970bba14238a15bd9b3c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d2b4e2711bb23d849d5be013849d16b159befa17b8593bf2d98678dbfcf346d8d788364782bacd9cbb995e2977f5f05eba0bad1462946;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bce19a067cd4f6bd6a13a8cab8320111d08fa8066bdd002b220b9df4edbdf2c3682768151125b0de1c52b2114808a38255207b0b80515b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61f3597d3cfe73b481d385de47484f5bf0d687dad912f760186f66b02d975278d369b74b5e0924bda7380504ab3f1f802e379b57c99cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha87f36f38e23a2c1b73fab95a326d02f3a7f84f99a06d49cc8124034ce3dd7fe21c089d2d86972fab7b10da8653a575daabb3f98a843b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0f21e5f6b94fc9f1e07bcb4f4c7cd1fe0cd765719ce2d215fe000e57a885e478168a03996d49c2f3ed63ace8cbc1b819ccc5d70d402bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae0bf93d0aa3dcf3171049ce0fba68c667904311f203649c16b9cd61b833afdd5d1182b9b5c9e666547429ad3cd45d08a35315d7c0c8d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4754f1b06a4dcd1042f720dd6a022c819d2772d10f5695c8df831d55249033b3e3a71aa28017a15843fc97b5fea090ddc32bf3875a1577;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bfc30d7f9bdbed7ad7c2985fe2a63e760b4e0a586632f96657df0dd8ce8aa63193c5812a24941a6c8ff55c03cae3fd4e4619afb17e586;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95689baf0ef24afe7a0a3ac2ca2f8ecd7a3ac08f87dddc04673e973dd5e2a58ddc20cdf0d913fb5a7388f18e1c3b69c47a129fcc646cb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h961dcfd963d4d89033cd24ae9c20b6d435528bb68ff6ba90449a72d597fda0c106c00bff6fc8aeec3596295cb6ef7f083b21053c95e28c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfff76399ba990894298f4cbc978827baeae6a0966c3c07094685438a6a6a3cd9ba38121ae5368bb544dbb1df7785fd291df1c18e59dfa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18894cce999ad7fb01cd833551f907a09e03bafd6849eef4d3b07be7ea779ab7c7c9b21483dfd726f72dffd7a220a53a416d4fef683fe64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e729c92ebae0e8daeaefd206e99f0037bc37de7f7ed689eb89916fdcd32d66f924f450103b98e7477675cbddce1ce9656881e54f11dcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f5591e9113486ec437f88beb0ce65a0efacf7e967b1d3b7ab5d909488a80b7d1372e042689b37445f748a561258d9ecba3a7feb1b042b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14649aa2612c2cdda9b24aea66c676f7c2b680b1f493f7aab9ae7333927f2fbad337c1bafacaa8d969a8c37fa9a389ef16ad186997c8978;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122131fb190baccec210ad2bfeae7276ec48829025c5973b51de840dd7b5c1ff18ad0982078444c4721d593f0e5a6ab3df37411b6355c24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c36dadc930170b8e02a10017e9350504abb422235dfae86fe678f60ca7bcf1e69b851f4b4855011cc55ff29950a861e9a3bdd80df4140e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdbbc20dd9068ddd403f92da3c8de79be91adecf647b72e99b42578de2b8b61d494fd835fc6981fa3f3c28cba8c6bb38e6eeef1f0fc51c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f926907ac98d745d951be5a436e3fb1454cd72b3758a44fe09543befd0940eb9c0898717048157742455a831820df35f7a68e58aee91ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b895dc4e0281c6bd5cc3445f378335a077cc94a0afe1aac8434e983cd5114affdc49729e6337981ec767aa2e4d1bc34f75343fdb30196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aeb35e2cb8991706fdec63ce04fb8966f24aed3bbc71b713cbf01511e7f1d9b68b9527e622f4f4b0acd6ab127f960726af4381dc18246e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cae3e857881adf354b68207e548e08bca216d30fe7674ae15ff343b2da2d7cefece8fce3b2b34da506f1993df70b1c721ca589a2ca7f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0d66fbd8fe0db2d6c654858f6af3cf0cb6c23cc9f35fa2eb53fb07cec4e79f65ac62ef2161a080f7f06195ca6ed6f7c5854198057a94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha03f19bdd94b38a6858f3218d4c5d1247a002e011e165adfe499db450c130a0eecfb386ae9f831d764dd40496b63d6347a0973fdb071d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87d1db41de97f15ced6ad02ef17c0cb9f574ff15c8f45399239bbf4872c79e7b12c56f79cfbda962705159c3f0f77401d1397531bdeab6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd9ddb1d52e6a4545dd15da71ffa81258c517fb77b061251aeb69d5cea04f98c54cd438b363911be7c335af235c886a43af292d0b1b842;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he27e5d105694d39471569ac5f48ab348bdca6ae9843c436afe7ea66c4e5e1b0ea96d28f45fcf7fffc4ac65608b38973a7256d4ddf446ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14736e023c73914252cef113e60ecfbe8820fbde0fcf84ad19647df1438a1d6bab0006fc212bc0ea881d1cf1e2d212688a71b86b52ffc79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1077e017aa970e5dd166ba38303cc9e206ddfed859b559e3333cacc17d7f3f78451a7cae3c6deebd35bc3db3715941de3d0441650d74a12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2e687c7fe271bec915c0e389a57864f3dd668178b9c3ec9807168bfa2ec50df8e89f0c29b1704cc99ac11bc5bb2c0a9d5edfe45723828;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa0323d2f80f9b61e2cefea237f2f3ab17b1c01a8d96508ed39f6c0b406dc47946d0edd3fb7693d43fcef61a9fcb54e38c4ee0615ab293;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1920a414fd125205a5e53dddb87c7aa55eadd1a2aa60f4ab5c158cd6dd047662b2d181be36db1c0212847d2e2ac12074d823b35c52cedd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1489799e6db1788f6ed113dd2f1a186a5ff42216b24ab9e579ed0c54fe8b78946105b74a8509b4d10e6052c6c7274cb7bfe6dc6608d7ddc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d5c346d5a7f41f6223abfabc967449bbcfd57d6229f5773244ec3ffd81634e68cec747cb58db16d23ed38b655770225b887bd298160f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d308d3060c32b51c163ba12efb86d49b60d93aa9dc064c359b94e0ad5f9cdbdf588c8f2f9310d62edb40cf35328b4f166f46c6f6c8b85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f20544e6bae6ccabe5c1f1de386829bbb2d68c0214d8ff45a0ddc83eaff9941b687e7696e361615114e6ca4f8ec7660af1275597137078;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0d35f702e41efd2bd177b695cfb4569bab6f61ab089c1b9104c4e845c19bc159776818ebbfd6de2398c326860f64cc3a08351fbd44a0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b9a3297d7e050de7a3d17978cf067788c1c78d72fd79995c88b637e3070bb43dab900f65a14c72e66a72c0d55aba82858beb4a4dc1db8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8a823e6573511e3dbfe8cf1840338f9fa8c75b9b52ea7930de7213d1ffbff8ac2894cae407215a1a27a9c66cdc3c41604c500ad03ccf5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h215dc3ea077ce88ad4bca70414b7bf35108936de70c9984c684adea80e80bcd7f5bab931d709a0e82bd3ed3f09176f938048eab2bb5c9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8ff92d9d302c5f0fcf04c0b2db553ce8e943ce8e2463bbfd4ce65edd0265b5ffaeff4bee837dd316165d46e52f973e3d5c32e95a3d377;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7126b108f2495b2f894b3101f30a79b381c38cb507a9254e628ffd5d5604298585fea33310295a2c22dfba7f7fcb439f86afd0bffd5c4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c1feeb0b7b44b1d388005dbc722177714936b532c3e5c1e9e359ee152bfc009348fdd2c2c669c3507889a5aaaf61e21f766900b74c0b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39e16ba1d3152ed2fd3390db3ad6128f91f33e7e7b20be0ab305607a6c97adbafcf4f92934092e7dd23c8d1154b1cf355662df3a6212dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h681916d3a7e1ecee77073f15465a6e235bb002d167d9fb9b8baf5c3e16490b56b295ae6644246f6f4ba27131fb17e5dbcad70bc08098da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1179b2c56a2b18f14db13d48a816510acb21621b9345cb7f0d62f5e1c3627c0373c02033ec21296ee314151e0303c7198ea6ec269085953;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ef7695eea635bbce31612c842147538e9b1435ec2d6585f90c8f84f48d6901a27142b96af1ff04f2b04308af8b70800e01c96b47cef08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b3ba8d705a23aae7b7d028ee7651b4ba7e7da0643658553e8b6fe46488d8e907fca00f914e2727fdd51cbcb527906c9b4a5ee2af5d0e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126da5777f92f6071253e19ee7d1f7495d3d246efcb7f6c45171939fd5d847e0ae4ae840484aae016cd532dcaa7d3887fa4f0c5043506a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c6cad2450d02b3babc26a2575a773b673f53fea3396a15c5a8b1836a00e14386b6ccea62d1c8263586b48be08e3daeedb8e0af7ecd8a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1041b4447164d7f749fda99c082c1c98f26d53deeeabb99f197404ddb349a1a83bf43a252ba163005aa5ef9724698556ca8fe3259dbfee1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd99131ccfbf3a1a5e9acf2886c44223ed561a8298405881c5a982b56d6ae0ebd304ce275aa92a10d0cc8549575e3c20755f6bd62e8297;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1782b66e865fc8d167e2720ca34b5fa3a22135af0e25e4b8da1f759ac917b6b7d13dc5237bbc224bc4ff66d3da128daca4960b2b72d51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d2f064f3940722090f11c5bde442cbc87ce88edf347bc841e4e5ce26dc2cca75a26ff0b727cf814f7947ef34078bb96013304a5df6034;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae3801dba46230bffa215c7ff2b4d91a9eee006d27d7020713074c79643820d20ca0e443b0e59ee482dce51d270bf8db5ceb8e16ddfbfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b81c961fa8b140f9a92b4da8f3e983aa30eec8d9c76025d090deeca89d675c982bafe1b4fb7130588aeaeacc0ddd0a68b49547a9e19f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h887a1f45381ea41a5073dfc64df242f6a8275818f799417c99bc06fe005a7b28bc91850c27871610a1003aa339076175cfaad5c1e88858;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bad353db45280498f75032bc2d168bcd9624e59d26c6045bd3ddeea1de6834b956cd3b9e47e753560b2ebd4bfc6b7de7780545a847e52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169c0cb86207ff023e17b814675f091d70b55696d85f49197d4d2c7b7f49d0b0abd6350137e0514d8b257e160dbd402b3ffe304409e5a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h606d4b4bf048c5c244b2987117bb668946c6032a551ba522c091cb4589540bfd36d702b7eeddd1a35152a528ec5523dde344f9fab0b63c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha70d10106bc0d427cd7baf2a30b6e95c26da924e65925e100aff67527bf86a2265c5c80db9a1434a222ac021326553b7c28a844903ed19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5e0fcd6a92470b87f6e0309b98d34617eb31e64aea0f3f01f16414a888555a6166c55d1eeb3e7ae11aa5bd1d5fd22777ed408216d4f10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde2fc25ff9956c902b59dffdff7610b4354e8c0794205fb72ccc62d82adeacaa09a4563d043d376da47b28456417cd370b5a07630678ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141fe4a81d932a5400246a588b8190b00c5ed2b8c9ee6d99eb6cc9583941ba04825ba62a7d52a9b296d9a1e072b377c3742121104e8a6c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb2b279145d9960582d5acb6002ce4930f76d877f680833ce5e8163e1633e47f4064ecdae64d5f0b773586c71ee8aa890ebc2ed64b551f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106378326cce187618405d93bf7437ea51833e8eba379cbe4814464e32ecebd3922c66d9d73da936e2b18cbb40a126f0d46b67fb56a2855;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afe7253deb71652b75be090541b440f4030cceeff62a38e1f9a9d913e2131bf8ba2f8aa97d5c97054eb0dace96fe9af205b630b5cff4f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18497f179a69ef87cf40a29b750d2869a6445b1d9626b22e2d060f49dec99dd7c049eeac00619aa9598d686acc324c8ecff2eff23132fc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb437eef8add9c0c6053fb6fded829d258746a2f0f905349d11e65295eb330a1e8bc4d73acb812dc148ace9dfa7676f1a44c44639ef2254;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e050c4981e392e8a7f8682d433fe697fdd411539c3dc8599a40f3b21d07bd3735a57c45e6ebe37da744d7d680689245b74d22ee539eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0a3df44eac63542170843521c642b78eb748f9a8f12f792f7376b16d3d651ccdd08626ec022e670393dc2aafe3f19a25c52959fcc120b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he57578944a9a5a8f773a0778a238c43de0fc979c4f4c666f6b1dfccb98ada03372054dce2fa82620067110de1d1b01b5d7ad321fcffe24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha18bb8beb88459cbd88669a9cbb2fc6ca143411644d19625efdbf0b2710345d4d15055e7cac0bdda2f97a459036b72c342fba498d930b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166705bf5d0512442cf16fd2f17a196da9a001ac297bc94ec065fc1a75e6cbb4f946ab87767f69369e0c1b864fd2d719b033e67b1d8d77f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he182a6e973f405e8be6c62b9b02a017a1874562f001ed0d95a65942fa238117b30d6361de77cc15fc79f98436b82db2f64b3fe358c849c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ebe01da1a5e5fd3a2579b7dab89fb4f06071a48590e2897a15ac53352fe07f1a4fbced8355de7165e11ce4c6a5cc8b5c46ccfc55aefcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc72d175fb10eb2070b315b34481116e8d979e9bea1cba96f5836547d2249c21d12d88745b0663a511d7097cdb32a029f104e793379d47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1590435e87a38f9f55dc8cdd6074b271f84fa37573bcc97aa0aa109ee6f1d388925139d8867cd415dc6d9e9e2d64381bf13674742216004;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38b9752f07840f236999d19bd556a0b25b636dada939d2a8d1c1ad627af44677acd76b272e3b8c70d0a0c5f4f54814baf62897c04b8150;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161d224f594ad8dd9635db17faf730099b9ba305d194e2dded0db35d69edefe82307bf7f235863b27f6cfc4f142d29fe1ee2f6e68e5214c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cba063a511b71ba315e2d83089437c8581b4005ce3b21433ed059c4cd72fb5586db05f664dab94e0716b8ea261ff7879ca6524dd0721dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76a8a1786f2f46f8a7d3e6859fd115bb377fb30d989914794858d09200469cb7470cf7a616096981a358ba496704b8f686e7c28044e70f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f99eb8a6c20d53bf31ddb8bf8617a0c449dbdd20b6f22d8dde8b42479d3086f0ca4a7e2a3ea7bdaf4da2244d9f1125d8e4aadbc4f75bf9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a8dafd0344c02b897fcef620f5bcd746e2233215f8c98bc7d370b23d63b861a863f3be04b1c7e695cd387af0ade69464d3827dc1e5cef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c174b92971c67aea4c2522d0277c7b27a8840283b68531493c9063836c957949764c3c400f040e5afd7e6aec6dc72013c28753d610de4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a903680d7bca40425c2c37afab98586c188b1aec4d85fafe49842067fdb64d04e23cf15e4633a92b0ccf53fd5d95a3fe67f7483d271606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a8a66e0d305241a7b4eecaaa90be833fd2ede81691838fe5b6ad78d3e9cd0ba4e726f56fb461fe3c465fe76e7a8ad76e1ce6a120138b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5bbee01754ca7628018dbb03fb56b61942c9d44e90171462dc1fc4aa7148611ee11db5a99d0e0b9af3b965566821d87ee931a4bebf45b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ebc52b2dbc8d5e6713c53e6a6146cfba71f43835e7c21f1cd4e7e2df2f3a33f3e74cc61e7311b475b1ad4fbc6ea03a72a57a0859b542a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1905c1cd1feae2e47b97ad478b959769fb913797ff61fc72435c0701721497ccaba00ebb11fa425e5dae129e818ba46f183555a52adfcfd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1994913f5c7dad9d3d0ca71b673a64db4063555a53e950492f55608e5a42b691fb7ef63592aaffad17191f9bb3cfc1e2de0f6b8f2a4be9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93246523eec878f653310b78b9586f72e37e050ca1957bdfec5a22ef7bfd5f9dc0683291ccf1ca0fce4426082350a656e74e06c5ee186e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba54ea16c4b867ae1d116d269f6bdc6068dfae5fc9d70a4317b8d7bf4eed596408100954900de9c548504098a7ad007b947daa6dae97d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c3e2bed62531cd917cf9600a8ba8ef55a9b6759cb3dabefb6da02e3059c1b6d4212d0b71cd96b6f3a560c473c65618d3e24761a383a39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6310132a6f66f1343409a2aefbcbfe6624bc7d3fe49d26ea097e965a75cf4151eeb61374b233f807d80849d5c0d538532e1af02f4dd935;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he463463beef45faadcba72a600155db6ab8eb9dc6673dad30b59b31ddbfba34970be8fce38cfa92b0a2debb90215180b3ff32a2ae6f787;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1953788945f5126eefe9be09da8bf17e3188181b949f09ca5499f1e676ddc44f8f395275012c0b673365fc538bdda59a3030cc7d0150f48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109ea0078eaaf3cfa36f24a46db6d312cc676b897aeee595e87bf1d2045394d4a75f1f583177f6f0ce0238ae621d6896309704ee7d4dd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d60ebdff5db82a86a74163bac29807a401d3ea29b52486917e6f209994717db26af71bcb0f13c73b8f8b5812e136d59b1baad1435d61b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f7a133270c859fd266a13afe075a2bd7a0c416a20c1fa25a36e5efc5e845c83849359eee91217b411f595042c64009168191797181ab1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1340a9598e9abf0d034afe951457f57ca0f5297c414108cd67781ff36109731b57501389a9476389966aee635b61b4145ac34bbca8ddd95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4f74dbfbbcbcbdfa72a531b418fbf8648abce3907182cf79b5f13eff368c06a0841c1cd9ba90ee13c2eb365edd2ce9beb6671ce564524;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa7fa783c3d713b47138872f5c6e1a214bf0fe995e7d64615a318388c7ac52119bb041ce7e010245eb8b030fd3ce26c1d11e4b3e7484a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24047f4f8b09ceac9ae96de5059fbd73ea1137f504cce005feef7df876228400be11b9eb3e41fed72f29649064926f2573ba598213e4cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5e3b879831f683e47318971929551bd81879e2e4ff5dc1bc34953e5be72fd63ab87ae6d6e31e840b6828f2011b332961723f80a3d0f71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b365696967244a98d8556fd560bf6baf43407af439af1c2ed6e8333441661e8f42adfc8ca0e79e29f8ad111c465d0a78a20ddd4f474faf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1f487ff523815034f27c013ebc323a3b02fd488e2d4ed08b917c8421ab41b8f64db45ffd5b58cba3acd0a6f0b30ca08eb826bbf643694;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1018b00f17ae6242be122d72caae5ed60189be85a3b83ad0668fd5fe0fbc0aa0e78edcc267bfb7ef9ee7872a032059d2af554942d92f250;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h720f1530386e978a705160e034ec486b46c0847b18b4dde2fb012adb5f555c444b401e1b833113f3a416637955d25307309adb657398c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha29c95169b77790a8db00a6cf54b53873eb1b4778b96e524c9cbfb6ba2c8b7b5eddb8c43736d18741a2afc85f8db24a5d29cb97e144b17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ccec83285b2b981aa35dcb91270aaeb935509147839ff0a082245fd527b39466b8ba1c9be48afad2d925a6f18b777e74bdbe4da75eaec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f59fc1c75c7f8ab2769344c52cdee9851c301a54e6656bd09b824bc3253d5c9443d7f6564931c15db2a6c2a77ba2a11a4f9b6c71e4acc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb03b5081aa59f8cd40298d6e3a2da7400611ada8f38fdf9cf4ee0604f8bbf4f3e2eaa987498df439e421f8d7f6887bcccdb7931b77bf4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f59ea1b96a01297cda1f09606de20fad896645c5a6b32232311dcde4ae19541003f019fe27b998b405c78f2aacaf92c017fde8eb2effed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156644e8876c7e0843bb825514eb088b4a8847943899727d62e4829dd24bbea39badaff18a8b33fe551ddbfb506d944efb32b6a2b90ade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13086aa82cffa909b2132c5b2a9994d6721b45815d631cce64c3bf780421a1b858e047c59a68da77844f152d81a3b2f8b3d71ca67a5c5ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d737c2da4ea4a5e35b75e3fe8607801ff03071c4a4225bbd1f1f97abd60d434d78e11668e4c1dc6c0fded48e5d56756729bbbe256b88c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12654a599c1dcf46d11b14e38fbb8f445532c362a98fbb71598390f3a291f738ed818e79589cdbd57d37824ac51c8badb3667d596b5fb41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ed208ae40a51efa5e54dc0b0b2e412326fedf8a63e593a16ba2423ba4c79c04be4c32e5c82e0e18cb59ca5cb371e75a99222d559264a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15624ddfb26cab6e7d1216329caa93f6e813e44162a95f78862b33ab38dd5b1e87d2caa6c55df441698cd9b7a4465072007675119396e35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197b931e3623341205ed0b7758155cfb1f9a62d4ed591005be174f9c2bcf36907ec3595a8fba9dfcf9ec36480ec82c76e671ec791a9eb90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa42637abc8b117a1ceb05d315ca50411d7b2acfc9c1641cd366c8e8ce6795dc2d6962e8f8869a78cccfe1982dc5e01fdc12def23d8086;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f774dfed00e093719223ba88858414186b4eb8a15b82d8ee7e3cf5c3165c724cf2a227d733de6f4d229b197279c4b624ab7ab6b83e169;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1c05fb9464fc32294ae1d823e14de5be87649964f24f7eb7efd5536d54206a66c9117292f1708ca660d931499b36dc95e72541427d128;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4aa2a537d806e669ea9b5c56c4a3b9bd2afd55b1017050cfe540e333d1a841991df12fa00dc56ff627e9344dc0fbae05240767f6b2399;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3aaa5000b6e3c0431d88661e58e5da787ce768f6e704328c5514d004740affe03e5a36d4e9d7e2937fe3abb75058709b0f6758b8dcce04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187e014ef6090af9893e152735775faff455e3ee02400d8e3c8cddf30ea08c2000a05e5ca9832df956ba09ef107b253c3e39af8695da7a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c0c92d39cac8cfe5e0bddb2ddd0c4a3c4d6cf81a8ed2aeee617407f200587df3dc46c5d5d96a549a1e6a5eb34cdb6c6d7f963e7b6d222;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf73f07059e60a808dce0bc12dabb7bb17d2325e90329bc575ce43c4fb739bb99293d11120bb5c8332d41be0b5a6b5fe75b8c0a4ba92ba6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1503d80bd09041a2a1e127ae46a4a08772517281b6dd560974ec3ef7d81db2b7fbeb9f03dfaee504d80d2abc9e012f73a0500a00929162d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134cb6209fe04c68aa5ea7705ae3e94264313a97af6f1a3620a5db0df5f86d38e5ba55fa218a292576911e2f6efcc8d111d7e7bd8877f88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dfc0bfcb3a997e3d3215bc9ad9ab1b0a2856e15d1772b8c597a1569080b8f650d441dd6965da502e79f5b57b32352e1a826d4805bdd82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb17e7f40e89b5c391dac3de38aac25d6008542af77970eaada56241d08860053da88e804f6d51a1e51f29aa2303eb542da87f9a2477aca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23cda7cd48f9d75a6235b8393b8bbf00fe6270afc9972414103c5c1d950e8b4dafb24993c6167afc6e241bc98fa62595ce8d83733df9e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7e599d77fca4b0e3b47ed368813130cae5d548794328809523904f9014af2917a6c3113b45fbb6b2214afde6fea0cb80ae62b890c27e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111526bd960496a02a95d5bb575bf2773e0833bceefe12093c99f3c9150827ca835d337d3f3ca9348c59cb988bce27da02dd7de14916a9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha288c9baffec4a56f29c94c4074249d54ebca7d7567f0af7c6f966603670196ce890c3ba558bf9d3a8c2001c3455894a390c2bb29f597e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3da8273cf71bfff8316fa42b2a37e10a66c8b99d485a7aaaa46bc89c655e51c1c99b857b53613f728d1a79f155e8b5cfe26f7f728616d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1972b3872cea48c29fed90604dd962d93c8fb22005b9b54c9ac629648bdeef2e0f682ad467d06a3a1262f86dc2d121909a5bf461af6c264;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb55cd296a0e5940ab47d0ab441676895c4f95ad9828dad337f247e98f8ae919bddf4194467721f826a4622cb39734ac00ef3d3c49f6e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha073cacb7a03c212c76e0f0d73735aa247ac7dd5ada2a8c91488336fa888e28f7de543945b36834c0ef7eb7c8d4d0d1f8fe3553c4b6e34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e985c65ae3aac487d70f07a54a36112d2dd532c9e022eec90b4166d34997f06abfbe03ae07e5a4d3a2a8c2371d5896b57f47ed502ce273;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67f8cd45f49e77615c1931cc85f5967592867be895b8146fc6989e38183564eb57cf10b9da65f1160a176a59bc0332d89dd826278352b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1236d46009a23770b2eaac150ce3812f6635c7e3a016fe0fa55158cb9ee4416abf0430e550a8651f163992ec6d01ddb0d70993a36b878ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a1a3b94d09812306fe98bcba0da45c8a59d121abe41da69a0517583baca20fb7b3813bdf09bcc8a83ac58d423b47c258d757aaab33bb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb911b20a667957cfe15325b1f7d8a3c7c7a650656c5e0803b4be191530ab9003917ff9cec5667f014c6525b5a338997b79640dcbc48454;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7df747113c71cd2c3185495f3317eb4887b0316f6c8cd155b1348e6bba9457773de60068f37361d5ad926e8f551cd23e2d57c2f4ba9c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf7561fd9c1556eaffd857bff4f465791320a7dc532c8b4303bcc9813e749e371166ff1e591b70b2b4e765d2c881008b8978e943494069;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1424d34458d5a4a24a0250779818f43e48bbd6caa4b05d52478c44a763570f80e79b730a51bfc228ac36e2aad5ce85f11cc356f99de1759;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbdf270d19cb4af904f78d350e6d7489a94a50eea1822e824ee97253cd2363d00a1af581115ef38d8bccde939e4e7b84aadd51e839ef72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea3313adb4f9aa3d4f217ac382aabfdec4de53c86343a68f4f5458ddf91c6d440633cce58f42d4d6dca8f929baf169aee1494b38f2a68d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127e4e77bdedc97b792a0dab5c5364deee89519b4e8eb98e550ccfdb8002071a2c7c225eaf259dd8564da44b36cc5a5e1a89ec02b1ba21a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e16acd7489a4e5ec229d125082c8ec9b8beba82732540e8ff838b333d48d66096fcdff3164a765c663104bb5a6c42ac254bfbcf7beb666;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18355ceb0655756bba6961f342f3bbf0c19ff396db2197ac0211122d64a600a198166c26f0525c0329d62cded618c15c1c3c75156186c53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h115f9048ad93fda0f4d81e52454a78819092ea6d98eaf2727267f7ecef345c02c893f947b8a6897a461cff5c6fe18103d44f70f481ca13d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9262aa20b6800b81554cc57a1211e0a97dfaa99663e0660d625035816bf390532b9957e7efdb51298392bb1e7ef6cd6bfeb48325e0fed0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h393495b6248b7b65c7ce228db6c2e42c18847405ffd77520315af0e6aab8d6a92e9a63b46196e8d9ae64a213c85204e6ed86cb35f25f65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b6bc5bf223219da49879d926259bb1652f2fea2b7deae79df631ed9d81bc37b4e4e7be556e3e60aed3925aa7ca5d056d24d561f523ef9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce34c212941a84e243a4b4cbe57a81a301e236369c41abd52ef9183ca75812e0ace5e62ec573a047ece818e329683bc7ee4fb119354853;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14593f69e87c0c8aba419b2a368967f227190dece45458d2f341d4c6b791b95af99b69e7c7808eb0a8150c0acd69e7a30eda2226161edb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h320d1b0b363bb851d0ebe04ee7a9667e4e298c6c009970e882ab9b1ffda32768134519ed8cbd6132c84d1e4b7fc7d045fe76e0d94b85fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9648eadd50de8fdd94f3b20e4d773594ab02f7d973da37aca05b9806be4904980fe35ec776d5c5fb1ec918f40148c1468e213058f6a9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5c994e5089e6e478f3239a64147f55f3b27a4b50ae502de7fc6c980588b31bdffba2837fc0f32b816b336ca20211bbf8c73275f6e4fd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca72c01810aea822cb8a5829df6d060097e1d002a8dbb8725e6095ae50acb3971a3a94ba12248bb21f76f98df9d74ec10f745a2b45b44d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d2bffbba367d4d3e0fb31bc29e2cb0ab5234653bbae54780a89a8903f842060a05b8bad277e7b83ae3ebdc91795d1585a3b7567c9a311;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186d7729c9cae89ba6bcb78f7c4c16658da4931622df31100c8dacb5b4014074dc4c9dcfdab666fc89121e351ffc9e665b224bf39b54ccc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ecfa2eef7b23c89a1b06893fdbdab658c9e718922a5a071d6eaa6198bcef191a268196b583c848ebab0ab697a53158d8634fe772cccb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199f7cbe656bb73f1d43f39fcfd836e16318f3f4449db0cb3d4295749f5a015692fc6b59038830492483ccf178d732fd392d96c1cddcde2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1022dde38780b6cf8a3b03419f74a8e64d5e2c0304ac5d9a1fbb08309774d5b7a153e0f43700dafa61fafeadef0f26c60dd63d56c79b8c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b7dc242587ed5dfa484e3b8f093a6e180739827a4b4ee3539cb1e9faec5551346a2efba8d919203cc3843b8ee05c78fc184f1994cc334;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c34a2e2816075d44adbce205f3be8b1bdadb6e19be68ccbbab607a1bb602cb9312b78d9ebd44bf0af2067762080372226ed7b58215037;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a552ffd356f76819367dbfb76f8b094e594c7cf18321f0fb4db8404756f1a9fef815759a73b32c0b0d8645311832d2d30d1bba1216e9f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8629bff0368dcecd37a938035c7c96919ec8fcd6207c1bc74b7c06cf575a3b9c43fa1577a0cceb5a0efa67c0de99de3d619b5e788c0e53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33e5659c7da52f231a352fe799a4eb95463dbf738f5f4c37ea58b580c87f425d8dc19d3594e696ad5b8acbb9b920731070131e9fca3f5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a1e99883dc9c122ab6ecb86efcc16cf3f4ec1110a3e2edb50a6b6d39ad16d5ad0fa782c422d2a3fc902ab41541626d94ad2d3455b48ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc0b643aee0256f449e2c6b060da5418102ef99c6ddc76d279683a596ff93d520b77b739be11ad4464666b001488f9dca9f4f00e1f7e3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81c7ed19b7000d5e3415cac3b28c409a276ed11f0f322d0c2900d80d47315dc97e41c9b634dd013b8eb4e284db42628585bd1e956bb6c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4861ac1244c955c73599743ce720be137da3a3b4eb2d487c17acccde5db575313823d3f1fd0aef67f4899d6bab2a7187296228c2cfb4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6c4a60c72f35075adce1f9550be4fb0bf931e22dfc474f73a2e7a5bb1f5f042fed629a54403312bb7bb0a05ca29e2b3cce609b130e3ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125c9bba99c2693655259f17d56527df8dbd23145f19aa3e0d7e1f440348766f4bef589cd0fa8445b3b1969d29c8045b92f9c855dffca9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c96db664b468a68b7a087dfa4148b601a3c1c645fcfaa5f1dc1a4eb9bbad0a10351e11af5ac5bcc5da09fb71cc8d9a801a9f4d28c583f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f7ee4aa27ea315e24a7728238164bffa75be63f3b71ba89b4188a976f452e587b54f4274eb3328fef3761d825ad8300ff13a3d07698b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5f5d814335a179f01e79caab2ced320527c03265af96dceeaae37868d916c09b9d8807a83668a20867faef908c197f09bafb5fd435d05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95fe4f78ca6e5bca16a6063d6d6a3f822437772d6140d779e83f83a7489300cee1000daf0255b693c3d2fc2abb6548dd5ca0227a03f01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16fcee1453daedb417831a9b55842b451349b183830015a735c05bfb729b31aa7a2702475dd7300caa293bffb4da9c282032fb634c781c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c42a600cf7a75129f5be5cedbd6e3b6f8bf0a8cc406df74a523ac184437b9bfaf9d8f9e5a4ae6f306ba443d439436338395b24fa61a6cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1109f39a124b513189ffb53c30772c72f55d5232ab05f06e62cd77569e671724c3fd2a44f85997220fb0d9b14a016cff8441b89098bbb7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aca6b5a297fe8507902b3e06b5ddfb3e388f11e59e44c955e2faa96eabd48cd7d96030eb7109d3865b218914f72274cd91b3f8ad865b6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1914530ced2a30ccf28fd97677695ca60e3c062dd658ddc21bc15e9c5b39330623cda96f26f59c6b662bfcdd2d08abf1b038e2b1407660f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc47ee949f84fc403afc2104c73287a504d7d2ee4f345985550c37ceda5db223d1de6c6ea47f15b1c06a59735051f3b070cb3a1f5ba97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21d48206f7b64d9c4f4a626410cfc4e61f065d99387260f53f7784b77cca109fa113e5e4c6c240f88e6aef754aa088eaed1caa845acdf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b68077bb70f76862376432fc3b94297f983d9b12ae69cd3641c970c4120bb45f2965a8ee735c5ef946691271ebcf34c7c332824b6d387;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h654cdf666ddc2aa96c5235c4e0cfa077c076c79110319a31193487da0a13e6da4c3b1dcdb4cd5d37ad81bbe908f790f6c4568f837b31bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1df46c3f9c35320d3f91634bc136d037f252db01ce96ea426301cea77561ab040e0c31936989e1d0102f9fbb84e564447d8f3a4170185;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc623c9f948b7a8dcbee10c7b2a709a19e3640a94636a8147ebfad88f29d68f838d1c3c21c259e680ae9cbf69e4c7dff156a77aab5d69de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0ec9720118ac060a8cef22ebbd1309745e1e3e64d0e6ce127f49548ae4fcce8b9b94eb4b797d8b32684113b8b52fb1e5c6598b62f3980;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h143ed3f1a84e28fc62d82c165f5c50fb07c177d9c403c25bc0a428b5fcb6cf6dad0d5357cb5edf9db5340293ed50d5f08bfc5bfdc5f68f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b57452a4b9f480b9196f8159bd23379ac1a66897b5487da0ffb8ee41b76df0ff3f80c6e9548b649b1e841ff89b859f75ccf78b0b633a9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e60dec5f47c2cc7ef771855401171d81cfde3e2b3c343908266b971fb80284431043733e62c11e5262a8acae23ddf66e5b149718cd4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ce130b5bd15f7adde17ae3e43d9b8280293a1d518175953d35b2d123ea6932118876f5a764437cccc01255116dc2c554c930a5726cc05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5efd0a0f80a6100d6dcde803e913a3cee661b9712c9363e64db098a74e76b2abf4c39298a74e7d21700da3a22b72f47b3474e39c7c36e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178b03197f5167bc03c3a7e5414016377f48e78bd7016feab2982d81711237c691a657c5ff77500070d883f6c61daaa6fc5f8abd8370e29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8d1dde60b7698ac0a5d5df6150e540d37fdd07ad3233504cbbcb8ff1330cf47b6eb0b3113324d2fc80ff2874ef028a60a17544736975c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ce2b1e4dadebe301ba21975368535d2c94fa0284962a207c6b3c673270501ff3bd2a821b22f2e269207d141595d2ebb322277f3f33818;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1513193d4cf5e0216465896dc1ad70f21c4df98b80ff36824df86e6825ef2306e498d09a33f863d3c842b16f31093032c91cf2fc75aca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1309ac726985461f7684f15602c7a1a13e6f45b8a734d329306c020e68745a123a92cf6160b7a1cb9c15da14c767bcbaa18ea221dc788ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10562003198272702c054dfe572f18354f0716fa724b2f82be7c5bee25e534338e563020ddd87b32cf0c8e0a1b65522908cd1944a861583;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a834a8333e8c8df200fec20ee0c96c40d1e4716d47e139444b09305054366928ac01ab1cdafa99060529d0d9e39c1749ced1c5bb94c657;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64ff2123b3d5d2518b2640d5cc45a04b2dc09e256ea9003bf86474e4eb2bfb1da96599928c3cff747757f20ba855f668c57bba1e2d3ac6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9165b4f57b810ed8aa1ca5252a4fa485bba3993d9f7560cb842bd85da4b974075a574de0d4482e94f576d48d0070d804da27329c99cf96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c935b179d31f78d81f81c84d0faca3ea7cadc9db8939d9bdb94434d2ecc3b41ffc92d67818b6d11dc77380e01fe5d2a5fbfd4f48fab37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1530cccb1b6333e3a293ce776b317ed6dd06470981443846df1ee184149df4d37a0f20284b1490a998d43878598b46c3551aa8cbbb6dc1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1092a936bfbb817e0ea75195b4be4dbe41701eaa3b5c3cabf730e28e255a61743b5220637bc12d42684a1d2547d4b764ed97767dd5b1e8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1412921896cc94c71f3b3228442ef4dfaaa8dee56e7f1235368c39f6883ede593bcbc5cb7b13597596f21f85358edad27349a7536fc3760;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150bc69ceb8d3047a053cb98aeaf784c4fb27cc6029c0251101c85b15dfb553360e7cf0f897fd4ff414dabc9fb77bf4046b3a9010b6c571;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd72626db085c1a0299315dd7f1d914463923c0fc390a485f53150cfc10752bdff83e797c31ab5f9ade6a946dbe710693665d15f51dfe2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cab7607a77a5944045c8571cad6e9f9c7c5b51858e71839a44e78020fe76bf0551dbe346b2fbaa08118b0fc8df7bb77d556105fc9a2d05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9206741b5b4d2f3c57f6e92c2508899e12723a997d39d938ce99207ae93890d44257a12f10d8a6a134c3d6dd5f0460ca63983e315e44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd097a8c86f6e8ac3056c5075c200b5d115d5ce7124fbde8c0a7619988d6fe1202589eede4bb78bfc4d3721a632d7f9f17acd8847a1ae9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5e3bb2232fbc3f422a5dcad30065e55329b0f24ef9acd22d462b6e7c7df2f3012c35cbdd4293daadb607b84219b6b2c4788b070577bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h378ab37186408dd41b6f48d9e10c6c046c7b77c5a3a69fa7c1c9461ac2bb158da2bd63c3fd285ecffd1cae8479657acb14e12244a12bf6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b259413d201089474a63989e8c16b697539886664e089d25372c38be9f4b5f7645dc08309bd972974ca1f3bc2222542200929f10dbe024;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46034742434487e455436e695ebfbeab90adfdb7f317e27fca289e8fc0d72fdcc9f8d7d8c45b73604e7dde2326e345a2287c241201f64e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16abfb5a597bfd17d2b5a70d5365229848fe9a887bd4fc62ceda03327b6aa2700fadfa322feb2c7c44f7c7c374cacfe64e0c48cef627559;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he672921e6f3d3a6a027b21b6721f8ed8cca42ec735a0c8bc7f580d24c5a03644092805d8e278e9d6f79f1b1c266989bb0a4b987ebe08cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d173f5f5d3e4337f3ee3eecd45cd089418897804c439ef11d6a9fa353d35844fea9e990941a1a39c6cf5a27935ec97949de8fc12be28d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1357a9412101db25f9b7530a402811a26d0a189a10123107fb266243d788affc7865d2fe0b30340aaa9372e31e0b5a01ce0d05693465c1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141302e6a69e9c7c40ae4c0fc76c758ce4aed0cd2a477234589259ebb1715fb316b96cde1745e5ed988564974868ad77f2c9cc9819632f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf35183540a0511a242d76835029adacd989d1589b665cb5353a496e255313ceb8507975b5b6da936ed66bbc78d61ac10203fdde131148;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34e2a2d265fea50f124cfa833b0422a71396437c5d54b904d3d2040947a8f6e5e269a3f42cac36f6b4e6fc1b5070196f36282d530484ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbb34a38875b9563bcb5ad52d981b50eb62c45be339f03aefbc6c0d54d841b9ae933b8fc0655c8b6fb51eccffb6556df2d3385f518055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166ac800c98000b058e29532a694214be900cef5459041dea0c41fc75058c4c0a60a91a7514fa3008af926cc753c2a310204471f8b661f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16869f07977505fe4d5008e1e4541dec637d1e2abf50942ee7d37cd7a449013b58ac048a4a9f08967dea2ff571508c7f818c170b0e48f55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56e622674306b603dded64ede73ad95409adaba2787d305ff5451b38d3ebc185954d4c4ea8fc1789d363a460a014aedd6693d836aae144;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101637aea8cd30a85239ccc65420fd9fda0af96482850c97ea54fd63dde258b67e869505b72501405c50359637c7dc376ed57def4cfaa75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5612e33fc2d8063e7ec953a371fb5338483774240c3945e2b20d896433d19db99b629e8b7824683076719f241d6e653f428a0bd76098e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e216e1ca89b12206ec57264af7a4944923e8b60d480f462684d3d51d92c74b357e459a11e78c21e9431638318c61f49dbf4ef1e02c5281;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193bfbca6c872715202e27e6241d53ca7c3709c50167efbe7df5d6ec9f80d0d24ecd348b6fbd03bf6d4d11c5a8614e5a0d695becb15c85c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1016432b54107430db2a891cbe94b9a33953c6765ec2dfe3389bee04e5e765781d32627dadcabaf84120460ea3c4cc02d2f30c1a22eec47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62a44396fa7420a6dfc0970bdf7c210055cb04abf3132e8198cd60c3dfff0ae0913c3d3187cde5e86effa18cfaf34f5f5bb3d897596f8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177711371737f4018a6c4ce104a0a1f7e08c5a8abd00db1eec8eff00e05554f7c51f0e1ae0f9d0a2e033445636f860896a72f991589ae90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9c561074ba8c549af2a6eb55e7eb981a2ee6bd0ee32b57451e42a46e5329c14773a339bbb934a2ede75401664408d1c3a41dde0ef2434;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4371275accd000c4e495be003abe94b8534cda8a6910a9e95575ef3036505552a77803a75664798a1901034a05948436bd1129b1058584;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9834dac1485c456fa4e2b8f7d3b7094d99a7acf1683fa5423d3e47e0b5f491f01eef96484f29ab0cabfbf562624f56dd2d3966a035da3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7884ff5e33c2aaf0866f6ce6f7c604981dc0a5cc70bbb7e6407a6b5a3a573d0515d8f90a78bbadf233b60c23c3a6acaf402805d7c7042f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8736e6fd6f4ba4a893c127b35238e1de88fc7fb5cd98de5504023585ca68b3011f483c606208f5d4eb5197291e96a67be422924f040b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h431028eb93592f7668c1b654364caeb2cc864607a762b58bf8dd45bca06d98fb8678247fee33c3a1ba955c49a0a28b9eb07679ee92f79c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1624475657a0bff162a310e65db00a8710ca9bfa4afc7df45ae5e60bcffc597e45bb4c7f6f961af84c4ea07002cce872af662c4d2db8f59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ab4d828b8a8ae8ec71e7606ab47cb5ea33dd4b5b79661f94c56e62d328c14475d8e7ac60a2e326e08d9c96a9e99242dee7a795c095a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba31ee989dcd292e02d8c405bba1d7535a282108949e31b411a78270f8d3f0141cd5f8523fe75254fa72bf202005b7a85f9dd1978bc481;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h294982e9c9b158eaddf8132e215dda1030a73baa1bf2958af52e0764580a9642227e0055812f81d6ced3dc414ea0c4b7f5919c6e7034ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb93f56c51e1eb7f9b9054bfe3ae18c00df46460b2b7cca85112ae61f2202f14e8b116f0f544321a7e74dda36ff75ef72c518a011e74825;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fcc5f99f601e044a47e9ff4f80cd91653d6b15a30fc9c5e36eb70d0373bc66dd0241349ba762f7a9428ac5a3b7565501d669b22b48377;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c6b6fa175add2c9a1822a6e31cbb009c7f906d2e84c291807daa663324c0d0c57d4c02e15256a968eb03f0d535335ad2cbafa0204e17a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104b16fcce302b34a05c4f2fb398eabfa5ad73d6e44957bd5ca76d6ef5f2fed5536f790f8d961196c8e5a16fd58e414ff71ea2903ff4e12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9514fd2c9ed20482a4651d522f20f5aaa98eb6fe6d56c9f9514f4c536fab1422a4614df5d48b6781dfe0a71c5313c577205fde67c22027;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha285e19468190db8218c185c7fa18ae3294825b5e2c8000694cfe84e57a0cdc40a1df6c0e7d5c7e66dda825cbbcf23b85afd7475d544f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120c0fa61dff527b93556aca5a9a1490ca7245c526e3a43b1ff0d4218d2ea15a21fb9dd50c6f43dbe0a0fe1818c23267701fdb559ecfe29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11184e9c475a67732b43bc9f5fe29db0f3fc09d4b6bcc9da8ade2eaf003c18c6eedc6533c28851451e7ffb3c111721b21131e81a3db349b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8a2a3dd639616e12fe7254e5a595ab54b5ebe6d5f75c86f90bf5a31e679fdf1ce8d589ce4993054e0bcd7c25ac49cf2e3fddc0b2b392d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1326a05ef685e14f2a726bacbb04f7ef76cacab738b386ee874755f403334b6d8de9080787827cc5f156429913d0fcdecf21c33a875727d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ade0e3a56643267b931a535b60e5d3366a2f755fc1ad122faaf8171b9bbfede5523e3fd8d4995ee452567eb5e05516b0721ce9251c8ccc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89ddb610acfa3fa4634e716e447c197fd7f2f6bb8ef6325498cf7b3f127c6bf29e8b5cffcd5b2c3661a1d531f3328f1a7754db7dc62627;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39050dae866d7f279d14fe6fb9b936e69f975a0acf811b169905656ba64d17d22c044b22ae7b53f9e5ecfea4d411743c192650cea6b3cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdd8f1c2135a5beafe2377a5015db02b5e52cef75e3ddb56b7ac186e2e5e1d9afca0fb6f81a43dea564b55f53754b108cc92d06ec49de9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he053200197288dbc6ed2b44ca10430a4c321b06f5f4a939e89f1d607f6c2c6c8c4c9404829cd81e89a3b0ce89accb0122a004e52f370ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b4ebdb93c121ac82aeea3b48405f92cbb1a967c4ef2e6ad08dc8dd9021edeb0e5f55dc11e7e07fed80e887d1e3276a1e232c299c97206;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6bb205c0cfcce29a9c723dc2c8cf115f03f4364af096fb60fecad25c845fdc8b866b836a3bce2d3f5e8bab8459c6d3a5e8233328056fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40128f7897b8637c20ef5ef246a86312217524b2e6fd33690dae1659aaa6419f0200af62370c23e98ee5f016af9a1ae5ba254826c8d19b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeb5f7bd48bc458a52f1daf977c1bfbb07d0bad5e6f8cd7146d191b2ef3364191d5a66cf71e511d8d4dbaa8acf87f86ff03049047bb9cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1996ee1017435f8b5d598f15639616eb6d5fcd8941a1c41e8809c75588610065e766c229674bc58c3620a0b9979e874773372f95ee2508;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b7855032076a61be1db36b75d0d5720f150ae3345b5fc79569bf682919970f8949f184763ab8e38b37f6f3895b1e8e08b38b49f04d358;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16600dc7941f7aa5ac96ba64d836ace706ea96e5f25df546b7bf86a0fe7ab5152d90fbbf6f04047408442bc5325331d274589fc58dc5282;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed5ef6cfed2ba57b008a1e0cf2f990f472f4822f100ea69f0bb38cc848d05754d055bf0dbb4e8cbca5cacc4c73847437528c48386a53ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176519d9d091d80ecf859b436126f87e7fcdc27bcaf12370d8fa020f26bb7e2d9bb1f0ebf0aafebb413fecf16de6d20d4cd0a3bb4dcc63f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c48306dc2f6f16cab6eef8c476afc48e207b84e382cd20ebf77a80a158a78b95894af0acf72aabf2478b6cd88d1208b5976aa1f3c2826;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfd5ef09ecbfbdb502753212e09954f7b563949335e2ce3e98bb545e7434559a9e214489c778bd57d541f10d5d9f3d6a814ac35a421b18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3604f9fe40d2255e64a17ed4afd6cbb3ff7f9db2e9e32e5c587eb2ac467264bee4a041e463f563c45672b2f617116fb4fcb069b57f71b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0bd187dc4cc31d29030a9cc62a304f07570887734ceb71f4b09b4307d108cec3a20aa8729a11dd1d917b4dd339664b195da3effc4989f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2f33b7d17d1457eaa2d0b3f888263d14cb94cf2daf7c852366b73ac6128b5d3f0504f5ec03e54546a0be636dbca829fcb379387898b0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fe0214513b16d5de11597c06e72fcc99977751e8c0dd74ac4edcab11fe5e708713e7ec22ceb1ec12bacfb9e1e49b70c2ccd09a1c27aa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14cc2388addf9d9ce7f5ea0dc01f122391853c795373106068bfd8b2961457a465f48d17b6a388630330b4c0eb5b9e03f253ee2808cd773;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd5dd72352f79c962a369007b499f13f87c387b3ec8b95adcf8a9b76f315978b9c8fcbc32efce1e6df8d265a1b2115a8c7fcfaa4966fd8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1932076524d7dee2ee4fdb2f697dfa7deb7375f42f0fd5a2a870822ad6e34f121d9e229895e7efa5f3edcfe6a94a75a98c46f3122fa48e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fada5ee42b85c5d730d8f6ebe3cd8c83b6fee436085a9d53092d5d9bdc1f2ca2d11a153e26f34ec6d45b0f0a9078e43cca22ef611fe3c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1dfc8882ea769c26398e0c8549a756ecfb225d3298871ac78fe02b5a5b245d4e1a29c2d0bf693310f709b1e8fa7781ee7eaf73f28a847;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e36cf0c9cafcf75e04dad319bc505f45bb238042538e392feecd6a00dbb78cb66794dabaafdba6524116768647a89f8b14dcba2c9b864;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128494c21dc1e427710921e2ec1d6130572e7942e82b52ef8f2f46565939518a1aa432a3a2f29fd04d564561d633d455d6de8f045e9e34d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57237f8bfc48c3d0a2204f25b8d6b02ba00a045b822ea28d7c71b4cd5c65c3ef93b97996bbbd4f3cbecd6760c8b7bf2effe24310b532a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c076d98d08d5bebf22db2ae68e6457bca9705eae7f98318797e7c1b35d9bd36f358d7f893ea0e5bf830130197b56bd1b938218dd7b96e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c74406ce8cd39a4d17aba0e3aba3c3bc70d0d83e4b9707256920b96ffc9d53f094f66300cc8ddfa21ce7cdd836ecf9502c490bebc1ac9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18becf36eb3a2f6a1bde81970767cd46a7f0efaf2413c841d3654f583cc72a97bfd6cc16832858544c3446d489b5af4c1bc56b55a6e0a8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h167c6e9e36fd284f2192137f19557429d496ccd48cad00d99272ea91bf5c5e25f03a6bc03e901c1a4d8ffcaafd97ebf5a946a62ef87706a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147a5ace8ce9993eb70968b26ca478a0b2e63dd19ddf9212c00166abd6be175c5c49beed5bf9bd1ef53b4acc82971a105c711755850a2dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ab915731dfe280dfab32d415810d8a7f577b56341404e749243909bd9f50934059204f21029f530b871f8bfe905a1628e07763976fc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cdb5ba0baa75505026e33418d229f1dab85eb4b3de7c0f8e295373f2430913f0f7afa6829a41802545be84022c1776da400535eb96512;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e7ec8d8f1318643b8e48ac5cce2d0c38802ebcf38b26efbbd1e8803399cd5b5bb93f6d592c74368d3a7a640ceea5f80faeba62ba906af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0128ecadd9f43a5a473e3ddd29722977fcd364eb1434609981c71f804226d517884afe0bfa279976ac99ab1ea59be329ff2c1c1aeac5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8075dbbdd9bef55c671ff44e9e92de15f407d4404c68e84293e1cd76a6311e88d58c92f5f38e962c6bd1d6618ea5d849170e19a7fd8fbb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa5c1529ee1ad5ad15a0558b43547b863134260894f6e130edbe8dc52c65cbe4aa5ae38870b579d21f82ba60325691513f32f205b48f91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3f432fb7961fb41661b8e905084cda184ca698cead4b42918575097c756588f2ad250234f8c3b276710b85c50b9578492db240ccd6bde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98992c21d5a864111736c860017abc3754776b9584d6c12054e91ec36082d00891c5ae10c3dfce02e3ccedf97b738eee187d4fd683e45f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1410badb39cf9182a6579dfa614b9dde39c042325c74069180f7c44b85a4f5ed08cd7150851083ecce8924fe1642a9d84a3d3398a23ebf2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9a96eca09c4761f4899b50baa831a83e19e296a29a121f03d782a6d052b6638a730753862bcf6f0ca591ab4eb6bcaafa3f85b451882f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeca4f601a1388df6f2469a709007195ddc00dec3be0205565bcb5a60493115760c2a99ffca199acf0ca83c28bac9c424331a063be1331;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcee89284eff2a47973b30b26aa86e76a08d95c551ed8b9dcd428d64e461c9935c5a972a05abc32eec31a4b40307b88c1f2b2293cd40b4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e7339657bed5f671503b107abbf540cfc8d3b9dba45ad7843c4fe2e7a2303cce6694072699961aa803a86fc62a83561e81bf35da68325;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e8764d567c7fdc21343cc8a33c7b51f3102adc91173d80bfb87e30496763cf488eec32fd633c4eb476c9f268c635d4873612b0b4409ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b30b30a9b6352bc829151910cdbd78e98208af296c3e80fdab9974d6d3f2f476944572e95198106a39c86e67457874530b97ec0cff6a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ad751cc0f4488238bc0c4625e9d5fb8d949d7130315697c76661e27d16be1b5a15c5d4773c94569532ed05d62a2f8f178c679db95cfe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccfefe285db00ea02d808370fe08399f89dccdcfe8f7598958c0ebca6dcc24da18e4405517429515ee1c01908c992607b8ded56a922ff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da192f83c8cf2021beb061b7af28eb87d9998296cbad6ff71646bc520511f5c42bc986d7a3fd570800c6a25c1596bb0710b877d88ce86e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163026d84a94eeafca000ee27c763f276d29803904dba5e0f58d424ec81e3c2b18f9ddaf20ef8753f1b5723ad7216a4f2ef82c01032cb34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142a4f79bba3bbcadf4b16a479bcea3ccf94bc3a5cc5261ecfb262f60deeff79ac73b841e243e450eb80c2b7362b8610d1c7d34a910d142;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h543d90970c257af37bcd53df60080eac0ec741ec62fac1f2736faf7fe1157e21005f84cd73eae520ed14ac833b07744d9872aeb68b45c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf981afa2c17a0e7fa0e2249daaf24d2c0bfe2e41f5b258ac3d652953938c923c9862fc23f81d1d1f9bc4d8e91cbe12df32486469f4ed8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee425313027a2623f28257491bdde13226761c50bc9d3cfd8635b0f92af35bac66698f610b1420d5af9452421dddbe7d0801f5cb50747e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e19ce58fd3d9c413dbe79a928eb81be1f5ebd5b3ae1367c6cce2bc80da00257dacd89fb5aceaee52bbd7d391c078f18bac660fe1cce52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d083c42d71bf7cbec3a163b5dfe955e6b0e265cdcf39ee54870605f2e896ba1f60455f056b44c06d35886c9d30d594a7a8f686b23e96e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2024f8834cb5d1e056982e6c0774a57d7049737c2afae11b3e5ad1c2141d09c2efbfd26802d252be83d02336bb2fe852d0f79c8dffd1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176ec6ceb97f6bc9d273cb01c552c7f83962682399ea7e3d815c2f733d23c32725cad9d5e253caea64beab474c1db1e3eb1581a3bb76959;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48bc8a9ecaebcc5654d96bd1dbd53f56492e09ac46244a1b7fb569c6252984bb7c32f03cdce58d32f4a559295b5c3c6ec90546aa9a73bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h502db4e648feb2612868296f40a58ca75e20236d545239fcddf9dbbf6a2f232a3442e2f186ec0fc7256726559b29cc4bf9125a78146818;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2eb7111c44d38034a8010030af591f8711e727c901d6e5225a84ec44239b7077f9d94b1a9248bc5aeaa74f25e91749ed883906cce1600;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcf1e2e7db54216c74339be2744a3180a1209ababf31524f1d3ff043342895c3dc512e88d7476055cc94be51585f930fa3199eb683e2dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15563408339e9f9072f1ede03cd513f4f9962c00a87af618ef183b333de345365239fc568193068c6e1dd785c09ae7ea8d354f53f5f4e9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1de9ce19d311d985c83c8637210ad8670f4b457749d99ec549fc4967b6fb2832236902480e92a5fea2e71c907a89b1807fbdd316a4efe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5e140aa4b6a18acd839dffd8981bcdc24adf759261a6d317041b306eacec74701c248dfa8b2d7a51e2a4d9e52e53b31381b2547f6a306;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1938b0fab1d918d534bbfc08c650142723dc140954b32cf35ecf273712de918ea0a1808b1311a84b014ddf6d0997be461c72355357504a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfcb022cc56ffbd3ac6ecdcf2dcb04ae271989a599a4db0fe1ade8bdc3fc6b5a4de28678972016e1636182fec073381e9751f8aac0840e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c68bb9351a1e53c4304dd5559648b361f4156cda5aa658b4e3f7bb3600f5ff7e68e4a7aab4381be9a9ed7fdffd169c27367f28b63d78f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda949ef91c37201a73a7fc02cd7d1dbd431d796374d1281ce8bf9f40cff67708ec2622560e765f1e956b72346a6397d022f690f89442e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a860e8a402f6533f4a42bc890c9a44d85f80bdecaf718eaf49ee0a2e54a90bca179cee071a4e0b771120b42c8464bda69312e0f46faba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9974f1221703a874ffa8471a4239a91fceef920b1f82d9a0ea27491081af00b571bdab03bbf7ed13daf8684efeb2f0a4ebb5c860270d2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb1477d2436cf237723aeea84151a87764f9fc9e92fbf43d8905f85737121b83d29c4afea2bc6e66cbdadd0c840b27df3671fabdd8aac9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178565e5f739ac40707149df82c420163491f48f4665f9d27dcd680b34379ea8e0c29c362e5c59818a7f6c3df38a6dff042357129655739;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a175b14512d93be63dfcbf94242140b2f9ce53f94769a25170bd1b97ed4b2617bd318fa2dfce7d35a499a85e64fe96e75aaf277ae0f591;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e1ea9a043b0d114d87bc5bf2939455856872821b8863064df911beb0e6a31a0876d81493d1b894ed33db985d921d7049f914268a3a643;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152f9bcf774479ff584c98bc1a6be0af9ca96a06526a9032bcfbe9241f501ee855047689adb0df6b0b1a024a9d3da8a37f9f6ce562e3f5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1093a037a77bab6be3a1eede1e96b8bd8ec57ef78f49c5ce78f614dc1a81856e9b7b19f48fcc2f7447c6d31f959a351ebe9c6c283371481;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102bc3a705405a7e34a5e5f0e4cc5ed3d1b3bdc4fd9b3ca9734c4b02ec3985792840e0dce215ad21845f553a4a3121752c3a446cfd25065;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4de4e45e10fb2e8cc7e8d7de1e516106a9205620054f247173e08a09ba8963eeee2b163381a31a08ccf1400068788e575ad1ca4e243eb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9076d328253c3180131df6a2c765df362d11a0ef31f8cc7be35d38d2f7bc8368f76ffb87e00487b952b92a0e0f7f719790592e4f30fe47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a8ec000d7f08346bceca2e8b05751fe3222e43a8657c1fcb1b12fc6697a8828efccdef30a05543845acd193671c82c60f8ecec6185722;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d2a24b27e552a084296a3a386ed53365c1a4fff6abf97f3bb91de14d7ce276a63f4ce33fd49a7db68e22b98d330448968b4850ecf9654;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc5498844af929e5b6f6c9530f89fb375e0a464310381d55d745600bcaa7848ea2b74210ab75e3261f410f23083619b27a67457108e773;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87f81daa4166d236db358508a8f2348107233857c5126c1c72932a396296825dbd67b01c2b9dc82e7cd49a5e8aab3866e6148e3186a68d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd30b78fcf938b47a38942f2ff0c19d075ce29a39ed5b94c82c6a9cdcbb54eb8a7bcb578ac2e11548026cb7163fdac394d0b6b5793b97f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46bf6e5607994b4182ef89cb3c0854df39d1e9c542dda2d7a5f728318f40eac44b4a0c486d0cc8a3e614767225332e411cff30f9741729;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d302a398bfb839bf2bdb0af46067903314f9d4ad455b3ac25f296b309c70fe0c15519f16bc4e8ee672b3a10408162139faeb0932bfa82a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d70718caa0ae42c78b1a9baab136ccd1768267fbdee3a4a0cf463f22d30a8572ac6df83c8c84f25fd8e601e3c38baf1f30655e13316b67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f81b4e004d64cba09c04b8b2c254d202e09e4a4328bb787379569a28db5a1dee212bfad8fbde7148db51746f6c76dcf637be24124fc60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h917a3d2d40ce029fd045d8929db524d82595efd4dd8afc360e91aa49806d112025d8b732e90a64aec09bcd64c6a921a57df3d6a8b2d069;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1511c38525e91e8a83f4dd9ad4c0ec1fd5cd812e405565fadcfd8d76cddbc9ca79f83cc6cb686654fc990ab71799d2f028d61ad1f72710e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha81568cab92cde1d4656022808a4ef8188c0c7155ca8249f3d8cc0c26c91647ca4bee61a11659bb0c3afe0c2392094a5c048b497542d3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbd037891737480274c91bfe3d02a54a619999f5813f13bd595053c8345cbab185b404564bff5d98036da44475b10795fef0e1c8e6368;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129790de731785c885c3c5e4f83f5ca1b97efad37a9266445af2e3bc156f8831101cb29239b7d447de3ce2d550e98eb44f218c9e38c3e74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1e6af04bd8c6eed78b4c2e5ad3a30f09cf35ca7d5bd31d878c54476cfb8fb92a06ab49d2b209c5ea927a07079d1f91740eea1f570ffd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14561c45594c0fed543186d411ad92c3f39fa72e10accfb2cb3ae39b99b2fd108f74d110bc7d36f749d895b0cd06b71d52f21c66e51903a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc4b20dbba84456dfd4d237888cdf5f653a338c7148d858e6ab98709f8cd8190dd4e67bcfc97b1762dbb10d69e5b091fa2b298c4f59bc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd3161fb1c880fb874bd464972f2d6f35d1f81d79063072d574295e963f82b4bc4fa14fa02e8b0587b6475dfe7fa72a21afe455c6484b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8774b3d18f931add2570d81dbb2bbd9a1b6b4e5a2be81f6eb9577ce79a6234b06e161d7f2704060c0c49bf801b62514bc24b9512b781e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb8e154e86c311db4e867abefa8cbcae77ae6f6778bacce010b653d5798d57403514acbe9f777e3823f0d8ab7b1b47cc647235b4bb622a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbd936ddea0b351e597c19745b6d094175c98c166fd6e3433ef5b833d608087703f87b8135e1a6514022ca009ffc7135cc984eed299bae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e2045428d8f573d645e3b84588bc01cca59637dad79e05f7651e4e9a3bcac7e210c76797d419e64139a62dcff5aea737120dc3e1aaeff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24de9a6dd6acf3d5f44d2877ac730f2938cd877bf5e29c23d26c87362ef8afb33a7b4e319691b661795b295bf8621ba7ae5621fddc4ac4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d676839e8de987d307eeb1d1597108e94dbb425c16357a988cb41bddacca9cb1f7a00de38fba81837a2b431f1779b5417eb7e421ef684;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19875957a489f94d125a6481f9a01020999d53f2a4a8575a29b01a9264bf149354c3ca4d4e579350edd8f603c64a9319ffeedb827cf6f19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1455845f33c700a997c8a8205de93f54edb680b313db17f08d5588d034d84f1b13869aa9532a67d0478f5418042e0e49fdcac7b5a053539;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6de63e4229bf2eccdb2175baff09e357632fd7b6991711b361e822c41b2308638cbaadb9640319f3a22efb46678fa2ce12a4c6df8763a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac533afc1cc80efa0ec31d4c5d5faeccef3d4b9b437c72f04e907e505835a77b24665272992d2a6fa823b2d4f49d651decbd87a8d5a4de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d5c9d9870b355281666e889cd8afd04ec70016d7ed6cfc837976257ec571a4d39f1d771d5982a58e0f60823b8d383e4448cca12d6a021;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7329e34549379325f764d76bbb70de9927de2287861671394448c6b01cbce89e894ce8463366c8d7916a37f5e28d6b0d6f85f70e9bee81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1373d8f78dce7da9440ab3f0fdbc18b50d64c155be2742b38df402ea530f116397f1210cf039c10348a774bc3db43d9695a09a5fe1f1ec0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1655354859b4b00a83a2b8e2e50b46c87bdae064a09fb107ac6ef14f247671d67a4f89873f66de58f6a01bc4b14829e0bb4487c1202d8a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4414648bc4e07caebf45dd6efe4aef002861a3fc639b70c6525112135d973903642c3185dfe4dcad3bcfa2e3bc6fff4187254dbfaa679;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179bef0391c403ef69576a347bdc892e6576d210a27f3fe0d906534ac6775bc0843bbfabe74faf3b54293b7476432f9920c21154add03bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7395349583288d3d24bfb3069b1d431cd52a0cd3a231850620dd95dff0dabfe9225c82935fba51291715a539a852603ce91e623de185be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec5a9b2b43c8a5d8077247c1ee9dd86ac91f6ab92f356804c3780dac67a5caf22d8a08d287f88a95f6c038f902146aac663ef2bdc740d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b7ea17a822056a0a457cae1906391a7392a725eebbe9d6293e8e2c9b263e876bd29957c802dde8812508b5a51c1a54b12ae02d9fefe63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fab570eb35751ca9014d24edaa2836027579db3f7d72b69f3b587d6241d132fbfce208166c42d5a0a17e13552460f909f5c1f07b8f9d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa5dfc9ad48053a8fb1df7d536a0843572468e1a3e4d06269d3ff04f2e086ac25a14086cccc0ed45114f4d6703bd67a2f9b0f8ca1e60f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d013938e3dc1e35a282498bdc5f8b3062869f7b0c04a03198cda0b4530356752a2ef31de9cc126c5a25de202ccc3a4cce49e465bd387;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e6e4cd2d5200b0f687d1677607dfb66ed2305a9f59a844a93874126be1ea7c14dabc33fe695c6fd6904e9b43da2b3ce75c1e853ae1951;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h770df2f5280e9413be953a8f25e809e9d56c7397c726ed810d30449c488e58d4ced2c4c9e7cc7e7031eba9b395353768e9b186176aafe2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12efbe8e8a31a9a4fcdee633869a3aed84a8b31361ec5107bd7a945521c5704c0e3871dc4f032de1c91bada5895187633304279157f6c8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h439381999077db84df3c1fbb0d7bb635d34b25d858becad5dab8ce8a6fa3e7431e24bd3084028420cc750a54c4c807a8c25e9617193bb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habe0f483c4cbf22b5a4b05a83e415c93a3eca79703b9d59ec3174808612f8733ee1751447610367e90cfb810d7036390daf40dc0a35ac6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16681485b272051170d902374d175f5687609e072353dda868ebd93fbaedd855622d6a30960e2eee751c0b28397a022f1488f77777e663c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110d5d0a7214f7aefb280b92af384c2ee143d027a941bd2e5dc0f24edf236a2977606a55babff41bc3ff4bcfd056e4702b909c3241ece76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bc9e7783d0b6b6f7cf51b3f5a278a8e8d1ccf400fd7818b589392109eeb16f56ffd0215ce4fa0211b689524d24087a58cbd44903c8720;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f61767bf964bc311e8712bc661b7d155c740de9ea5a2de7cb054c3e1b086294a2517b086c649c531bf4758719be7a777274c2b69101f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97b7e77c9fc60edc95a4e98809e9fd00bfb0f26edabd1ef612f384a7f3d5f6e49d3c57df4c02279792c51287bf2bf5e46c9af0623fc3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he37fc858f3d7eaf6b4aa9de5cfac0ee701514d18801ec70b17325be5b27c8f9ba6b330a5e28ea27e8948f117dddc99763470c204d0ab5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed71e39626192147d0b1000dc2160316647c84b6184a01afaee1c6514a172d1354dd634b0a0d93e0f10abdb5c794a627b623d466409ef4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131fa9ca42b4d989de6462b563c7fc5057deb78fd907c00a3dc984821d724d993e00f1d91f4d1569d3792e0f13a638e74b2de12b4c8eae2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b6773a1ce3792985352ace741df8fe0da8f514e23ae4217dd981612c8b46b59bec1ff20cc9406746421a5f3c8d057f1ae58cbf6dca1a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c406322c3f5006c56bce2ce3031b313a7ebb6d44a5f4ed1eaae0aa2b71e71689f7d6ede64eea1f98bc56bd4514bd754f3d7ae279e79c6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc83945ce4aee94803debad4e8e2612a12eed495332b0c84574f36db3135eeab7f07605b4e095e1c667b4939656b160262ddffd6d88f96b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h206a36646fe56be40be71e83b3e37311f8c7ba6f8320e612c1fc2b2be293efcc41e7a4667ac977446504cdf6bd176057c6b07cf4d8b60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fadc0300e901cbc8ba71987a3f76e91115beda4734861108eb9b1e21930ca0d06f761c53ea3d9749409b68deb90974a69cd279ff2a15f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166f2376c1f5dc4b796dc2c31dd2175e347d9fda2df056365cc60d93d2b87892b55b9c3f5846e53f787a011aad5e8fcaa738536ac4c186f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e96b780f316a93c60041984eb22fd2d10b2e0ac6c86d2be521596f326cca9f9d6d68bd1bff9ea2f18f9cca9e88e94818541eb53ef3f32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17dde799f73615eb0d28f6e6be0107012d9be5dfdbde3a1188e5949890daea546c872410af0646440847e5fa79f3c4732b49bb6a4f5d8ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cecdf49c91f9efa8e77d19dfe5198755e5d65077170c11b012cd5855b7f3afadaa3ed77d12ea3d77f93281d72386368ad3ebfaf600015;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142db461a1913be0d0972d6577299019bb45af3486fc74469afe1dab446e44ed6824a795e9b6ae621a8a9d1457d66f86734a055b68b6115;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4fd01882a5c2e4f8a394e50f3542fcd5b988b997a5919d0d5db50f926b57ebdb065b1bd9bc4c94741c0d6721ebc1729db005f5f219940;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128761d12ee25ad0e08c25dcb92a96bee6dd61dd48d414cd3614949ee0509363f1920e771d1fe069351e56e0773c2e8d757269642dbc826;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf728854f4f2ecd491548443f3a657f1a2bb0d399c977c1ce7f7e46f37c7669c9f730dc2435be17d0c82fdb03aaa22018d9cc63bb09f327;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d79c8f400ee333b7570041adb7f16045b95f16eaea92d657691da1685244370745d6e2c74ba6a3ab5aecf79bf91c2be11f68722d8fde9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7130ab904245919011fd9343f35b4f1a044b4d0b03800ada567a85f94b0ce81a75416a15e4ac8133a13c6f8d514d98a50a1400050a2814;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfabead4dd0bbe35d105b1595cab1ae736a5719d73551a830c7664ee41a616860785204a91c5128618ee51ef6ecddc0cdfa64cdf3cccc9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd361a34604f6105229e205623be6b1713eb797e3dd9832fb16ce8fe9141f4bb8e785e0090ce26821f0559393ffd88765a6ac5a5ec5e3df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heaeeeadf20008fe8f1ee8a7ecc3c33205d06b2453fe8d5628e455f5b6a308da5c65db9824e5de1f1df940051718ab19f7d26a59fa45c4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4a4020c868ef5efcc04bcf41e7dcd8e44c35e7e5020b9380c563dd251b044faff5a591643c57ab73e476f2894fa7c615c3927c55c48df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h467fee564b23ae7cc505b9727893a5acb44ffb7bcb4a70d0545ac44dc6f72cab2f1f0097610600392ece0cc04da837b7f3bac7fe033117;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7a5a70987ad1e7478ad7f35305aee76896285916c0c19154c7ca5e62e437c8ab02f9d5deb2db96a0c427082db5c416a290a59888c3521;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcecc91a7838843d9ce14aa70960316b069bd9aea09b1179ebdba05511524afc4db664bf039079a6a4b46d4ab91f10af5ab5fb2740a85de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b0244fca47c85e8138e88349c6708bc704832961196280b9861dfa304a020fbe055f531f299db7e9d233300be1ed79e13d3f98a23f676;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f68d9ab5b79b63a2eab2c25c94f42ddd6b0f8d024349905eee5362e4c12b8d5a57c101d86701d564fce8dee1deb2ba4b3cc27047289da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144ed10ad5cd0c812cdabb25bb94c3c1dafcd12e66b9279f6a6cc351e9a57249f4b2d9e6b2fcbea0489f3d7a20500eabca5f5bddb6c36dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1714a120f854b5f5ec4be235c4db23b8d190688514cae7e5b8a8aac5b333dfe7791a21c761e19d41c1e0385800320fd0d0473beac00457b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b33ad7f91aa9b941dafa4efc13001ecfa622cc8dce55def5474bf3e9123ed8f359c618428103ef20bec4ff2e88d0d8b44dffebfb792626;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138eea59191f040fff97077e91481aebf9576a02e2eb05aeb060dbb973c6b0ca988f7eb8347d8599a939369c2de230404f122a7a9d033f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4948cbc6493a9abb7c009e36dfd0fd488c478ee016f465a2853d634037c07b324dde73890827b265df3ba419d62303776a1cf3c472a92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d51a46a2834e69f8ff1568ac5f3707a464714ba9c2fb62d4e0f0313d33a9994713215263464e299788a5a997adbf11a89d5f0af7cfb7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce68988e14754ad6b8ec863c5a870f4f3728b80d7e0c1f21721cd91e385f6d954e64a5d5667c37be1f794ab800248741481c7b7511840e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4d1276ab5cc0220f64fe0f61a5d32779f50ee664478d79eec6720c9713487f640762e9cb1e75a3e0b6493bea04a3e5860eb23562ea70b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94a812c69987c7659b4edc79e332f0d9cddfa63a74b117f0d4801b6969da975d87871355ebe685e285d12ba3e843b48e876bb98cd86b72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141bdba0194aa594ab64c7030d099889b9417275c95311e9cd6d484d76df1d59877a8c315100445dee68c327a9f8edba09e36b53e28a1f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec328e0d0a30243a33c5a1127b98b69cd2e951cac9ba4f18edd1913d2afbf660c6ae09167621fe0ddc9e2bc7ced37f2d30a4a1458b59c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a61020fe7e0977a8250b0e7b796cee8c2881b36e3c2efa437fd834912cdf2288b6ca7fefa7f8a751595cd07673475dfeb1116d44cf03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c490e5e0eae8ed09cc12c29f4061728d111ebe1bb245920317cd6d8b119ecc4b9bc57824b6d97d2c40c78a1b4a00c31c5fa53177f6b014;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb34f511d481c7ffa5ab1a583e05a1d3ac69352d0a14a1e67dec6763018e8322b5bd119d3aebb6372f2fbf3865d6bbca2501293f0fc822f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fee6db6799a157862e77fae6ac21d6a3342858fe80b6e5d8cf1e3ec9d5d0f858d39d90cd782af39dfe6aed45ac40463cf45cbc81cc8269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d99a627a1b96e599fc1d236470444a0c1e9f66873c21b3075ccfe68ae926b8f5696786375d32fa14fc0d99ad4d9b2b1c34a1bec34c6b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15970c992e0a394cac0b61a270dcdf27f74dc145a4dfa700ac895067ce88654027456e1204a4e07185671399a76a891b7b8d8bea57604a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116711dc756e004dfb7155cdaf55de24babd127ecd7951484982d79e663709083b4afdaffc9c243f7b369a45d31d4bbcb5fd4a23a412040;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fe653aa1c6c0f00e7ead29ea7e3dd23a1784f5143eebf785d8887382a90c1e10074c10242ac8a331a001869d6a4908fffd95a78f71ea9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c31b8b8948a9825d60c295f0a25982db05c6b8bbe087eb37043bea20ee8a5385b078c404223f76cebcd43ebbbb5d71682483e759aaba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163ffa83129293eff59f5b9e261f4b474404b51341c38176e6939fba8ed4afd37e5449df97a0770615800e1fb0b45fa17f6323a7a6d4184;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13173ae9b890139c32ba0d169ca788eafbfd068d13792171a8378370202d99681e414b03d024f4887f090ac9deab58bf227e2e772d567b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e34e97a5f067685d0c17a2ab19edb709d27d33871631a96d00d09c892356a96bbc493f85db70e13bee6363031904db537bd491b8e956d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52433bbd50e48a0b307487769bf4e1fb090b26b3a6d58d8a923a0d432d040fb29af6634cf99b5fae49e3171e2a396aa48a4113b0d204e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97bb4cfbea5d4bdabb9887c68b53a281124874490eac7a576c5c54f5da70c9ae804527889a7171d91d0dc34545fd8a54fae64f3fe4778;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h777ff7e975c1055a3e96c7e2079b2a37c17f2d8b58a9367efb4b10e85f3c3884e4662b96af0f36299ca639140e6ee93b81f29299193aa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c38fba0c7047ce0f79bc8bed01324a8ef313cd31570ffcc30af9e840f11152ad91969cbc960d7894acce181895ea9a109d29d820628022;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1add756b0a07b0741dafdd9b07b553def647d2fd1e1a9eab9419f881fe47a6285c71ebc19059af7a342ddd1596a2ce636f3a5d29c8fcac0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e4b0cdb099575ae84dcd4d34a85386af25172f1b21f29092cda6cd9044652b6052db2a3d91f8c7bfc9ba5014103d9bbbedef647445d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0fb3c11ab633c62235e77c8f31142a5f9101ab6b03641342e336d3c8b37e74d885ed6325da4e01b678120ec1bf8375bd7d0abc79b3942;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123f299b0fab8bd634747ca7e9f83793b454d27d884d8d8c564219ceaf36df47c2472ff8eaf52072618959cc62c8811c5212c0c1ccb0d5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0a6803b716bfe8f09f5b1c70617cb487b147084ae20a9e5d61a959f908b4251a2f1f7eed8b59db0376933b34bfab2e335c758e8b0f9ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e52e002a2c01c93f9cd63556bca59b4e15f7383de4e4c51ba244617a871e900204a5347a96ebb8be107fe33a1761c924eedc595533011;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d346436ddd8f6e25bc292cd3787a303db26a2c138a6ba9a22382accd0722fcd826b86fb235f417a30313f24a3c3056d6f4a0320961188b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbf16d5f1c0eeb8cc4a7ad90970bb0d9e8deacc0a776cb40ce975b9fb6fc99792664c6dd4913ea43103b334bb66b72631b852ab1471051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57ac30158f9310ba9c2affbdd9cd5da225f0c1de53e05a751d302e35989c7ca53659dee63936db2f77b077bb922b5d0b5e7a3c218341e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he718995d66753b395769900ad7ab57a5b236e1e0d97858ea249c4abb532b2ccf2e132849be05486fd747e161d6bf31557e57eca0af0542;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2e37164597420824a532d238f8e2630fa42e074853469f762806bcfe9b81f7c21502969c2499be810dc2d527afa6456a6d8fc0020dc95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8fc91c781851ee68a89d13f6b86cd7c49a03bdf1308321229ebe43710962e37ceb8d1bbb4e59d4acb1659a9d809b71f6e13f484c74eaee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h440568255cbdc3b4bd0fa4204839b60e3ebc865b01d76e5fbc7b64a1c04c3e67fc665af64236f7ef1a1ffdfecc730831a0fb51caa30d67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a126b470d5e862493f29a068f6409f23bb92ddfe25c596ded3408ad5544babcfbbba9e85c4b50b8221f4d0b7b50370cbefeac56a04dee4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3f45ffe43f5b2940baef9af260ec4b366498ccd7787dc5bbf364dc73198d173867acd5890b736a42dd467f8a6343915946fc229b76933;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4e339369f9baec8450fd7a751b01f7d6748d6454a6b26c9f34faccce107d1789fd97d1b3a092bc63416a318e5f467ba996a2cbb0c90b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8d6d6ffdb5bdacdc2c00da4295179f646cc6202412237922d5938bd5190e772c39ce8fea03cb239d396446978261f15af75c5da86f9aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e22aea8013f64c2d12341b10daab02432f6adebabdf0fbdaf14d5e9f051e60ff9257f75e20273dd0e06ee5a8002b7bd4d5936d75e73be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h766bcefc2aa04309270b382be88128afbfb7da622666901c1f7f25bf67a4cbd1c0adf5f3ffa735736be664dad46d24ee1e7c232be02714;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7d3661fba853a5d6637a4bef6ac4c6039c134fce2a15477f736b48707218c6b952660e9fbbdddaa20dd2d196eee9963daa165b2fb4c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb67f6b9ccf18f57be217437de3af29e0971581817ee65440d6e8f200d8049f5ebb1bf4a73e104f70c56e2f175803f054aa13a5dbc4c8de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h493bfcdf23b713d957cc7fc9a81268dee4046d8cca86e328b0cbda16dd62b999753c635466fa6556eaa7b49ce1ee0830d73de5a6b222bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10dc407af3f3f8cf94266c94c2c4c2dfcd859086a2bc307996021d0bf62f3e9ef40dec71217a39885688780d3b0024e6e31bcdd403414e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104a368b15de1ec65e5184747651df67878381d6b95bf74e9555bd88fb0ce92385e03d75fa5743bd341e7fd35f13968908d6569d8625d6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9273ab82eec541c035a90756694febba38d3b1ff930e0c47b777dd7514c10eaff9ac3dc96844f6d94d3041f873d75096c350851e0385b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d056b773a89ed863145f7965a0ea35769e7ef2fd701e2e033411e8bea1f75712e9d37b80f3255daebc772bd064cea2ca4e1d3d61df2f9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f37e25d1bd0f5a6dcfcca20f59c893c617fad67030fb879493bce7cb4e352fe9ee8d8f32f0eb1ed977cbaea4b4fac8ce26f0a2275f47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe6574d876d0f558a72b50ec8ac652d4306d4571bd754ca2fef9fa6d7ad78096b140efc8d4e1c96605580ca68e7990293c442c91679241;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdff5b7fcf29e52de19c24b1d234109f8593fed0d4472c349dc0d4099aff6ac7410dc36c9167ab293e6409067d889cf723812d6f6dabbd2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8a1a29590252120bd15870e94f0891944ba6dbfdc6cde20345519cba892b9b9038737f7d036d80b960078fe8ebc54bf535a3309677bec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd755f9e2b727dba0571fd3a26295f812497b0f31dbf41579070cf1cc5863776c1b85332549be532a0caea4da5f08cd326cf7d5958f49f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf9d6dc826261617c24abedf35cf97523cc51ec41248dead623d3c333e7767113fdc05fe8635c36214269744bad66ad03c0912fcbf6023;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1942944f3d33f69cbeae9c24dbac43c51f88360812b9d6936ed94e040796dba2823d91e88d3e67610ceb5851521ca1e5cc648480a7f6d39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12abe9233a9dff810a27787dd296cebc832ae6297009d7d275910e49f7ce6ae31fda5a61916ac96b20a0590283d15ecf73e44b632d8b483;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d2f35241fa4fef7c150ac298d6fbe3e8ae7f00bfad1705273eee7a9ffbb7fdcd10bc6916e453f4d9f903e67a8afea77d474cfabb4c1da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a0c31cea677c600be3e0b59af47a9e644148821dada52e546696f246010a4a8e8469435984e7cb20f966620dfc1d049a892496426bfa1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107a76c71504d3cb81ed141b00cf4728ac9e03d102a32f67ed651c68fa62df62a255c01ebe8cee9a29ba479cf748db55faabc4f810d2d43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h586a28a5b112d6abe99887f0e82569dc1697292c3516aabaff136c11e3094fb3fc63966da40b81f83e4519b0afc923ca5571199f647dc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39aa9a23a66f0a23460dbcf439f76c4fb9a52eff9977a86005adcfba69f790a18bbf5e2660aae839b4b75a1a9143f32273d0197e37857b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a254249dc422900602689bd5b9f7600386fbfce665194554d28de74f05bb013aab6588747fb211fc9c6b61119495113da9f86f8cd80c56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ef602b181710c8fba3a84730bcb0d085ed80c4a4f069ce7b412f8050c3e1faf32455f3c7c2d12c0bacdd137234e1b825577f8f4a21ffd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184c1caa4a51b4553ca6f65652bf5d6b23a3ba8cc1b4cac31fd35450441c7cb87e460e9325a665d2f9a16ae5a997f7bfab5a46d3d72fed6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ea064d0460161d4d523f280f8a5ea7ee6e2098f88b833627c45423814d7986df239bb569206a9cbe2fbd10dd912301f8a1cb49d7a0588;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c128ba7e3940f1815b78239f2087a49f6f8f3d38626566c89630b80ad6172724e71a2d864b226ce45dd8fd2d65654a51cee9545a1c540e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ae7434bd0ad2085d1fe2395e43ea79e5b950606ac0869daf35f2acc9c858b4e09857bb29c9c53bc22bb482596ff9a03258d0a5c0165fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1711cdeea53c80d90bb3844427fc4b7a615611d05a434b94047fab32fafbff9f230a40a788722d49e68d17fc39fcffe9be2c925279ec79c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71381ad011bd9914d2f35c3e0a339d59a071886d10b5e3b5512479ff7157c729d8c380d5c59ad638f3fb810e7b3f7b8af9d9c7a25b41f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9730907599a93076ec627c74bcbe74cf13eb862b6ea1632931c00cccecafb0597ab3b60b6a735669ddaaf6c8585315b75c2813083acdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2afee93a37e6c85c31fc1afb78d366e4a8c5612ed86c04cb350e907a610784e2e14389af5bf9f93a123dbfae354c3ccd734678697118f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a06c233a30ba03be3240063d7cb6b3bc2ba392b1fa9d4b0532f7b785b824e13e4909e752aaa66697a8673a44bd410bd4deec42e34953c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb27fdeb252e3eaf331ef5ed4390e180c8bb98d922011a2fcfb29313091a8579e7ef456f2724f654b50748c4102851048797b52c52b389c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7afdaa7880405a6e31b534028464d8ef9ed650aa866c3b71e2bd43b1d22f4d700da757a612977066c4e01943aa9e8789530ab0d2cf721;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9f0c255a0c9117c4dec214d8e75b7fbf0f9cdfc4a02f560c24a32b936d779115ea42087703c4184d71f10e8d7c2012ea5f89aa4403cba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1238cb3867b4ddbbca814ec9cdefa27b84e17d47b2476998181bb93b1b13791a3862924c506a833435ad33762e45d7ebfb309481bc56d3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1025ec664b6b6a1bcacd7ff4bde46983ea0aa11921da7c5e5bc9114f5cf5593060b1866662cba74bccefc64da959a26c466213aaa0ffa8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84f61724d6c7ae60fbfa0f223f05ac3bfb7adeb817d189ebc164cd28446e6fb97ccec440e440e60add2df963613495cdc3f30a1909b3c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12509df8b1207f561af424351d76ca7ea5a5954ee270f55d8d286eb8b600b4b10649e0e8e6640e277cf36c34bcb404e2bffcab6ce407b3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53204468b55fa98d77e329ebbc9636bec4ef8d334a06d2ad610c48942cb30271773d830dd2ac2aac193dce5b31d55a4209d617c0cf7d0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38de9f4ea62866a4eb8ca969096cdc88d654c6b15cad5159be84579cf3a259a4bab9d3abed5b8e82ec2d758856cc47c1b6e34533c90c75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ad3b6abaad1c26243155e35de9b29fa4c601cacf555553f17a5523e539a58ef1dc6eaf57e943d10705fdf9d2e1f037672d9beda311d98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1009192275c9901353037ec440b11f70d856866ffc1199e26722dbacb38221fc766af4f642a2e2574aa04dd8429c6e21b03621d02a6032d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c3a630ae139506fbc4575bea863112426ad8070e78cadd55f6572962677817512ae7d144442efab1d5929cdccacedffbef08d006086e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a128e3727ab39be7d1905706db728e0b7a9d28160a89db6706182193252c0c9b91dbccf48aace4178d11817e468eda4681a367691730a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb549e050492f5d2309ea4b7aa0bf7ad144ce162e47b0ee6ad29dc67efbf5ce9d2c0c9c6984d9b03daa9c02b145cdb20529ac5e8c72a58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba2e070459a20f87131d4de47a72bb98c1af3fba273316e5ad6cf52e0a47868a3ef8de9cc04378ef4ed8908dca83277624306091cb5857;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102a8496965eba36bf9db34938c48caf5d2a48d515a2bd7ed27c0f54bff896e2c95b3132758aae9f33d58b0315d6f864cf3e4126ee2c585;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1498d0b31bdcd9769a33732893b4fbabe278fa09b05634b9aa1c5dce3a8b14c1f6472ac39b9f69563c32af8534fc84c974cb6c410a50de9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfba5d664f5d3fce00017c9204fc5ec7037a3f3d3e8b1f3781474676bb64e435203db2da7030ee11bbe32365b22ac537646f97a59c573c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a0c2d35720c0af9d3c20d53515bcb237c9013bef6031482d55c628364a2df99a899c798b5a979b44a48c3bad74f51050b75bba9e07c55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaddfec66254d3f2246399d298e78c4970e14c4123047bb19f76dd637c2fba9f4947aa99655e86f7f1892db84949319961f958474f9131;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1184da794e3ee2b5e515de7cf81118a8a67e7499fd61ddf2acb29c2a9a12907dd613c51a61084f17cbc8e386cd8996a2f9a933d7805303a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1747d975b0c92da66025f80770ef05955c95fbf92a1211d3c03ae2bf9174b086407ca1b16d1dea570fa4deeb4cfd20a5a2c28f0744a7269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e07653bc8113ea642d944280c61781f99776a46f7a7f881db5def44d11bb89211b9fd5867e05db8217b5ee29590838e094c9f36d032dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1baa60e60382491b148041b96873bc3f9551a0bca618bbae9026fdae2cec27ba28734dbf606e081e665a7eba2bb2b0e0d3da0a0c4555a18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h460235e175f58f789a1022beceafdc997c5ee34dc52614cee9a914146f6a230f7f453a3f42c83b926fe2f1ce6b3820cdeeab0a20e178af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ec43c8c31b4fd3e63977da3fdc0846f1148b65508239d8cf8677c6f7dc83f420faa6aeb72cc9eec5aa3050bbf5b5dac7badd52585d8f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df7c52b574dbdbbc325a73c599dce7569ddcbbf7b0bee2cf3b1d57b3bdbf0b404dd7541e9b1cbfd9891828869623fd04c602a68cd36269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ed4500a66d73d5f5916dece6fd99540877dc2f432eca5fa2e71a10638a84cd4eab967ae17860476e36bfabbef1511362868c8e7480b96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1e09ff70d6f1747b3ed3907ba9d7378485b588acb6b3e932e331c160ba0934e8521ebefc3cc90acd4d265438ae44057a3c1b0d2fea48e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f2f1b2ea81162eff75fd3ab1588497b137d851b4cd6b1bec0e02b0ec402e93755106e7d2ae1c69e8913117367863be750644cdd2e73a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb301f243a85703de9fb22a3871b8fd6af3015a9c6cd9489a6b691d3a9a99d0c8ba03660e2f2fd6f3a648070aab1499dc8a3d26013cf32f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12817f0ee60a8de9e4cf087fb9a0851f61aa9aded8a6be8e999617eb46fc07034f32e813d54903c4e614d9bcde827bea9fdf68884a1cf0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h393fa8cd3a62009f500a8f821d1865f2e5ca4436c4c00d59ca2cb793e3a54e1180cef630072997a8d537881a527f680f4230133e1a6057;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4dc6464a682f5ad323570542fc4e3ff4d9ba6a8b39178f8735697ab96697598610fd4b96352619851b86f5c33e445a359eb275de62e02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd5f3de0b63e3576a3cde860b1d4eb5af89a9821ae95e6925bfcd9c6c238d7d69043f58e448eb05849fbbfd4287972720e7fe2422ff618;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1044ad18766d05b5f21484ef02586fa652469a001f64fd11250621a3950b3465f5d049c431ca773890a1bce16fa9af0cdafa34e57ac47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71608e5cdf73f71aa289729ce7bcbb67177cc711c136b3d3b98d10628705c4bc47c6d8b1711f2e402ffdd3092e54813380340e72779cc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149141105dcadaeeb2fc3d56eee92e7bc2773764427fd1d3197a2380cb7e9ff371ac35506e96a2f6a21e6a9e05a915419b3f9a5ed748965;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54715624aa33036eab3ca5aa8fe459189c621581f2a63a40dbaca1bea0ce1c3c6f646afafdeb7a35f9aa9b16bedbc8f5eb1f9dc9bde5b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc208208491d26b4b5ef21cf2726f8a9978df2b9a5787f816e9b11a85daf9571bbbf91fb3e7f8642ba8f5c4947b748bccb2bbc41d36e5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49706de42d096a9a0975ea2bfce7ce288914ba402b5e54c93576eb3130b83246559d58b3884e6b1ecb6aa1f8af591846a709c0878334b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196af49def02ec979404859fa3dc749e761bc9a6bffba1857d8871f7811d178dcda04ed2c65813bb173e1fe3651f9ee80b4d3030e43e96a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d822fc551add4a2640ba58e8f72c8960839e39448c9264d82b0d8501f2cf801ad5d1a4175dbce27932c3d281ac72029311c14a485e771;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb05ece9849226ea5b9baf70954b1bc63cdcd9b8f9c842882ced5a39468cce7dc2a96e091b7e7eb8b8c729c25ad7f409552374c67687df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c921ae5d2b71031f674a0604c72b4f509452fc73ced2ae7ed2757ba1347a800b3661f4e175903a3ba68b775465abba1bf97ae0f079ecb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a49d7d313e486df59c20e43ad3a7da9d0581185bb706b89219108ab9861ec4a4259d0c511039f0511f6377152130991b732034526bc0bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c7041a1a0a9add9e65bb52c60a89352ef5eda2c7732ccc64a18acc283b805c719d1a2868cf096713ae634aad1d858903d8c7a2f84f29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69a8a48328f5e0d2d970d1b2c2692b886ea4befae410fcb3daa10de6d0dc178ed88d7be53a41f9b790458586bc5cadbcb8bd0190dfe0e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h257c7a4f5f171e801bb5ecc460daf6fca55e33e2988ff748d6f2c825c1579335bcef165eab8abdb65c5661b0d82be61f099e112a301716;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1056d6daf96289aed32759b4965859b3997b50834dfc010d9b023a354afd5dbfd679e92858c3da733f4c85147bfea468b3d53ba03424e52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98fdbb7e82ceb8c623129c20f41e32138a06cceae77f72e7bb2f70e7a117299e1ab341412542def079c17fbd6112ffd506cc040e2f4d99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb26432bcde977f5c2254e7aeff6e0d67cec7c183ff85fe0e9ab441a50c0c77f61d55153bdbec2e074d5b04f5b354765ff1e682759bb2f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a945a029629ec5f836a934ac04fc64cccd13950adb22e985ed39d8d061ae6c9e847b212fe77980bfb8f2f19159c23c7f2357393ce25e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1014482ff7a908309ab44e8843f8e18c40ff44703360e1502be734c70656e7c7a173ce8e2389f616c5d26278b442b583326fa4a4054a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfb838ca39f7fba957c74c7f03c81f236ca9a3e88dc539a99ebd12edaacc629cbd268456d8832167c039f0faaa7405079c6e52fc662be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103d4e8d869e1c0d8d371ef24e43f94a6067343e160a0ccc8aa2f684e86a68dcd1fb6f7a88e809d7c0e7a914ac7a05a5c10c0bea860f597;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afeeafe800538a0d70c7b059900ec3ae57fe0359eabca3bc09d93ef12b543c2254b91db1ec3337816e183e8c83ac19096420d31b6f715f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h697546f89939555bb1450b64d38ad87447680cc8f786b96c93628ca58ecb6c01d733695001c201fd1a0df6f4b3fb38d375c14207f6e3ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78d84c7d0c96edb096c70ca7a06562d176426cae366e6c36136f4e8dee32d08f074e2a991fe72e5ec711bed8604589b5720adc684cc054;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc920dc1905940357f41de46b7be5130439662a44a7f1e4f53aee9dd2877bfe24c3e3d46ae6139c93f7961e7983afba2da924084d53cb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14971f3f624d7672d67466e1ef7defa2709014dbf0460249519c26d9a64e80a6cbc6538f16352b9b8cf797b0c80b780615a02128f97f68a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137afb8a3c2e256a3eec2718389c7f704cac5cfea7b57da1b05b7846afbc954d2e87cc06e6184b14e33280d90091136b874514d064004c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd2063012e0539280ce6dfbc027559dcfdfd4f33c689d56458abcdff8a6210fe72dca08dea673ba896650ebabc5f8a6ff83688b02efb03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c0655efa546389c0493a579a6c65d51904d6c167125564b29154b4cff8f5beda53a08bdbbbe65f8224c6dbe45fd089b71e9bac3668b7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a708f87bf546e57ccbfab9c7266d12e6672071b3514f42f1d1c110e307d4c865800e3bc2add71ca08c46d6ec80dca29758d7d06a54090;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125eab0f3732ddeb184d09705897164cc690764ba9ddd2333d8e3f0ccb892e9197ddd9f26e289b6cd2c4f7a440b0073550e4bcda51df270;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cde2bd7b4cc2341f740d6a20b0985f55950347f824a811f60445fba1613f9d87bb105c666644686b65650ca8b465c918adcf6518b0c26e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e37ee1f16c21843dfce0c713a93a364148a52d8184598162268722024ad2cc2aa4df0aba750abbce73bf839bc3657afea30a4f8d05e676;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129751c9996a6258e0b9788a63475fb2e962f8ce8defcba72ea1bdeb4bac9fc53dbcf73aeb836fea5c4be0bc48e5392b32cd255ba281528;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63bec21a0b9e1795ce5c336fd0cdc17e5cbbaa20251599d8b500781c5403d57e6c892e807fa1a8db9550ce480d12d3d26eae94c2546629;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de63c06a9048e13f6421b6b1860b884fd239eef4279355ec8c152f7c239d9fdcc60274d83c4d4861b4b419ce75551ba94a65573fc0ac76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a6a3ddf86dcc06c6ab1b8146bb7d96bb3431312f8fcda77191da18ee13b77edddae835a3bbed4ad8249fb2b46fdfbecc9c4e1a2657c32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c1e5adbd55bf5ba07dd71fbe4ec76b559aa3f41b4e94d4a5382e0cd16affa4182a82756f7acd12aff6ae92fec896ac7a41e72447de060;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bff13a61b064282e113dfbea496eb6c01217153b335298df9a47bae0910fdfeb651e425223578a64b21456da31199771a1ccfc5057740;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h258e509af86fa4437ff1c7b4d594c687ea7176c31cd724016d84343e8c40dadddd57188713e4f17524681813422443323e577a7f063fdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18585959f6d81c4a06740a4dd40b66617f8c375eafb4e642083ff696d7af5213170c9e85d1662f5b45d9e33448c9898b87aed3231a2a768;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8a9afb228093ccde58ff53bf729fd78d2e92edcb692f87d2f89a7eafd5402d5365a4b3337eda08f2ecc3b0ac636361075db3a42ed52ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c19f0d7d6403447332911df5024f5ef543b04769a38c8622c25b06c6329a5cba06ddcc3e8ed3fb4a84bcc5cbc6f7304f23bcd74c78fe95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cce232fa64327bb2611d828bfa89fb350d33cfcd353853f5a0967951aec65d3fd69d7b79da599db9cb759c647c08b077f5b7f06b5b466a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135751137a083464503f66952fd64da21f272c92afad8bf52a8e8ae15b9c501507936640d1cf73afd336eb37c43179aae62c69c1ce9c154;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1980215f6e6abba90de63cc2c0d01d53ab8f00c376649255ce18aeee8983afdc0bc5052696a21ce4b35fbaaf1a17ce734379b4f24ec2e1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf786cde2afd4f738dfb36d8f58edc181347fb51f5d77d17d5fa56514f903e2de5174a6d9015ddd196b4177dfe6c658f3219c33a77143ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h924d3610cbe9e3b7b52708f74f85d28e32ea28b8105d20b2828bf33f613a642b8296bc5c706e3b5021fca2a2ae8405f24e65c343ee1ed1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b9dd2c270de6dab3b5715450693705601c55396a6904b4bd92c44587df9c0c20ac445ebf87509076f9c2d388adc5300e0a3ed71510d59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcccd4c14a2f955a381c5fa9ee772832d3ac80ad1a5ce96334cd022cf8dc04d96bb075d074d7cd26373991fb06b00ee79d1f307d45548e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4fd0067e127e16f6cefeadb7cf970b22fdbae5eba9b41e6b89257f1b3b8e1278768a3ee7f73a2b27781a80a520a016b42bf08b9cffe52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fd298f0b323b044b8688874255cb26fdf97333664ff79edf20e36f8d4b78afa3aec9cf46179255afd08dcad9de491244b44f3b2dfba5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1793a0b47171c7249a6e2c302cd9284c36535943551c65dfb5648046c97731a9bbe59d6a1b7cdf2b85a49c898ba35fa025a4378a0aaecc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c15659ca966852217d23297b9ff728b8cc7aae29d92fa4ab7f55a6521f20361e98056b68d37ac2df8c456681b4f1b6e56315d5336d9e7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30263df623945f8b93f2389e6ab69cb4b4eb97e65d56bd7a457f5b9741ae95146b913790dab4b9e20e14469ca3c8bc26694087538d72d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he70a3ba38614e6ef12c44993e4c87507ff9d85729c636e6024df643fb9e46a29e3c5d901900b2941331da9e880b8d584fb698a578af1fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54ca31f086c8d37e220459d7c45e469b253622003dcd5eb2238c3d0f4e11064baaecffef5acebf68fb77d190a7c01bb6d53011a292c5cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb59b192de57cbc88554d84ef43809e82f557c4d94421cd0381cb4a8040736b8f88a2e613d4d52d2f7bf852b446fc9b41907bc0a0506f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180fc5edc1de4aa192627e3e70b90b5e55eaf8c9442ea6fb5716a3787c556e40a6af8f9d400dc6a29e6b27f6a41dde3cbfaeba2a67f23eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbec9ac8f0740ab0975dabfb05001089bfd21c8ae1dc83574419dbc832bfe27290dd37073cb2a14d5df44e25003d4cf832eb5b1260b0430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18954e5b32f48cef3dcb0c0a0d3be3c82ca3fcc822903f770e9dcd23c2ee737ae0057c5cd0221d0c0c5fd73c6b4808f47f37592d6712c18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc14eb26207239adca401a9947a285fed0bd2733e5e3e18886e57b2a3212218bf415f7919c888a45bee535b3e77315cd8cc1f72faf4f0f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8661152e8324fb9f5a2c0b7663266225593751168e50e8eacc9b93a89b4e8d056cc5ce0b6138aa41d0acf5868be527ebe1d1da67de0e8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1496777ecb9a1e5b6f54766dec456620abe901761325416a8711cb135659c2786d022c3a697d67b635a8464d0558b0a4c29aa6d63e561e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he092c67b1335bacd586ae0099378e5e8b186612cfcc4075312555f0139a6b96e4aa8094f272eca17073d266ac3a164a806313301d92a79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb9a38610ceb423eb1afe57256928a28a9f5097c0a52a2b12ed44f30e86ccc9ea7ac3315d74e6fc386fe5b1131cd59e99c04b31d49f5e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fad640be0d4593907474623696f1e5c536e37a78dc5ecbee66f18082f9d7c536a4e2baf8afb660af8ce695b8a27e0c0c013a7c9640b633;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19663583e901df7ce88525257be2a0d2bcbd63468846f70a74da4bb6079cefe094a253d750c1109c2ab5accf448a14c29863c3796af0b52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1525e36332eb6db0ca93cae2f2cb4622b84f90e999dcc76c4645fc48a41d0cd98ae98bcbc48728177d7ad3c6659ffd6bf5a3ec2afd9c402;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87f96873e3313a4b76fc86a01a40081a8330b7fe3190eb74021fd6289f933ffc012065dee7ec96e7908c597f9b8c7396bfe09a5ff6c316;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52420c2587620c585133a91d140c1fc883ccab6f5b1d69f76459234a5637685e2e80e606857e2545ac12d479a8f7f52d3708470f5a3edf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a046d0fc25343d0d90d70d48bc7dd9ca51be535eadaf3e3a605ff303aefc5306b59da111d696f247d734a729704145108acea240c3112;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1100c90bf44a7aca8d9683e6ee03e9697562c373362d1505f4c916cf5803da9ba76f563b22e0f5abd119b6742390b1aa7bb2c85dc4612f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1379d7a117a400cf70b4b00af7f8acafc0cac1b5f0b8f1c016a911094bd748cbdffcb46ed9c5495e459d1d0d94f9ecd1f7de6f4b987d454;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e6915bd06a2660516403d1cd33d328773e5c5f8cbea38c4e1cb7905afc8447552acc9f6c9abc0b736e1033f11d92ae1699df881f63f2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191e32f63c12c439fb52fff53c2c1a0a59f0bfde226805bbcf2322782cf972c6d15be98ada5e83b6e00482f6d5d1b9be312c2663f4f8fa8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12086e8390e1c4dcca32f067321efcda46c892361615719b5b2991323a3af3f6e707368a722ae15d1b65378b0dc3f86c338a88c342e3bf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea65ba3f482698e07e0d4ded359ca797fe59d5f01a0a25fe938dffa1653e9d99b9596dcfba852d51194e7a3ca6c7a048dae41c16e49a9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b5561aa3a83dfd446e64344b3c66c48ca148bd2ed2e7f97ada42447521703f9878f6e60a3f77f80382c5123f2372dc5503bf9fa1a35f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5830305a3162b94fb72b23d3b600e0ba089438eafd82625a4fad0555453fe4febd0f7261efd3012ad2fa52a635fb671bee4e8a538132b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19da1c5e9e4f9fd88ef6f25232a1752cccf4c68e16ef097d1b268946eaa1e906227039bae1202dc3a6931d5d20b59c15e556032dc6264c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f5dcb8e54c39ff0f8a1c2e0975dedea4024132cf87ce5d1d12a2584de86a66cd050c7f8778f981ed7c9b4311dc9e1935a73ffc7a96e62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee2d62f8f50b75d90cc7ab507009bd656ebddf127c579d6feb9550635caa511a73010f6f60a177048c4d2abb721b5f65a1792f3c6e6055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b9e8827b5ad60ee7609345bdf7bcb0e2adf698816662def8b0d321b5a3cbfc7c5e89e8f2ab71002d36a6fe6a523b738712337ff98ebdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fdb40d6af6505ad557994053a779cd6b304d2109831caa1fd40aec38bc8e868667e18ba5e9ad842b75ecc5d65ec46147d2314faafa626;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h260a5ddaa2684994aa1797f61e970c2d0dd3daac7a2bb0744926c82da7cd72116e39ea946d30f3b78d655dd2b9d1c2714808f63f3011a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1162c8457449cf90edbd269076306142d107eef859eff64b7866ceade93f27a942dedab9fb58043a86d2d5ee717069d26a155767610a9e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf62ba04f7cc312e5ae425a545ed77b75066c5b6bb3249a078994ed1290ee90fef97d43038ff3ccc5f4fd0fb9c6d45e76caf7952101e247;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46510c9f89f20c545074afd0accd94f60d0cc638ee0ce091d39d94b816ba2b7e54beb86bf6a0bf097d7cab24779deb3302515b511c2bd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7af3fb01a5f7970e3a11a1ee0c879b50079e1c09ea532b1386c079d89e415c86e3529efc2251202cc960886bc0152f740521c994659909;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b29e5c41de0ac1a040eae9c83b1149f1c29f680dff785954e70bcffec3d57b3f90564ceda2dc5e46ba3102d442600372136525f3d8b63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d71aeac031e66346ef6257e512b3e407acb1a41b4a603026cfe81c25322cbbc4c56973d0957b39b90d1e8c71961a55f24d1fa4d6fd931;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4055c561fff56fc444ea499a64b03016aaf52a90e2e42718d86be3099548474c9dddafbf86be1c598846b8e459688e0913fdfc6fd73bfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d73bf3ed5dcd11a00a12749027539370d38038fe6da477ee77ce74393a99480d725eec34e84d435cd2383d16e38c17e76e8d3514c35c20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb26a6ea9e70fc1597a1ec2884af67eab93bc909f5ce08f171db7d38a4c7bee9c079ca48d1d026004bea23321e42ff739b9aac2607b294e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc8e644c00447a39cd27dca51f6e6e71f61df40ffdb9f95eb22913e833fc49107bddbfebd0ccdce242e598d9d1cd85c1cec8046eb64a86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha057ded7cd059ff341018e489192bf2760e9dfa5a57a137c301512229786c1094420424fd7bfd916a3a6a228a3b39b9228433117ef359e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e4ef448c97ed7b5988fc0f2894357b158971b0c9e9d6bc0f06c2d84f016ecaed367bb430679c9afaf7c1aed66dff94fde358c4ac7887f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139d2306bbc29ff8cf433a8e5b8c3b14c483e394a287c39b27cf00f31c96c64572468c3f822e57b8a41910146fc94d64c31ded2e75b789a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9d8df739417f3a9acd0877dc681c86d33660378cab6cf29da14eaf9f8e3457f1f0abde8fe4f8f82b3378fe0a869f33d150b945f97b67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1942720339f30c8a492f2d8ddb75559e3ae4ac7ad1f64630583cf9473d2082e35962f90af154cf506c5944f541648106c7a2b68f489ca74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102d8a6db99b6aa71751254bd8fe1a4a3f5799a61b662871cfaefa66b42532cd6de2d5d90c009f4d654e0d8ac1349d0637e997d434c0e67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6a2b6149225f42dcfe3df06abab813d7e306bbc1703a6bfcf8aaf56ac727137d55ad58fdccfef3701a412cef0cc327cf66954c6751997;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155c9e9174cf9a9d603efec643d0feb9d9ef21e2a5bb4785e3c39450a07f143fd1aba45a18370f86f27c05ec10d88e3919197de66bf1361;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a788f85f8dc1a9bd8a439e4082039942c6140a84fab1871d2ab5f99d21cfe611013c23cda04279a9695d9a11ed3f1290d0b1a214258ff7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18003a34e843c75b1e7f47ca138a9b04942a8e8d3fc280bfc1ac0d0b8aa94b4813cac045cb0fafb8221a65ae4467318d019357a480cc75c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e8ebc4654f0ee413411e099530826195378a7c81bd4e3bd8c422bf49ecc49d49d4db45f3c9c37e746efcc1e8afc56b31f94b4f402ce3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a50aa2dbc435a86ccc41a5abec32734ca10e34297ba31e27deea4210542afbd43ac65cd0fdd532086b99c9f18cd1f03d9973b75d6892c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f731477875897490d69b1ad9783297838454bcef3b0e0a20b50ba8cc502ecb0d3ec585ede252e7ff6a922183411794c350a875e07eb56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1340ec79dc3b2c07f64afbdf98322942230f184b48de0fdac4d65cb467ab748beb374104573f401013ec5c8d022d1ca21eb4e4d13370ea0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1959650e2e6500842af27e0f6f48216b2a492aed53692e33db6adefb0ec791744733331393fe711fa994ae5d3f3240d71dd88d83f3050fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e01bc0046e92f457b877ecbba58a05b2168f7c1084b4e8c95535a9859fff98d0e28d889535fa70f9e3f224e0363d21b19d6ccf26997616;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19886d2e047e134c14ab1f387f8472c29b8933689ef8aae6a7aee9462d78cd7a3a8b066c59d8bad355b85aa280aa54cf0c9498834c7e411;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h991b3e491e19e2bea5a7bf08bd8b257846a6596b83049f1e8a21dc7d5faccfc699943780d0c4e56bc99052289123110f77006b26c98609;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef67895a3ffa936d08dd87fcc9a3c54f546f0aab67905582f2a0ec352e2ec882c240e3c12fca79c423ccf00256c48af1fcb6dd8c52dced;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e0d4cee1fa89a63db5812940352a1b9e3085071f7ebcd828e4f30ba672e0ce8701e56e006eb7f78a21235b80df040e8022a18bb289198;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d5ab5b5ef2dad33fdeb0e804c8244ed9abc0a2fb0bf7dce684e1fe9b30ffbc5ee1a8f7f61420aa55f833707602552ec72bb576db960a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5516bfc1f86b02d55f80e60b3bcc0b59610c7be9ac4e94e89dc9485a099f6bc4ae291c718cdd476df0f57686b02ac0920415c4a4e01d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18257d5f8143afbfb06d055ee42b63b84a635f386e08b1d9042ab5748ba9ac9adc5746a368d48deeec52875e2e90d4a0dc0a7c43c676d1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47ae98b7b0e138db83a9c00e67d92c657fb59585bd82f4f121e6596140fc80d153625081e8ee976f4d700cfc99db7bceef0f8d3f03dcb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb49064eea80b215661909160b3191ea093ea983e516ee58e7fb0eff9319096e56722f7b3fe5ac84d243ae18d1e31bb9d3d038670311003;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184b6d7b9cefeb8b0148c73b780ed2ebcff541581e0450a8c28bd4fe0775f95980c4053647a97bc9c2b5f9a564967838c72b4e3984290ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130db6f19211b62fb56ce3dd55fad4bb867dc211e6c7fb965201688a5255f1e0ed297191d6abf93cd4f78228bc64a859d8f0a176bc6a3af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19128883ab3f170847eaaab5744a3ddc8671572ff2933f84111e0fbb6ad00748494d0bb187b5200a95056d249611e33657dd75227e419cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7ef28eb9bd2e95eb72067a5df75d6c08983e9103993530f745d803e77a4097f730ffdf3b0270bb57262fb3d9f98b02598f7fefc6d62cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb2386efd8fc559caec750a545a41f1aba0d5f3ffacceb37bc78897f2553e763dfdabffb595867c5bf4ea17a50e8916d4f5b618299f03f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192c5dc9a04076f6359ba3fc222b8fe0ac56c4b07cd5710c17a7e2cdab1d857a05e57f00f3b9dc4f94f9a6fb7ef035bcd845648b358a070;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1797e938bc03a10ec766e207d752765d236f7a071a293817eb4f4fbd29b10e3c3c1cd931a17abaaaed269a82f0368014a75dabe424fe6b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7f925bf7562ab527105ac3422ccffcf7b862d81345e189aee1f45a5f4f718aa8d7929f2211040084d6d7ecbd3efbfa0971700304838fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h340f1d5e8512918a03d2ee0cf371bedfb1b5eb87d1d54df5c6315ffa029084f42ffd7cd3a9c174dbd351a0f9759e9c5606e92db95c39f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b174a3d81895b312de3f2016d9178d63dbf956ba6f6ef42c778bac35f7f2da09bfa2a0a789a8c8d1e19aa53b52ee1c07d56f7c122fdaa6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74620114b5cbc98f20353014f72feebdef7d915da93bf2751ae5a12124848f8e5b548a147efac3517ee5e500dbc3d903337ede5de5cf1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15308ad2d407b3f77c91ed7f2b3fd0adcbe549efb6339accb36c6b69b3a5eef9ae07d9056825139558dcb442640ee502c36d27fb3e0ac10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a55652fc00803f4be3528d9f2fe2960ddeb5a55f166c4d817275c7b0b1c4bc115d174179deecc2b3abd0571036d2546e9da50a43d68de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c9840a3eda8bee229a28effc82e6e7f99f592098a9ca5f068b906922699c4409d5b037991e969a1df2547aed7037495a087002fedbe43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c3f99ae200bd86535f0c708fd4f85ce1486b757fd664e5d01b15ba8b03d46bcaecd7137fa613d92ace016fda882ed9f8a7b493b39c9611;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa1c042269d698072a099e4d332a0795fa6f9a71213785bef353c87eb835b009659c1ec17a705e9151572ca4fee05f17ca5ccedc0687b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc932fdeebd8acaacbc73b8720b2e73d8bb675d505f40edf9f5606fdced49fd7d8f413c1813ef3d848418e71b0b3e2ea84f5f9edb41c99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ed955b99d8649e50b3596f8ce4d1cf52508eba6d9a07effab9b7207d1567d1d2df7c3c5e6db42fc14541ebfba5fdad220674e5a03e70b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182ca2f9ca2421a9fc6186deaa92742be7f042c97cada30d391d6e026f701210fabdf639f86a1b04c23d67720049239bb7c42c62f6164d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h676dd968ae4d395fc228626bebbf60737cc4912cac63b7caf349b101292fa51daf4ebcd1e2ff83e0e1e22e328d7225aeac1cc93b147122;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4e67fdc3089c9c14bfd028bed4f89e9eba74bc4cbaa3c8abdd042ad7d7ee1d30196ef0b975d1e64f923c9e231a4d1749e4f52bd16d0e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc76f90f8a5c6f3da867d9d7351360dba2b87310e7698940544bedfae00023fbd43a00a59a3738686036775b4a709e835cc16308eaa4e54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129a00c1d48e33d983e11c795cba906ff5765b2b6b3e46b296d3fac92c4df885cc34ce963d637ce61f59498ba6b2ab0981d2b87c0991def;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h948ee737be69514f60815a2d04181b48295c89e18bb194b39818e68eb8673efdf70928207f8a23fddf2d18f0196b3865731bc99b410552;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f04b6e114bdef41f35b925fca92745893f9a5f660f20d030c213828007c8161311802876fa36c9bde8220964754b1dca756a5c2ede83c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52e6a39b5ff9f3a8e5f1ba83024b76d01cb5f2f58d731be3e98cf308174a1b889373f28ca875c68675914e1990799660abb4b8bb3f1b1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha6143d0f386554c021069795c070af34e0bb1104eae82a55efd81bef813a233e5ec39d981369bf0c6a7e63c5b7afc978e297d6c1a8e65a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce0b6d040151fba7e3c3cc63a6091352a383ef3a8143dabfdb279c85fd97c3668c75e60c090e13e44c192b729381a94551738716b9fc18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a811ad4adfe23bb13612865d8fd50187f3eb3344835f3b1b8bb928df4d92f91a6a2f78fafa30943328528eccfd1c93d8e2093aa1d209;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82525a251a2a47abc49f35267ad879a1da35836d2b9095ded727bc2e142c17fc93d195708e50e83b059dcb2a708e9cd2eae645c545d4f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a71704fbf5626b726f0f80e44a09d1e5542c8f8dd9365d112b9de7f45733866e2cf7d26574907868830de3bef609bcaf7653ac164ca178;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf71554627e745b0f975dbd2246bf7dd7523787a4d9d3d81ea80693444a0a83fa43baaa078090baa0c86c82205415700dc62443a86bfe1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195389f5741d9ffa28b95a73de97627cd281915ef3151e68b4b3f48112db929b0fed68c93ffdd89063fedd8195ea0638f77329895b2a050;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b24145920240e6636f39d710dc1eb179c6c60d7478d57e5df3ec0e21947ba729820fbdd7e8d0a8a59e58b4b430b8e0030ef3ead766ed51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h311f731110c2589c4ccd2314e20d8102e01af3de98cebb53ccd351296d24b1630c044e60ba3208988456e08bcde4e0448d5ffff6d08858;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14382b9e1be3afc3db6ffa084bcb8e0ee5381432516924037d0c1c4d1b0bec9b0f9ab37e7ffb678d98d82f9541c2042073624e1c090c50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4ed97c6d7c0ba06bb5dd1bebc6de6bc4ee7a26091a6236f2c06a2461ef1bacdef5dc9beff714a60bf7f5680d9db81dc237e6141a197a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b85d195191e41fab826b21942fdb9b4f6b6049aafcee98d6a368e5de759a17388099f79d559658b785f4bbfc2aa021aecb5fdfe2120b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b696232a7e8d9dd5441323cd354c92637b8304b02b1a5b20db33a5896ffe5588c6fc29c354b7b6df2c08e70bdd6033c089c817cd486d4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f835ca1e7e681cb48f1528ffde923cbf317558b3ce071bc91b1bc3028579627be5d74c2a676d4018320fb1de64159ce4d12e22451b1b7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he075e0fc27f3626ac47638205857ec13a4794c841a8d89998f9f4f6794aaa698c9fd7c7cec6ddda6a451af94b5c10f266d243e1cd16ce4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1241ee0d1bda43a4b19f63b13cc9053ba90a2756d083ecc69918ace805ae838caaffe6822b6cda674c6a8b3eb0d6abea0c1d832667077a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2746b060ac7bcc94cd5f3b59749666aa6d856bad29146f2125de0b20e136cdca4c8b00939ed105c1e54cb664f5fc3d4b0026dac224a347;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172591a5441fcf0cc704a460be923768d3364d4b9ebe5d83906c0025eb212801b7937bfdd0d2e2facb900fc6674cee9c9f38b81a686ff17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc34a838c1d16b708262d0f40e59b5d803e1a1e02458fca62846e83df2161224418383542b956361c028225ace76da69a34246c835d94da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1254c1c0d7b7eb8f3bba7ec571fbee8f8bde996998901a0ee1b1c3dd2a6165bbae266c915753123b5bc2e4eab73fb4fa79403758f9378;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h729e0837b05b30c53b5023c64257633a80b6528fde8eab3f05690654e19e9c81cdc15a487122a120fd2ec454495545d271161659e4ef3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12236e56302532c241b8a4633d09a381467aba0e6895e97c463c74ab0e903f4178d1bcee8a844703bcfc3b10aea45d8a672460c61a27a22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52ed583e42163bdabd1f16aed259a78a782e4c398359d932cde440c8648237eb02ccc3e4647061a9d958591993e03c93d347afc7f6bf36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106778f15d1dda93b3af3e1b60023792588dbfb58627700858405658fd858e0c8be9b6465921716d0c4540c62abf95290034f531cec8968;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e29944992246514eb6fa36efe1617772f93b4e35bf05536791b6cfd01a937bb772b82ad31fcd49734d18d38ac958a5a1c64dec21af31b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aedbac9a04c6df814466d069f6447fdfaba6c92b71b181dcc8525cf041a543b73740e1af9d2dc9b1df61f0ab21ad3e5d78328f426e258f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1015be8c555ab91f303571616089baa5552f7946e78be06a6f47b2a0307a8432fe98c9225744e3c4e5f27f9516f5029997e0a2150883075;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f883b5b7bfd68b41e82a94e369870bbcbf69577c1beb349e263c67e18ac8b7d0493d32cc344f3e8736621d4e5b660c64a2b950f3f174f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e5f87e96329cf58ff1fb62f08e8dc8d96d46b86011a855252fc80d6ce19b9c321c9de143511180e4649a72d831f78ec0cb16bd97fd671;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habf265c6ce46fa9d97949c739640a4a9d6c005bcdb7db6875f0123e5f9d1fc988e64da396070f4c2c48950f598972c7daf393b02535e3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb7189ef64da9ce752b0ee5d31023ea1efc0ecf11f556235cd456769ddf45a357187e48f21454f9ee54d920063c7a76b3da607543bb17b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0bc7ab98c7dad750aeb974afcb3a774bd41578dcad70e203a8c55b26a17a259998e1129f0f389ae71736e0c14f664eaf2f4cb8742acf4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1b0599194a846bbfea966ad7b30a5d87b352a72694994b71ab90e2089166a7dd4e6daf5270b049644d9f186226715656b0b8d08452930;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd165a9d64e0d2a366184205ee9ee03c26299890b8d748d0fceac002ac350675fc7f8c81c8dc7c2f91532f25d4e7d86708fcd0e2f584aac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d9b348c97221bb04d368cceef1c1c4849d9d0cb0365a8ec2431f2f3d82f59a0a21b5b0ae392038cad0159310175d21cc65fd260f55e77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a5b413aca8110b9a624cd41dba0ab216aa0e73fcab62b859dc60cb115c5e6d0034192e37227fe72220d068d1b13f2586fd9c4bc8a2a91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0e8dbd3b25d98ee4cd5c2739cc0c55145c1de9d6c980b7e47ce1624ce8fafc0ab80231a1ca112a848f1d5a3c151166245f46be070412e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af5a51dc84e3c7992dca4247e1c3ad41da7c4b23a6dc37d19cee6771df1848487ad8f3845c9d7b8faa45f08e658fe06de7d2ad1ed680c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4be343ecbf8dd6d17a90ad28f8c722f9eccdfee890e94918704c77337d831d032c4d2e6a1bb9e67b4e58a3ef46599c1a09b31b83f81ceb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139e669430a8b340bbe7afe96b958dff05eb7fdabb11eb4b53806ae5a7adac999f9127ed1ca061787e7866ce675d8f645533fccc901cf26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abcec04ef0c5dd731532fefbe132671fcf643c51481155754654c6b35e375ad77fefe6c54a2fb75bc2ab4e76e162f143d15b70c8437917;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194cdeccb43fde2041286664f633778db087936a080ac5f65dc000563871f35cbe909f1aec7ec3bc1a1493572ede8cc9b46de36b3b720;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc436e1f8038125010a073ac78dc4d1b45629b8b69debb803e86e6caa482013361a426105daf2055ffcac9f1292575e67cda89b5c26177c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fb0e95683516f96948c77aeb6ebf77a965c2b87367c8235da7e005f35def6906eef1c73e3bbf67c6717493b2adeac559a071cca20730c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8d149ec1a460bb7b4863cc7ddeb4b280062ee6d0193c8c022c4cd3876e110346c33a0a2a40c905101523328635f8def5ae4a30577d7b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd60c897ca98b8a5843499229ec29cc279dc2b392e226a401da3a1da7633c7fc35f9c8cca1fa8873e8fac29b1b5a6d5065887458c70ee7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd111dcf0294fb305252178bd2c7f4d2e3882cf747ab337225334870ecafbcd3a7f10778411ae3b782dd3896cf428f16753c07afd10401c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h786f45dcee19f776a63ae5f62e66660c78442911d5470fad32a09c631cbf4693b040cef059847ba868a3b8771fcdfa41a46a026297d4dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heeb7c836e3ffbb0470be1479eaad125910e12e901f712b09998ced0dacf2926b0b151d2bdac596f11a6285dfd62e643e98b7ab3402d5d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15788a039d8fba9faa106d944971de556779d4d6ef9dbb1b21f39d0dc03a7f911a7835c95b40d2dd22d30b384126c2673bf29b0d3f0e3c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd0378b71f0b353a929f274a6d55031ca564e860ff2f34b2d5cdb46612230b63ab4654684ce1fcff563ea7d104adaa3869a7bca5d6cf5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce44c078a7805dc0ce67eba821bea1ddbf9362805017d973f1ae86e6e6f095d84e9903867f9e10a7345cbe2a5f66d5b9360882ea336d5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0d37d2f538f3c3eb3d7728fe7a876170892c03d528a6c299a75eb9bb45ee03f3843c1effb6445a26886e1406232f47545361b66320e70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf41b8b1bbe337b6aebd6216f2929ecc73521b779bb1ac106171641fc829476146533d3761c8d7b4d38268c383330221ac4133291e5365f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170738c30de373604d00578333bb093cf87ab55215328d5bc015d9c5a97747ccffd702177603e443d074cdc9a157ff6ad96a4816dc68a37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee67246fd39c2f8b914f850f9ba9c86bd0f259a574e7d1d351434851d6cd3d6c75cbee4a7a722c0916742974c1eab5e9e27fc972c6ec39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177a6679f611ba09f5ba797b04e562e438ee8da046118ea76e2aa30af8894eb62f497f648140d8c75294bad3d5c86e2298208a3c5bb0180;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b59fbf473c1fae8c39decb2115be12900445aee59d4d43ba3c919704bf39169176c018bb0fc16dce6cc012d1f8269512d5b5e61bfacaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1824fdad49bc5227d33218cd8ba7d07a6a9b1a2c05a63ab4bf88182619ee4112e067fca9de0dc1c28fe9e457e55637abc1c496faa1eba77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1051238b65b78d902025e6d00e853463cfbe3379635cd0bc156202fc6c60005b3245b2403ba4518afed63979e735f63dd5a2696d2fb5a37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38ea932ddee975feda45f045fd7aac1b6825dea6df712f09984a529d0faf8cd183f15d92a7cc17ba8f2ff6c78af47a137000ebdd78adb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d1217577d6d607a25d3e03c46e076ff187b5443086e3e5b563c6e048d69d50bb241a2921e8a205759f688600f7559633c08ebbbb9c0f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8217c7abfed7bf7e845827da5c6cdcf251cf5b3d8538d8c06c6cd489a8f54945a2c0bc39fcf1a9c6fe576faa85103b8286d0910d539b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5de015cdc1ab3c2afd1eb23a4297e1ba80b6d9131da00dae95223fbd4ca7e92212c81808b65d9433c2752a270f673eec409d83a559f8d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c055ffb45c3c1800cf677a0ac36c8bf76d40d27e53a3988dae3ea7e9c17916deafe8c60b091c17ad30337061f410870bddd82604ba8d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc77a5950465f5b6f21d0d62fcd394d0b58c58dde97248c40ff266fb18e1f237aa64ee5f309c7a543784ddee56d625583823b356932281;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108b96cac0a4a52f05340e2f52c2a701c544ff37b540d3272f23af7ff6d7cc8c64bc07188180f342d9360eadb0f71f337170b7fe83410e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he528e3ef93a371a1e38ac54b15cc1bb077a1a888a6e40c56ce87dbdb8ea353c865fcea93f7ade107d6422488121802c7f21e1421f031c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a22da6a52bb4f61aa64c5f168fd1e76585425de7b9ab970235a6a535ed024b89f4e7a83baa53d9418248ddb8e5ab650295fd8857d6ba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a80a116af299b5f3072f5b048f8183881503d26ee3411769425b3c6c8cd57c141ea3004731a01836207dfa25584f836171011b4a90f822;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4f221fae6768268292c4972f553041d64319fb6ff0a2b59d5905ad0dd50abb2c3446aa6e3355795cddae011b5b54ecaebd5ea2a26d714;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1451190df4f23b0f489cf88c01fb91bca419d0a11d2ba43ab86b672e80851fe73f3eb1c5f0122dc2af1c45f972004f717703c66c1be4edd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d5bf77c5a6b2cc95a00e98a4b962411610b932c2c48103941b78e40be9813994529fcbf14b3404440ea74c812013b7aac9f25ac22d93f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd73a6c97a2b1f7a1f25d2d44a49544b136cbd3a85360eba4508f8785d2ad6a470dcbd19b4acdd5feefb67fc6cb47887c38d42d30df132d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5acc6c1cfc392675ac86ba7c19288e614f7da156600bdd4aeaa5203bb2638e2628e359c9e75635b97dd276cc71fdbca2252514db5cbfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6f14cad36f4f8cc9ccae01f918620ed6a739bab59fd8e5c6b250f7d98bad9ded881059aa41bffd08e28a2c68962fadbda1f54bc224ba9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8e4e2d9bf0043e86f0cbf1878aac9d5d6af1c7ea0cb50aaf27962730db64ccbce6e5a28a92541711985211d7872684ef0b6818a5678da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1120ab2f86be691fbacd684db4190c8b7fcc09b631c2a3e4b6d3e4ba26c53ba79fa75bbc69a14b0e358bb623f90d4b204de8826872c3e7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5be94e55080ddfb0eb036c87d9a04724099a10eb611b0049aec4f5b1e7a8881bcf35df52c75eef1306bd7629d8ec6cb93418633a953df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cca7d9381b3d8a9599ab3ffe67ecb7965a9131e390c3eff35fa40c5d86d5997b3cc019dcf9181ef57df2cc64d259f756f097b4a0fd73b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bc548af8be98e0bb5b8f3e266a07044dd9d4ee4a2d54b38612b2a07a405d0ed7414ab52e9fd9aef0ad2489a9110b1790517eb9003ef69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f523ab1f8e6277e60d9259614e39e0fe5a74a9db6a6660b2e5cf0c981c53a27153c3557bc2c8556ddaa3daca14617ce178e1793407e618;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bbfb65c17f758e47746531db4bfcbb01914cd0200f32bbd5ea2e44decae0b785f81dcf49e8fb4e08cc88602a56ad27218636d12fe0b08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5cb7503f1ca82b9ce9e7e9a5e606ebbdd54fc2dbbd535541aa597a258526a62bf11b5d2813d914e7c03ab53d22c840919170a4d2175a80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7da0a00bf49fbe884f9b30ff2b623c1d224b0d0b6d680cbcae2dff0abbf79a4656d8934c03e0d7adf73914d1297075a7d72957384b052b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd05c2b2651d2ff07959f44204259eb4e7ebab517f5365d325a36fde24b7cd545c32e9c9a3dffe71fe9870c1f55e521dc0dd85dfe1c60a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168ff21fe790e0d77b6b6eef3424864b7f8e2f41d8cd8d544bb887ea8248a6b3852dedb0f599e69f33b736712bde445e137888ec834e3ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h989349ae39fce15de0b413331e21dc5ed34807deef45e375f1062e907174cc3c085dbf2c5c540fb0565568b994c1f21394a2de5269bc4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1771d5a7598ca0c33e1cbf4e4a3017b039344ffcad21fc7b25288d873ad53c2416edae94af2db0dd6f89603d25a1344592c4ecdd19607cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2111bf9cf2680329d0d21bc175c06eeb728dc460dedddfdd803a963765ea1009ea9b465da8a5e4c897df494eb7c6cdf85636a882100a04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147d1e549ca0efee26f10bad3ba92f1174b552d2518aac0bf5cd507d4dd40f45361646d63509123a93104507ff1dbdc1a74ac79d8f580ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7aa9ad949b389dc26b818bf08ff0a5f8662ff1453d4f215b347dea78ea873c91e84181143f3da95503236017bb0b93539a2b49b48ff64a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c91efb05f7924b0eedd336239d24484511f4186f024edf47b802bfcc21ca3fe161b97ae5f95a7fda378e336120b0090dbf33d1272b3623;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b897cd9c7926826a9a5f5bc3a08d0a196f072fcdca17b3bd3a3363245eb346a6c27bab6ea4aff6330389f525ac1770589c782917fff42b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125fa1e5743e11eae147134aa137056c6b04325bd838eb3fa3c37f24387bd6e8deb8520d961ead361aaae4ba6510f7169a7aec425f567dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cefc2ade4a2d7ecfb22d53cf6a00fa3ae5e45f80bff4cb584331d01eb77f3f1dd15b3758d17546d18cb078250bd619a465d0270c05d5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1d923103507787d35104b2f7d89a74837175e3f7072bd842e72bf183b54fbade0f840634c9c546f454dccdd55dcc6a87c58137e082a63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b79057f4e5e44dff9a11ee0a0344abb1fcccab371698079c8a4fc59552b5cfd07caf716f334d20f3af1581137cb7eb01d764fe630c031c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f39983ba886a2e443dc23d636f13866810722f9af032fe0ad3965ec0b1b70e56ad4a48f22ad3e0d2a6a5ee0e15e37f43f178ca0facc19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146f8f685fd2e9798a4ca00dad6b27c63c0b2e696035ce0a13b83a73d1fa06ae923b7d236ab382c5f93d4082f0c8ac734d17ef217a8b510;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65cc10d2216c663c3a78953d93324a4eadd9c2ac78340e6884ec720a24f6932cfe3af9c82855c97f0e9bdd9146e8803d7c2eee29576984;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6d68aa37be5d8782e593ca8a0289095d9cc1415d4bc44c4d2ef716c4772332d1c2ce9a1da296235e86677f650656b4c44a1bf9317c965;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175e90ccb6b190cde661101d1ce8f93358a634218ef297051aa1eeaac3a82ba88d3bfae1bd53723ba8761d135d46a1bf6457b42f906891e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2ec53b7073474f9066ad44cdb269c8ae31c7ea2b139a288dbbbc4180b5e0e1f64fc6d7d94834eec897b10f5c295f541bca8d4949236d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a4330e0ad4b03cec6a3fa04a1ce3a848caa317414b7fc4b49a226b58e2c7b56121de2112c6dfda368620214ec63724dc8c112904ebfda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28940d75357fe47adc958977dc3683cb9a0fa958077da60fcddd595385137397642da46132d3f6e0fc6c283a1efe82c6b3f1c7560b773a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h949a4ed266bad56c84756515f6b44b7c2d2b9cf887c09d20da39e38089d75186d7e94541ce528ced4acaca8f7b1ce379a01aba8f92860;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0678c443901543e6d5d643fa4bb8b07cf46aaf6ebd6e21be80cdd9873b83ee301014ab420c6cc5a97df721809e834710929febef8b48d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26799c98aa0cec546dfcdc8a0d130adea8904e70b469e19bfdcb25efc5a208702b36a7107b7ccac886fe03d031923144657de439d411c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e28f1a37816cba5b8c8b6b22b2ab460bede786c2ae7a14932b9cc5134a1a7999f77d85b6d9134f013c6fef22658ed3ca6aeb695607d32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6f10dff5b38ef4280bb5aebb409a2def009c32587d6e583255c5aa2a4f8ad4e822b737a669ed1e8871f3052a0986040174ea8cb60bb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hffc3f13f205d25670eb1b65ee2e8a606c8cdc6093cc0d084c548149303e101409b4b3068bd881b91fdef28402b3e24602bd47d3d5d602c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd005ae845765b6f44c63cb8622a5189e2a7f94c0d0e324f56920ac1bd7d895ea6c1618d110fcaa5e6fbe192d60c6a9f21704ebeea1802f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc359313ad091ae976f730b7605cddbbf5783fbeddbfac2313b02aa8a6e5084ffa3d9cd0f589cbf5dfed3016c14dc94cdd822432bc1e3f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d62d7685adb86a595d999f9071f32d07dd75eafe11a7ce9b80e1b9e17731585115e75d9fe9ecf76661ab56e9d12f7fb648b3721f7c6b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130b0e9c461281b8cbabc539cc0c2e081bc1a1478badab5bb66f5cd3208f897cbc2604016a54885267416b999389118f1a3e0e28ec1e3b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef3c898d16e9a016cfd6091a34d36eafc1163e8c6decd894f8cdd5ec35bf3706e42eed3ae450232ab041e802ef6a785634dc0c1b14ad48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac61f0d195ec26899ba7c6624768c819070253a61f155d98c33962a9ec034b5fbb1073846dfe260e5864985a4f01a8993222b9f16d6786;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f26eba1ce7a5222d25632a22d37c5dfbc6cf3d55e95d1b0ff05c37aff381f3fd2d4300fdcfc55082f7c5a6b20b9a6825e4b4bcd2276406;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13584576656d85b014fb64e3646ade696d318d8221e0cd80cb9ac62954247c5d29ada6f18efe54ac78f0b5d6d97e4ebc739f09cc75bf270;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197db1000154c5a3516ac02a3d89d0cbb484bfd2f6a043c7af728dd352d86de2e8c7758ba06d16a36697d6d0c8f5d0546b58fdbb32d7ff8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h525944bf8c1034002ad68e6d95bab3d21e3454a408e5ebbdb9d4d10972676f0913a69c5346d7bc575920ff0cce123ba6110d85f2c84765;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd94e213eaab09df775f4c49d9a82539bbf5cfb4caab5fb0be20b0f891aa47216845c26c2348f6bf7a60fec433fba4a8988ef9ef6c16b2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c10efd276cf4c1a17856a0b66561529f0692d27ca78a55a9faaacb55e280b7c60b85a9e43f9c72e16ce7ee8879388722d7d502acf65532;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61e753c56725c2f0025cee1be7c5e79b6b7f18c2da560b12f2a0fee7a25cf14e412403555684413682571a7c9f991138fe5e4b08e84d6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ebdc66a6299f92447f69c61c8863162e4a5eb400d204e9e5aadb874da87414f82fa462ded752a636db41f7e4245cfa8d741d330c9c8e3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2817d0796810e6ce69bf8e47268d52bf7f951c7cce85c2b41a84701731ec81d3d41d58938eb03ceb2b8b09cf0cb0ed0067062c2b68cbb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110a399a56f653c4a1106437dc25c131a8d66af5ada83aba1d6ded403b9c0e70773aedd04ea0d22a7f83aab4eb5cfbd977f4e6d34ebc0a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42efef9abead91ce5d8f7a36ebc680d533f75c0c6048af20cfc7e62b1d7e7f893f5d3c3f5f108155c752bb7f7ea51d61992de517e2a6d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ee316826e36aa19db39d6730da099d46462027a62e7c0f83ae626f3f1f2f771a0bc2036a57fcca88b6d1809e6ec26b7a8a49677655747;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15121ea02c850a467e713b4d9e1ad07845b3270ec53f0251d743106767a9ff70af6702f163c5858bb51f9e86a8a928f138c7fc885838640;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dd3ae760395d1cddc6211b3fce96803a3def969f975aee740829986a09599485f9228bc80863051c2af7dc97b269cec617a975b98ee20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161bbdc6a3805b47328b22d0f0e10b537425ee92956305e9e9d004360d390d6b256baee9f375bcb2f16a5937f2431ed3bace2b159565089;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1688942871523cd46c2df3d3ec88ba61ea8f09bece995e6ffd39f9b04ffd53fb2ea1aa77c36833130c5b1255d8b389486c6e0cb14ba0021;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d920eb69a95ef6de01c397137ab7a589f95d7670af523822ad2c4c040a83aa583e9aebdccdaa98091047200d67af2ba064371f32190aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae215fb418d1b144cd2a2135dc0516d46d0c078bcc01b331ea71b772e0a32c7388ad5446b8729820098f423ce2314a6503bb43a21ae72d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127c828a3039b14462c298712f36dc26266dd71de98bbd08c82d91a7357137d23bbdff3076cf501979d14d078e080ea07fe0cceadc015c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d0899c706fc54b762b794c2c7f0bcdcea462312a3483503023efb4f55c1814839f7b95187f0303305067d564ff2240b71d231debf35ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f42c962114d8916328cb769daaf442d02d7ce46e121766c572f725c11e60236d240d9eb5b9d77f95f0b68bdf1d9dca30272e3cd370942;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12419f0ede1118a11fd4feb566443b35cac762819b49dbbd0c4e7b6b7877d5c85467f13b0b44f621bd7c27ef94734e75f5f8d9b7992129b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106fde3292c484eaae6438b9c08370ad577b5abcd99296a705c9a5fce891bf0943b14d232c15b76682af29225c088c82450e9ba9c22ba6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166b084239c5401d75978c3413f4dad5dbfafc948c3bbc62ec4aa8255ba977e57fe5eac2813e5ccb4a8e2bdad82fe404d5d0390783e1ae2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd4f4cac100ac9cde593d3d5c859f195c7a253419dde91529e1809ee85d524eab333946819b71549bec35ee7480acaf1c7338173f08d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b1c53b1f4d5ccc1c48785b1d6cdd73edaa590fadfdfa715cc977215957eef1473e04d5d4356dfb4ffedb6fd177c7023da101854407b65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3be384b4cdb80c7e25b160ddfd0470ad6d1aa22faf6f78504bfd4b7520f277e2b4ba89f13228f2456bec02e0117cc6c7b507e126bfb3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf9f1de42c2390a07b1f7befdec1302282a4cfb17e419481204184ebfe0f13cb8add8481dbffb30a4d60bf66954168b5d7a7c85f74d4aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c60c1d8d1e0faa770c1d171f029c6a5bb16f39da78a77f8be1f2f768681eb8131ece159469bc4cb7fbe75dad1de61cb8d78e6c9ef51c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbdeb575c0dab47f69fca3260e3e0c1b5aa5c653c8014fd13706f32b937add1b58afb99b2a03e50edfa590ed1099f1e65e87cd3134129e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4979653913e7c81992215d3fc84cc06ae6ff3e71ca846b8eb112d78d36b15059980b03f01e3b89b3cb3ff9886399ddc153dfec8c3fb38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1347b26fc7daa3753bbf2ee8af7f59b3af95ac8bc52f24adc0c756451dad1ec96411c0a87966382562530d86ea55318929d957a6cfb9b81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9e984e99222a7d7bda23dd033f5a4c08dc344d276db46defd8fc22ca29727d5908face71302592ac8a6391260f12b61e2209ff4ca0673;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4988fe9683f43f2f551f15d74aec5f9ae3c412fd1d3b15774fa7e43ab4b077edf83de32dc76d19340362e97d25dde3a1b7acc8361dc90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1802de0dbc7663bcc1ca01215024876a64863228d8e6ac5bad363a9738542e0b815112c976bf7afe7a8e73eb6821c91e9fdee4de3511a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170953b105845a67e8fb7a96ded9338c3bbbfe3f654e6bde954a87340f7a177b99907026183f3ee40ddbe3aa524523b33cc1e6145a25026;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ca81bdc85e3ccfc1740727eccbaef249db245ed6f25d0692c290a0945b7e1a7c95c26488fb415fa8c125527bb8d80b2cc65c21e6a9638;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ed9d00ad1209cf79cc950a953d7c300011c500347d93463db1e18b1b3c3479e626401c4e1482d26ed408d52d2f787002e2f437b89c220;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf3e3fbd0d91e34c6341819338165220cc34c665fdf924730bcacba3f49f4a1f049979afe74704f915650e7e2c80b9ea9532627aebe0a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97412732cb764a7e5b2f6cbaddc806faf6f7c629aed296a76efa9e0c24eb18fccee64d8d9d78f61234633fbf93cf21ed8528fdd81163fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4ef79db9d7a730e0770a03ee12f68595dd4c473357a51fcba4970d734b708d0f5676e0775b89f5e23dc57ab439cede1ebb4507bfbe68a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c009662092c8d4ae5e9ab331378fb5fa6354187af8c848d4269fcd004e6b64d63b341a37e8d5bf4a41b7d3bd811078f5f4f5ab9429284;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63284ab3bc644732ea4d45093de610df01f4ea6c23a1099e3bdd9169c3b42229a3afe2650e6e2dcba8c337245a07009e291d91df3c9244;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147fc4bb3d2a8ffa0afe0864e797dbd291c5274f019f54fb4d1cb849b104f7d2c5985ffbf0107ac62a325a643cb0350d136ba887750d2c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2400c4b88a324abd0e26be7252cf033f56bc7adac10379ac6b47467895cf6d845c52426f9a82a08310689245b734ee36b9b4d67654f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h884b10336a21a36ad08784c5c2b1457ba81e9fbeb5c4d72975948ae395998693fe21633578fc406cabfe5e0e6b98a494d3ac7975034c71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb57518e01b28fed58d50809f36aaafce04735b25ab31c22635ed34fd2aae6481216988735a8c0429427e2ae96893fc5d2a3334902da9e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9b5d9934fb942617d959e496af8c7da1b9574c59f5a7a48e876d477dcbc8e283d0dcd718a1b73905f93851d1d4ee7b085579aab2ce5a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb023a9fa5b01a538e2b91972a19b42f2cba6553ca62bca04fcceee90269ab2cb96bb96091a76d66278f895208e740a51492e69dcf18f20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf4049e149e3cdf03acf59a48c4af21e06099c7f39a0ee0318e84e0b1c381ac4fd59ba14b722e66291df86e0603bfca6222c0d4595a978;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d91565d5dbd49e11da1e45f8fe99736fd5627583ab66eb6da1eff5e3d488777588231100bfae5587033abdbb48c082a98003a0f0327df5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hefad11adb25fdddc30505a301e01cadd45ca323dd51575db22fca2b4d5b5f6b223a50b363bb2938d42bccb37b2093c3b7c9bb7f354d196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164a39a26e45fa375e47f842d19e551e4af5f7f749baa8353bbbae8af33572934eeacf591dfbede318e22668ac7f94980a24f6f2161a7c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15aeef33733a98c626081b9bf32502d2195c34128e24a9f72c6660638f1bb76fd2a69fc8ce2703016611961f5c3dff60ec0be93394c6ade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15cfb7c27507d7d075d0af24c979f359508ec62145dfccce7aac54df7dfef15ffb8f2dd37b16755d4387f59c97f56b4deedae7a81d00f09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64dc2ec3bd93a64d6f64b007718a331dfe06a9373d4b38b9d61a6208bc08a3709ccaa59eb370d72e94b4647cdb7434093032ccf570369a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d46371bce8d771606e5d7f73e378fc0d18fe3f373743fc0f1b3c38f942cdbf3d4a4e8b31d70537e68f1ecf54641b78db1bcb9c99626a51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b427d54141c9e5fdf4f2f3f73ce540d6c29d3cf2892bdb49a5232c26f5b1fab8991a6c5b298eefbc3e91ded8c371c413cafe1a629d52c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1760cbcda1df55770b6484560527a628820e1afe5c67247b1518fc17c484e9195805e79560c9d4da2adc74c9895298d85776d9cf71c9b23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1530a530f0027b61a6640728fbebb6e27485b00923be435d71ba62d064d5c8dc19afd1eeddd7b6a272c2a04666a501797e555b9e21095;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8cd15725ddf73c182942c7b78a8dce5791ffea5b0945c30dc74917c6d3e47e2a9c732d0e4302be8e2a0e51bf5172f0f3ec10a91040a45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a46a8a3228b80f043c5d60fa8fb5ca3ee52441a81b79ed864b55627fb5a1d541b1b56e9b66cd361466043c78c81607f7ad03163cfa85e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b10c4110e83dfd6f36c60a5a07e534ccab762be00b4ad8ef2bde3e5d4db6d01bf83fbc4aeff3623990f035ef4497ce9a85fff0a5a89c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h638327fae57bd06bae89fd11669ea0ac086372bc332467d65d411af2d7b9cebcb9fd5e83ad75c340981128705e40d0dcfcd332ccb2e62f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h922647543c28c54c74e61d72009c14a2ae02b7513bfab3dcd8980781b55e0561f45b811799871334ccb9362a2b48afa2027e0a3d0209a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdc9752e8dc40dcf48eeee25d6c952e215a944ebfcd3a3b34b8affd9182711f7b8228368a91d33161e2853b319abb2a1d161fde796ff65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadd7715ea60e842f37d97d7c14081dd6ef8b47ae06d0cac5b3173072d8ed23c86cd9b80475218f254532f8890e5e0647cd8c7c07cf7e01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c4a56ce9757c0317c05d1fc05dcb905068cad5450d0e8003ca269b33ff86c3c452a9e52adf749699a67cc5a59bd855da591b41233e6bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6501628f7eb992fec89246c1bba661c7ea472776833409b1345b2e8b89d7d4cfdfccbec9f84fabd3fd1abebba3bfb0cfb544238b77db10;
        #1
        $finish();
    end
endmodule
