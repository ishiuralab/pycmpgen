module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    compressor_CLA512_64 compressor_CLA512_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
        src32 <= 512'h0;
        src33 <= 512'h0;
        src34 <= 512'h0;
        src35 <= 512'h0;
        src36 <= 512'h0;
        src37 <= 512'h0;
        src38 <= 512'h0;
        src39 <= 512'h0;
        src40 <= 512'h0;
        src41 <= 512'h0;
        src42 <= 512'h0;
        src43 <= 512'h0;
        src44 <= 512'h0;
        src45 <= 512'h0;
        src46 <= 512'h0;
        src47 <= 512'h0;
        src48 <= 512'h0;
        src49 <= 512'h0;
        src50 <= 512'h0;
        src51 <= 512'h0;
        src52 <= 512'h0;
        src53 <= 512'h0;
        src54 <= 512'h0;
        src55 <= 512'h0;
        src56 <= 512'h0;
        src57 <= 512'h0;
        src58 <= 512'h0;
        src59 <= 512'h0;
        src60 <= 512'h0;
        src61 <= 512'h0;
        src62 <= 512'h0;
        src63 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA512_64(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    input [511:0]src32,
    input [511:0]src33,
    input [511:0]src34,
    input [511:0]src35,
    input [511:0]src36,
    input [511:0]src37,
    input [511:0]src38,
    input [511:0]src39,
    input [511:0]src40,
    input [511:0]src41,
    input [511:0]src42,
    input [511:0]src43,
    input [511:0]src44,
    input [511:0]src45,
    input [511:0]src46,
    input [511:0]src47,
    input [511:0]src48,
    input [511:0]src49,
    input [511:0]src50,
    input [511:0]src51,
    input [511:0]src52,
    input [511:0]src53,
    input [511:0]src54,
    input [511:0]src55,
    input [511:0]src56,
    input [511:0]src57,
    input [511:0]src58,
    input [511:0]src59,
    input [511:0]src60,
    input [511:0]src61,
    input [511:0]src62,
    input [511:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [0:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], 1'h0, comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      input wire [511:0] src32,
      input wire [511:0] src33,
      input wire [511:0] src34,
      input wire [511:0] src35,
      input wire [511:0] src36,
      input wire [511:0] src37,
      input wire [511:0] src38,
      input wire [511:0] src39,
      input wire [511:0] src40,
      input wire [511:0] src41,
      input wire [511:0] src42,
      input wire [511:0] src43,
      input wire [511:0] src44,
      input wire [511:0] src45,
      input wire [511:0] src46,
      input wire [511:0] src47,
      input wire [511:0] src48,
      input wire [511:0] src49,
      input wire [511:0] src50,
      input wire [511:0] src51,
      input wire [511:0] src52,
      input wire [511:0] src53,
      input wire [511:0] src54,
      input wire [511:0] src55,
      input wire [511:0] src56,
      input wire [511:0] src57,
      input wire [511:0] src58,
      input wire [511:0] src59,
      input wire [511:0] src60,
      input wire [511:0] src61,
      input wire [511:0] src62,
      input wire [511:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [0:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [511:0] stage0_32;
   wire [511:0] stage0_33;
   wire [511:0] stage0_34;
   wire [511:0] stage0_35;
   wire [511:0] stage0_36;
   wire [511:0] stage0_37;
   wire [511:0] stage0_38;
   wire [511:0] stage0_39;
   wire [511:0] stage0_40;
   wire [511:0] stage0_41;
   wire [511:0] stage0_42;
   wire [511:0] stage0_43;
   wire [511:0] stage0_44;
   wire [511:0] stage0_45;
   wire [511:0] stage0_46;
   wire [511:0] stage0_47;
   wire [511:0] stage0_48;
   wire [511:0] stage0_49;
   wire [511:0] stage0_50;
   wire [511:0] stage0_51;
   wire [511:0] stage0_52;
   wire [511:0] stage0_53;
   wire [511:0] stage0_54;
   wire [511:0] stage0_55;
   wire [511:0] stage0_56;
   wire [511:0] stage0_57;
   wire [511:0] stage0_58;
   wire [511:0] stage0_59;
   wire [511:0] stage0_60;
   wire [511:0] stage0_61;
   wire [511:0] stage0_62;
   wire [511:0] stage0_63;
   wire [118:0] stage1_0;
   wire [168:0] stage1_1;
   wire [220:0] stage1_2;
   wire [321:0] stage1_3;
   wire [250:0] stage1_4;
   wire [216:0] stage1_5;
   wire [179:0] stage1_6;
   wire [339:0] stage1_7;
   wire [238:0] stage1_8;
   wire [362:0] stage1_9;
   wire [152:0] stage1_10;
   wire [317:0] stage1_11;
   wire [218:0] stage1_12;
   wire [184:0] stage1_13;
   wire [255:0] stage1_14;
   wire [257:0] stage1_15;
   wire [223:0] stage1_16;
   wire [217:0] stage1_17;
   wire [241:0] stage1_18;
   wire [218:0] stage1_19;
   wire [243:0] stage1_20;
   wire [204:0] stage1_21;
   wire [200:0] stage1_22;
   wire [298:0] stage1_23;
   wire [234:0] stage1_24;
   wire [210:0] stage1_25;
   wire [188:0] stage1_26;
   wire [211:0] stage1_27;
   wire [248:0] stage1_28;
   wire [220:0] stage1_29;
   wire [232:0] stage1_30;
   wire [211:0] stage1_31;
   wire [414:0] stage1_32;
   wire [209:0] stage1_33;
   wire [267:0] stage1_34;
   wire [190:0] stage1_35;
   wire [330:0] stage1_36;
   wire [302:0] stage1_37;
   wire [276:0] stage1_38;
   wire [196:0] stage1_39;
   wire [229:0] stage1_40;
   wire [276:0] stage1_41;
   wire [228:0] stage1_42;
   wire [243:0] stage1_43;
   wire [268:0] stage1_44;
   wire [188:0] stage1_45;
   wire [299:0] stage1_46;
   wire [277:0] stage1_47;
   wire [210:0] stage1_48;
   wire [241:0] stage1_49;
   wire [216:0] stage1_50;
   wire [226:0] stage1_51;
   wire [303:0] stage1_52;
   wire [186:0] stage1_53;
   wire [262:0] stage1_54;
   wire [225:0] stage1_55;
   wire [256:0] stage1_56;
   wire [179:0] stage1_57;
   wire [242:0] stage1_58;
   wire [293:0] stage1_59;
   wire [199:0] stage1_60;
   wire [216:0] stage1_61;
   wire [372:0] stage1_62;
   wire [294:0] stage1_63;
   wire [111:0] stage1_64;
   wire [56:0] stage1_65;
   wire [33:0] stage2_0;
   wire [38:0] stage2_1;
   wire [72:0] stage2_2;
   wire [253:0] stage2_3;
   wire [92:0] stage2_4;
   wire [111:0] stage2_5;
   wire [120:0] stage2_6;
   wire [96:0] stage2_7;
   wire [172:0] stage2_8;
   wire [104:0] stage2_9;
   wire [133:0] stage2_10;
   wire [135:0] stage2_11;
   wire [127:0] stage2_12;
   wire [71:0] stage2_13;
   wire [114:0] stage2_14;
   wire [114:0] stage2_15;
   wire [109:0] stage2_16;
   wire [89:0] stage2_17;
   wire [161:0] stage2_18;
   wire [93:0] stage2_19;
   wire [87:0] stage2_20;
   wire [111:0] stage2_21;
   wire [109:0] stage2_22;
   wire [97:0] stage2_23;
   wire [84:0] stage2_24;
   wire [122:0] stage2_25;
   wire [130:0] stage2_26;
   wire [85:0] stage2_27;
   wire [79:0] stage2_28;
   wire [111:0] stage2_29;
   wire [99:0] stage2_30;
   wire [127:0] stage2_31;
   wire [117:0] stage2_32;
   wire [108:0] stage2_33;
   wire [127:0] stage2_34;
   wire [117:0] stage2_35;
   wire [119:0] stage2_36;
   wire [113:0] stage2_37;
   wire [99:0] stage2_38;
   wire [107:0] stage2_39;
   wire [139:0] stage2_40;
   wire [122:0] stage2_41;
   wire [81:0] stage2_42;
   wire [110:0] stage2_43;
   wire [137:0] stage2_44;
   wire [131:0] stage2_45;
   wire [92:0] stage2_46;
   wire [107:0] stage2_47;
   wire [153:0] stage2_48;
   wire [115:0] stage2_49;
   wire [152:0] stage2_50;
   wire [87:0] stage2_51;
   wire [127:0] stage2_52;
   wire [96:0] stage2_53;
   wire [123:0] stage2_54;
   wire [110:0] stage2_55;
   wire [131:0] stage2_56;
   wire [78:0] stage2_57;
   wire [84:0] stage2_58;
   wire [139:0] stage2_59;
   wire [110:0] stage2_60;
   wire [101:0] stage2_61;
   wire [144:0] stage2_62;
   wire [112:0] stage2_63;
   wire [101:0] stage2_64;
   wire [67:0] stage2_65;
   wire [53:0] stage2_66;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [14:0] stage3_2;
   wire [51:0] stage3_3;
   wire [59:0] stage3_4;
   wire [54:0] stage3_5;
   wire [66:0] stage3_6;
   wire [54:0] stage3_7;
   wire [46:0] stage3_8;
   wire [52:0] stage3_9;
   wire [67:0] stage3_10;
   wire [60:0] stage3_11;
   wire [80:0] stage3_12;
   wire [46:0] stage3_13;
   wire [34:0] stage3_14;
   wire [50:0] stage3_15;
   wire [58:0] stage3_16;
   wire [43:0] stage3_17;
   wire [63:0] stage3_18;
   wire [45:0] stage3_19;
   wire [57:0] stage3_20;
   wire [62:0] stage3_21;
   wire [49:0] stage3_22;
   wire [48:0] stage3_23;
   wire [34:0] stage3_24;
   wire [51:0] stage3_25;
   wire [51:0] stage3_26;
   wire [41:0] stage3_27;
   wire [69:0] stage3_28;
   wire [58:0] stage3_29;
   wire [38:0] stage3_30;
   wire [41:0] stage3_31;
   wire [55:0] stage3_32;
   wire [62:0] stage3_33;
   wire [44:0] stage3_34;
   wire [56:0] stage3_35;
   wire [55:0] stage3_36;
   wire [34:0] stage3_37;
   wire [68:0] stage3_38;
   wire [59:0] stage3_39;
   wire [45:0] stage3_40;
   wire [56:0] stage3_41;
   wire [53:0] stage3_42;
   wire [59:0] stage3_43;
   wire [84:0] stage3_44;
   wire [39:0] stage3_45;
   wire [48:0] stage3_46;
   wire [73:0] stage3_47;
   wire [36:0] stage3_48;
   wire [64:0] stage3_49;
   wire [63:0] stage3_50;
   wire [53:0] stage3_51;
   wire [55:0] stage3_52;
   wire [52:0] stage3_53;
   wire [62:0] stage3_54;
   wire [46:0] stage3_55;
   wire [38:0] stage3_56;
   wire [52:0] stage3_57;
   wire [48:0] stage3_58;
   wire [45:0] stage3_59;
   wire [52:0] stage3_60;
   wire [56:0] stage3_61;
   wire [40:0] stage3_62;
   wire [71:0] stage3_63;
   wire [50:0] stage3_64;
   wire [32:0] stage3_65;
   wire [53:0] stage3_66;
   wire [14:0] stage3_67;
   wire [4:0] stage3_68;
   wire [5:0] stage4_0;
   wire [6:0] stage4_1;
   wire [8:0] stage4_2;
   wire [21:0] stage4_3;
   wire [24:0] stage4_4;
   wire [46:0] stage4_5;
   wire [20:0] stage4_6;
   wire [39:0] stage4_7;
   wire [34:0] stage4_8;
   wire [13:0] stage4_9;
   wire [28:0] stage4_10;
   wire [33:0] stage4_11;
   wire [19:0] stage4_12;
   wire [27:0] stage4_13;
   wire [29:0] stage4_14;
   wire [22:0] stage4_15;
   wire [32:0] stage4_16;
   wire [22:0] stage4_17;
   wire [31:0] stage4_18;
   wire [19:0] stage4_19;
   wire [21:0] stage4_20;
   wire [26:0] stage4_21;
   wire [20:0] stage4_22;
   wire [23:0] stage4_23;
   wire [23:0] stage4_24;
   wire [19:0] stage4_25;
   wire [20:0] stage4_26;
   wire [20:0] stage4_27;
   wire [31:0] stage4_28;
   wire [23:0] stage4_29;
   wire [25:0] stage4_30;
   wire [16:0] stage4_31;
   wire [23:0] stage4_32;
   wire [33:0] stage4_33;
   wire [29:0] stage4_34;
   wire [23:0] stage4_35;
   wire [37:0] stage4_36;
   wire [15:0] stage4_37;
   wire [26:0] stage4_38;
   wire [22:0] stage4_39;
   wire [28:0] stage4_40;
   wire [23:0] stage4_41;
   wire [28:0] stage4_42;
   wire [22:0] stage4_43;
   wire [39:0] stage4_44;
   wire [25:0] stage4_45;
   wire [24:0] stage4_46;
   wire [25:0] stage4_47;
   wire [21:0] stage4_48;
   wire [27:0] stage4_49;
   wire [23:0] stage4_50;
   wire [26:0] stage4_51;
   wire [22:0] stage4_52;
   wire [28:0] stage4_53;
   wire [30:0] stage4_54;
   wire [28:0] stage4_55;
   wire [28:0] stage4_56;
   wire [24:0] stage4_57;
   wire [15:0] stage4_58;
   wire [15:0] stage4_59;
   wire [24:0] stage4_60;
   wire [28:0] stage4_61;
   wire [23:0] stage4_62;
   wire [17:0] stage4_63;
   wire [26:0] stage4_64;
   wire [22:0] stage4_65;
   wire [14:0] stage4_66;
   wire [16:0] stage4_67;
   wire [11:0] stage4_68;
   wire [2:0] stage4_69;
   wire [0:0] stage4_70;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [2:0] stage5_2;
   wire [7:0] stage5_3;
   wire [8:0] stage5_4;
   wire [20:0] stage5_5;
   wire [13:0] stage5_6;
   wire [10:0] stage5_7;
   wire [15:0] stage5_8;
   wire [12:0] stage5_9;
   wire [9:0] stage5_10;
   wire [19:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [14:0] stage5_14;
   wire [15:0] stage5_15;
   wire [13:0] stage5_16;
   wire [7:0] stage5_17;
   wire [13:0] stage5_18;
   wire [13:0] stage5_19;
   wire [7:0] stage5_20;
   wire [10:0] stage5_21;
   wire [14:0] stage5_22;
   wire [11:0] stage5_23;
   wire [8:0] stage5_24;
   wire [12:0] stage5_25;
   wire [16:0] stage5_26;
   wire [8:0] stage5_27;
   wire [11:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [11:0] stage5_31;
   wire [14:0] stage5_32;
   wire [8:0] stage5_33;
   wire [20:0] stage5_34;
   wire [8:0] stage5_35;
   wire [18:0] stage5_36;
   wire [10:0] stage5_37;
   wire [6:0] stage5_38;
   wire [10:0] stage5_39;
   wire [19:0] stage5_40;
   wire [8:0] stage5_41;
   wire [19:0] stage5_42;
   wire [7:0] stage5_43;
   wire [25:0] stage5_44;
   wire [9:0] stage5_45;
   wire [10:0] stage5_46;
   wire [12:0] stage5_47;
   wire [17:0] stage5_48;
   wire [16:0] stage5_49;
   wire [9:0] stage5_50;
   wire [9:0] stage5_51;
   wire [12:0] stage5_52;
   wire [11:0] stage5_53;
   wire [16:0] stage5_54;
   wire [17:0] stage5_55;
   wire [12:0] stage5_56;
   wire [8:0] stage5_57;
   wire [23:0] stage5_58;
   wire [5:0] stage5_59;
   wire [13:0] stage5_60;
   wire [9:0] stage5_61;
   wire [7:0] stage5_62;
   wire [10:0] stage5_63;
   wire [19:0] stage5_64;
   wire [5:0] stage5_65;
   wire [12:0] stage5_66;
   wire [7:0] stage5_67;
   wire [11:0] stage5_68;
   wire [2:0] stage5_69;
   wire [3:0] stage5_70;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [2:0] stage6_2;
   wire [3:0] stage6_3;
   wire [2:0] stage6_4;
   wire [6:0] stage6_5;
   wire [5:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [7:0] stage6_9;
   wire [4:0] stage6_10;
   wire [5:0] stage6_11;
   wire [7:0] stage6_12;
   wire [4:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [11:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [8:0] stage6_25;
   wire [4:0] stage6_26;
   wire [4:0] stage6_27;
   wire [3:0] stage6_28;
   wire [5:0] stage6_29;
   wire [7:0] stage6_30;
   wire [2:0] stage6_31;
   wire [5:0] stage6_32;
   wire [7:0] stage6_33;
   wire [5:0] stage6_34;
   wire [4:0] stage6_35;
   wire [7:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [4:0] stage6_39;
   wire [9:0] stage6_40;
   wire [10:0] stage6_41;
   wire [3:0] stage6_42;
   wire [4:0] stage6_43;
   wire [7:0] stage6_44;
   wire [6:0] stage6_45;
   wire [6:0] stage6_46;
   wire [3:0] stage6_47;
   wire [5:0] stage6_48;
   wire [9:0] stage6_49;
   wire [4:0] stage6_50;
   wire [4:0] stage6_51;
   wire [7:0] stage6_52;
   wire [3:0] stage6_53;
   wire [5:0] stage6_54;
   wire [5:0] stage6_55;
   wire [6:0] stage6_56;
   wire [6:0] stage6_57;
   wire [6:0] stage6_58;
   wire [4:0] stage6_59;
   wire [6:0] stage6_60;
   wire [5:0] stage6_61;
   wire [4:0] stage6_62;
   wire [2:0] stage6_63;
   wire [5:0] stage6_64;
   wire [9:0] stage6_65;
   wire [2:0] stage6_66;
   wire [4:0] stage6_67;
   wire [9:0] stage6_68;
   wire [2:0] stage6_69;
   wire [1:0] stage6_70;
   wire [1:0] stage6_71;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [2:0] stage7_2;
   wire [3:0] stage7_3;
   wire [0:0] stage7_4;
   wire [4:0] stage7_5;
   wire [1:0] stage7_6;
   wire [6:0] stage7_7;
   wire [0:0] stage7_8;
   wire [4:0] stage7_9;
   wire [3:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [6:0] stage7_13;
   wire [2:0] stage7_14;
   wire [1:0] stage7_15;
   wire [6:0] stage7_16;
   wire [2:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [0:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [6:0] stage7_23;
   wire [2:0] stage7_24;
   wire [5:0] stage7_25;
   wire [6:0] stage7_26;
   wire [0:0] stage7_27;
   wire [1:0] stage7_28;
   wire [2:0] stage7_29;
   wire [3:0] stage7_30;
   wire [1:0] stage7_31;
   wire [2:0] stage7_32;
   wire [2:0] stage7_33;
   wire [5:0] stage7_34;
   wire [6:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [2:0] stage7_38;
   wire [3:0] stage7_39;
   wire [1:0] stage7_40;
   wire [5:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [6:0] stage7_45;
   wire [6:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [5:0] stage7_49;
   wire [2:0] stage7_50;
   wire [5:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [4:0] stage7_54;
   wire [1:0] stage7_55;
   wire [5:0] stage7_56;
   wire [2:0] stage7_57;
   wire [1:0] stage7_58;
   wire [2:0] stage7_59;
   wire [4:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [4:0] stage7_63;
   wire [2:0] stage7_64;
   wire [11:0] stage7_65;
   wire [0:0] stage7_66;
   wire [0:0] stage7_67;
   wire [3:0] stage7_68;
   wire [2:0] stage7_69;
   wire [2:0] stage7_70;
   wire [2:0] stage7_71;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [1:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [0:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_2[7]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[8]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[9]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[10]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[11]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[12]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[13]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[14]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[15]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[16]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[17]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[18]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[19]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[20]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[21]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[22]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[23]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[24]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[25]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[26]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[27]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[28]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[29]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[30]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[31]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[32]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[33]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[34]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[35]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[36]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_2[37]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_2[38]},
      {stage0_3[31]},
      {stage1_4[31],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_2[39]},
      {stage0_3[32]},
      {stage1_4[32],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_2[40]},
      {stage0_3[33]},
      {stage1_4[33],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_2[41]},
      {stage0_3[34]},
      {stage1_4[34],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_2[42]},
      {stage0_3[35]},
      {stage1_4[35],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_2[43]},
      {stage0_3[36]},
      {stage1_4[36],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_2[44]},
      {stage0_3[37]},
      {stage1_4[37],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc1163_5 gpc45 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_2[45]},
      {stage0_3[38]},
      {stage1_4[38],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc1163_5 gpc46 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_2[46]},
      {stage0_3[39]},
      {stage1_4[39],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc1163_5 gpc47 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_2[47]},
      {stage0_3[40]},
      {stage1_4[40],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc1163_5 gpc48 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_2[48]},
      {stage0_3[41]},
      {stage1_4[41],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc1163_5 gpc49 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_2[49]},
      {stage0_3[42]},
      {stage1_4[42],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc1163_5 gpc50 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_2[50]},
      {stage0_3[43]},
      {stage1_4[43],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc1163_5 gpc51 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_2[51]},
      {stage0_3[44]},
      {stage1_4[44],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc1163_5 gpc52 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_2[52]},
      {stage0_3[45]},
      {stage1_4[45],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc1163_5 gpc53 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_2[53]},
      {stage0_3[46]},
      {stage1_4[46],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc1163_5 gpc54 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_2[54]},
      {stage0_3[47]},
      {stage1_4[47],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc1163_5 gpc55 (
      {stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_2[55]},
      {stage0_3[48]},
      {stage1_4[48],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc1163_5 gpc56 (
      {stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_2[56]},
      {stage0_3[49]},
      {stage1_4[49],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[50],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[51],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[52],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[53],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc615_5 gpc61 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_1[307]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[54],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc615_5 gpc62 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_1[308]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[55],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc615_5 gpc63 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_1[309]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[56],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc615_5 gpc64 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_1[310]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[57],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc615_5 gpc65 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247]},
      {stage0_1[311]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[58],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc615_5 gpc66 (
      {stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_1[312]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[59],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc615_5 gpc67 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_1[313]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[60],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc615_5 gpc68 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_1[314]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[61],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc615_5 gpc69 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_1[315]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[62],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc615_5 gpc70 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_1[316]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[63],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc615_5 gpc71 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277]},
      {stage0_1[317]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[64],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc615_5 gpc72 (
      {stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_1[318]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[65],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc615_5 gpc73 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_1[319]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[66],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc615_5 gpc74 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_1[320]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[67],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc615_5 gpc75 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_1[321]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[68],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc615_5 gpc76 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_1[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[69],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc615_5 gpc77 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307]},
      {stage0_1[323]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[70],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc615_5 gpc78 (
      {stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_1[324]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[71],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc615_5 gpc79 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_1[325]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[72],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc615_5 gpc80 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_1[326]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[73],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc615_5 gpc81 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_1[327]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[74],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc615_5 gpc82 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_1[328]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[75],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc615_5 gpc83 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337]},
      {stage0_1[329]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[76],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc615_5 gpc84 (
      {stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_1[330]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[77],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc615_5 gpc85 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_1[331]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[78],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc615_5 gpc86 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_1[332]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[79],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc615_5 gpc87 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_1[333]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[80],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc615_5 gpc88 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_1[334]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[81],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc615_5 gpc89 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367]},
      {stage0_1[335]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[82],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc615_5 gpc90 (
      {stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_1[336]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[83],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc615_5 gpc91 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_1[337]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[84],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc615_5 gpc92 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_1[338]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[85],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc615_5 gpc93 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_1[339]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[86],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc615_5 gpc94 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_1[340]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[87],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc615_5 gpc95 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397]},
      {stage0_1[341]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[88],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc615_5 gpc96 (
      {stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_1[342]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[89],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc615_5 gpc97 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_1[343]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[90],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc615_5 gpc98 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_1[344]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[91],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc615_5 gpc99 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_1[345]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[92],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc615_5 gpc100 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_1[346]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[93],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc615_5 gpc101 (
      {stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427]},
      {stage0_1[347]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[94],stage1_3[101],stage1_2[101],stage1_1[101],stage1_0[101]}
   );
   gpc615_5 gpc102 (
      {stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_1[348]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[95],stage1_3[102],stage1_2[102],stage1_1[102],stage1_0[102]}
   );
   gpc615_5 gpc103 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_1[349]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[96],stage1_3[103],stage1_2[103],stage1_1[103],stage1_0[103]}
   );
   gpc615_5 gpc104 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_1[350]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[97],stage1_3[104],stage1_2[104],stage1_1[104],stage1_0[104]}
   );
   gpc615_5 gpc105 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_1[351]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[98],stage1_3[105],stage1_2[105],stage1_1[105],stage1_0[105]}
   );
   gpc615_5 gpc106 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452]},
      {stage0_1[352]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[99],stage1_3[106],stage1_2[106],stage1_1[106],stage1_0[106]}
   );
   gpc615_5 gpc107 (
      {stage0_0[453], stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457]},
      {stage0_1[353]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[100],stage1_3[107],stage1_2[107],stage1_1[107],stage1_0[107]}
   );
   gpc615_5 gpc108 (
      {stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461], stage0_0[462]},
      {stage0_1[354]},
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage1_4[101],stage1_3[108],stage1_2[108],stage1_1[108],stage1_0[108]}
   );
   gpc615_5 gpc109 (
      {stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_1[355]},
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage1_4[102],stage1_3[109],stage1_2[109],stage1_1[109],stage1_0[109]}
   );
   gpc615_5 gpc110 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_1[356]},
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage1_4[103],stage1_3[110],stage1_2[110],stage1_1[110],stage1_0[110]}
   );
   gpc615_5 gpc111 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_1[357]},
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage1_4[104],stage1_3[111],stage1_2[111],stage1_1[111],stage1_0[111]}
   );
   gpc615_5 gpc112 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482]},
      {stage0_1[358]},
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage1_4[105],stage1_3[112],stage1_2[112],stage1_1[112],stage1_0[112]}
   );
   gpc615_5 gpc113 (
      {stage0_0[483], stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487]},
      {stage0_1[359]},
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage1_4[106],stage1_3[113],stage1_2[113],stage1_1[113],stage1_0[113]}
   );
   gpc615_5 gpc114 (
      {stage0_0[488], stage0_0[489], stage0_0[490], stage0_0[491], stage0_0[492]},
      {stage0_1[360]},
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage1_4[107],stage1_3[114],stage1_2[114],stage1_1[114],stage1_0[114]}
   );
   gpc615_5 gpc115 (
      {stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496], stage0_0[497]},
      {stage0_1[361]},
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage1_4[108],stage1_3[115],stage1_2[115],stage1_1[115],stage1_0[115]}
   );
   gpc615_5 gpc116 (
      {stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_1[362]},
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416]},
      {stage1_4[109],stage1_3[116],stage1_2[116],stage1_1[116],stage1_0[116]}
   );
   gpc615_5 gpc117 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507]},
      {stage0_1[363]},
      {stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage1_4[110],stage1_3[117],stage1_2[117],stage1_1[117],stage1_0[117]}
   );
   gpc615_5 gpc118 (
      {stage0_0[508], stage0_0[509], stage0_0[510], stage0_0[511], 1'b0},
      {stage0_1[364]},
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage1_4[111],stage1_3[118],stage1_2[118],stage1_1[118],stage1_0[118]}
   );
   gpc7_3 gpc119 (
      {stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc7_3 gpc120 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[0],stage1_4[112],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[1],stage1_4[113],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[2],stage1_4[114],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[3],stage1_4[115],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[4],stage1_4[116],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[5],stage1_4[117],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[6],stage1_4[118],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[7],stage1_4[119],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[8],stage1_4[120],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[9],stage1_4[121],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[10],stage1_4[122],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[11],stage1_4[123],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[12],stage1_4[124],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[13],stage1_4[125],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[14],stage1_4[126],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[15],stage1_4[127],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479], stage0_1[480]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[16],stage1_4[128],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc615_5 gpc138 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[17],stage1_4[129],stage1_3[138]}
   );
   gpc615_5 gpc139 (
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[18],stage1_4[130],stage1_3[139]}
   );
   gpc615_5 gpc140 (
      {stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[19],stage1_4[131],stage1_3[140]}
   );
   gpc615_5 gpc141 (
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[20],stage1_4[132],stage1_3[141]}
   );
   gpc615_5 gpc142 (
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[21],stage1_4[133],stage1_3[142]}
   );
   gpc615_5 gpc143 (
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181]},
      {stage0_4[5]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[5],stage1_5[22],stage1_4[134],stage1_3[143]}
   );
   gpc615_5 gpc144 (
      {stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage0_4[6]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[6],stage1_5[23],stage1_4[135],stage1_3[144]}
   );
   gpc615_5 gpc145 (
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191]},
      {stage0_4[7]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[7],stage1_5[24],stage1_4[136],stage1_3[145]}
   );
   gpc615_5 gpc146 (
      {stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage0_4[8]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[8],stage1_5[25],stage1_4[137],stage1_3[146]}
   );
   gpc615_5 gpc147 (
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage0_4[9]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[9],stage1_5[26],stage1_4[138],stage1_3[147]}
   );
   gpc615_5 gpc148 (
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage0_4[10]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[10],stage1_5[27],stage1_4[139],stage1_3[148]}
   );
   gpc615_5 gpc149 (
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211]},
      {stage0_4[11]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[11],stage1_5[28],stage1_4[140],stage1_3[149]}
   );
   gpc615_5 gpc150 (
      {stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage0_4[12]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[12],stage1_5[29],stage1_4[141],stage1_3[150]}
   );
   gpc615_5 gpc151 (
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221]},
      {stage0_4[13]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[13],stage1_5[30],stage1_4[142],stage1_3[151]}
   );
   gpc615_5 gpc152 (
      {stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage0_4[14]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[14],stage1_5[31],stage1_4[143],stage1_3[152]}
   );
   gpc615_5 gpc153 (
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage0_4[15]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[15],stage1_5[32],stage1_4[144],stage1_3[153]}
   );
   gpc615_5 gpc154 (
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage0_4[16]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[16],stage1_5[33],stage1_4[145],stage1_3[154]}
   );
   gpc615_5 gpc155 (
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241]},
      {stage0_4[17]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[17],stage1_5[34],stage1_4[146],stage1_3[155]}
   );
   gpc615_5 gpc156 (
      {stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage0_4[18]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[18],stage1_5[35],stage1_4[147],stage1_3[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251]},
      {stage0_4[19]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[19],stage1_5[36],stage1_4[148],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage0_4[20]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[20],stage1_5[37],stage1_4[149],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage0_4[21]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[21],stage1_5[38],stage1_4[150],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage0_4[22]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[22],stage1_5[39],stage1_4[151],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271]},
      {stage0_4[23]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[23],stage1_5[40],stage1_4[152],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage0_4[24]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[24],stage1_5[41],stage1_4[153],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281]},
      {stage0_4[25]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[25],stage1_5[42],stage1_4[154],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage0_4[26]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[26],stage1_5[43],stage1_4[155],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage0_4[27]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[27],stage1_5[44],stage1_4[156],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage0_4[28]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[28],stage1_5[45],stage1_4[157],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301]},
      {stage0_4[29]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[29],stage1_5[46],stage1_4[158],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage0_4[30]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[30],stage1_5[47],stage1_4[159],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311]},
      {stage0_4[31]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[31],stage1_5[48],stage1_4[160],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316]},
      {stage0_4[32]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[32],stage1_5[49],stage1_4[161],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage0_4[33]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[33],stage1_5[50],stage1_4[162],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage0_4[34]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[34],stage1_5[51],stage1_4[163],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331]},
      {stage0_4[35]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[35],stage1_5[52],stage1_4[164],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage0_4[36]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[36],stage1_5[53],stage1_4[165],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341]},
      {stage0_4[37]},
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage1_7[37],stage1_6[37],stage1_5[54],stage1_4[166],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346]},
      {stage0_4[38]},
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage1_7[38],stage1_6[38],stage1_5[55],stage1_4[167],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350], stage0_3[351]},
      {stage0_4[39]},
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage1_7[39],stage1_6[39],stage1_5[56],stage1_4[168],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage0_4[40]},
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage1_7[40],stage1_6[40],stage1_5[57],stage1_4[169],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361]},
      {stage0_4[41]},
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage1_7[41],stage1_6[41],stage1_5[58],stage1_4[170],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366]},
      {stage0_4[42]},
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage1_7[42],stage1_6[42],stage1_5[59],stage1_4[171],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370], stage0_3[371]},
      {stage0_4[43]},
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage1_7[43],stage1_6[43],stage1_5[60],stage1_4[172],stage1_3[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[44],stage1_6[44],stage1_5[61],stage1_4[173]}
   );
   gpc606_5 gpc183 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[45],stage1_6[45],stage1_5[62],stage1_4[174]}
   );
   gpc606_5 gpc184 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[46],stage1_6[46],stage1_5[63],stage1_4[175]}
   );
   gpc606_5 gpc185 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[47],stage1_6[47],stage1_5[64],stage1_4[176]}
   );
   gpc606_5 gpc186 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[48],stage1_6[48],stage1_5[65],stage1_4[177]}
   );
   gpc606_5 gpc187 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[49],stage1_6[49],stage1_5[66],stage1_4[178]}
   );
   gpc606_5 gpc188 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[50],stage1_6[50],stage1_5[67],stage1_4[179]}
   );
   gpc606_5 gpc189 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[51],stage1_6[51],stage1_5[68],stage1_4[180]}
   );
   gpc606_5 gpc190 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[52],stage1_6[52],stage1_5[69],stage1_4[181]}
   );
   gpc606_5 gpc191 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[53],stage1_6[53],stage1_5[70],stage1_4[182]}
   );
   gpc606_5 gpc192 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[54],stage1_6[54],stage1_5[71],stage1_4[183]}
   );
   gpc606_5 gpc193 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[55],stage1_6[55],stage1_5[72],stage1_4[184]}
   );
   gpc606_5 gpc194 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[56],stage1_6[56],stage1_5[73],stage1_4[185]}
   );
   gpc606_5 gpc195 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[57],stage1_6[57],stage1_5[74],stage1_4[186]}
   );
   gpc606_5 gpc196 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[58],stage1_6[58],stage1_5[75],stage1_4[187]}
   );
   gpc606_5 gpc197 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[59],stage1_6[59],stage1_5[76],stage1_4[188]}
   );
   gpc606_5 gpc198 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[60],stage1_6[60],stage1_5[77],stage1_4[189]}
   );
   gpc606_5 gpc199 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[61],stage1_6[61],stage1_5[78],stage1_4[190]}
   );
   gpc606_5 gpc200 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[62],stage1_6[62],stage1_5[79],stage1_4[191]}
   );
   gpc606_5 gpc201 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[63],stage1_6[63],stage1_5[80],stage1_4[192]}
   );
   gpc606_5 gpc202 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[64],stage1_6[64],stage1_5[81],stage1_4[193]}
   );
   gpc606_5 gpc203 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[65],stage1_6[65],stage1_5[82],stage1_4[194]}
   );
   gpc606_5 gpc204 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[66],stage1_6[66],stage1_5[83],stage1_4[195]}
   );
   gpc606_5 gpc205 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[67],stage1_6[67],stage1_5[84],stage1_4[196]}
   );
   gpc606_5 gpc206 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[68],stage1_6[68],stage1_5[85],stage1_4[197]}
   );
   gpc606_5 gpc207 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[69],stage1_6[69],stage1_5[86],stage1_4[198]}
   );
   gpc606_5 gpc208 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[70],stage1_6[70],stage1_5[87],stage1_4[199]}
   );
   gpc606_5 gpc209 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[71],stage1_6[71],stage1_5[88],stage1_4[200]}
   );
   gpc606_5 gpc210 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[72],stage1_6[72],stage1_5[89],stage1_4[201]}
   );
   gpc606_5 gpc211 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[73],stage1_6[73],stage1_5[90],stage1_4[202]}
   );
   gpc606_5 gpc212 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[74],stage1_6[74],stage1_5[91],stage1_4[203]}
   );
   gpc606_5 gpc213 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[75],stage1_6[75],stage1_5[92],stage1_4[204]}
   );
   gpc606_5 gpc214 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[76],stage1_6[76],stage1_5[93],stage1_4[205]}
   );
   gpc606_5 gpc215 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[77],stage1_6[77],stage1_5[94],stage1_4[206]}
   );
   gpc606_5 gpc216 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[78],stage1_6[78],stage1_5[95],stage1_4[207]}
   );
   gpc606_5 gpc217 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[79],stage1_6[79],stage1_5[96],stage1_4[208]}
   );
   gpc606_5 gpc218 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[80],stage1_6[80],stage1_5[97],stage1_4[209]}
   );
   gpc606_5 gpc219 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[81],stage1_6[81],stage1_5[98],stage1_4[210]}
   );
   gpc606_5 gpc220 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[82],stage1_6[82],stage1_5[99],stage1_4[211]}
   );
   gpc606_5 gpc221 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[83],stage1_6[83],stage1_5[100],stage1_4[212]}
   );
   gpc606_5 gpc222 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[84],stage1_6[84],stage1_5[101],stage1_4[213]}
   );
   gpc606_5 gpc223 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[85],stage1_6[85],stage1_5[102],stage1_4[214]}
   );
   gpc606_5 gpc224 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[86],stage1_6[86],stage1_5[103],stage1_4[215]}
   );
   gpc606_5 gpc225 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[87],stage1_6[87],stage1_5[104],stage1_4[216]}
   );
   gpc606_5 gpc226 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[88],stage1_6[88],stage1_5[105],stage1_4[217]}
   );
   gpc606_5 gpc227 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[89],stage1_6[89],stage1_5[106],stage1_4[218]}
   );
   gpc606_5 gpc228 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[90],stage1_6[90],stage1_5[107],stage1_4[219]}
   );
   gpc606_5 gpc229 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[91],stage1_6[91],stage1_5[108],stage1_4[220]}
   );
   gpc606_5 gpc230 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[92],stage1_6[92],stage1_5[109],stage1_4[221]}
   );
   gpc606_5 gpc231 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[93],stage1_6[93],stage1_5[110],stage1_4[222]}
   );
   gpc606_5 gpc232 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[94],stage1_6[94],stage1_5[111],stage1_4[223]}
   );
   gpc606_5 gpc233 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[95],stage1_6[95],stage1_5[112],stage1_4[224]}
   );
   gpc606_5 gpc234 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[96],stage1_6[96],stage1_5[113],stage1_4[225]}
   );
   gpc606_5 gpc235 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[97],stage1_6[97],stage1_5[114],stage1_4[226]}
   );
   gpc606_5 gpc236 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[98],stage1_6[98],stage1_5[115],stage1_4[227]}
   );
   gpc606_5 gpc237 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[99],stage1_6[99],stage1_5[116],stage1_4[228]}
   );
   gpc606_5 gpc238 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[100],stage1_6[100],stage1_5[117],stage1_4[229]}
   );
   gpc606_5 gpc239 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[101],stage1_6[101],stage1_5[118],stage1_4[230]}
   );
   gpc606_5 gpc240 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[102],stage1_6[102],stage1_5[119],stage1_4[231]}
   );
   gpc606_5 gpc241 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[103],stage1_6[103],stage1_5[120],stage1_4[232]}
   );
   gpc606_5 gpc242 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[104],stage1_6[104],stage1_5[121],stage1_4[233]}
   );
   gpc606_5 gpc243 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[105],stage1_6[105],stage1_5[122],stage1_4[234]}
   );
   gpc606_5 gpc244 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[106],stage1_6[106],stage1_5[123],stage1_4[235]}
   );
   gpc606_5 gpc245 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[107],stage1_6[107],stage1_5[124],stage1_4[236]}
   );
   gpc606_5 gpc246 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[108],stage1_6[108],stage1_5[125],stage1_4[237]}
   );
   gpc606_5 gpc247 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[109],stage1_6[109],stage1_5[126],stage1_4[238]}
   );
   gpc606_5 gpc248 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[110],stage1_6[110],stage1_5[127],stage1_4[239]}
   );
   gpc606_5 gpc249 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[111],stage1_6[111],stage1_5[128],stage1_4[240]}
   );
   gpc606_5 gpc250 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[112],stage1_6[112],stage1_5[129],stage1_4[241]}
   );
   gpc606_5 gpc251 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[113],stage1_6[113],stage1_5[130],stage1_4[242]}
   );
   gpc606_5 gpc252 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[114],stage1_6[114],stage1_5[131],stage1_4[243]}
   );
   gpc606_5 gpc253 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[115],stage1_6[115],stage1_5[132],stage1_4[244]}
   );
   gpc606_5 gpc254 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[116],stage1_6[116],stage1_5[133],stage1_4[245]}
   );
   gpc606_5 gpc255 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486], stage0_4[487]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[117],stage1_6[117],stage1_5[134],stage1_4[246]}
   );
   gpc606_5 gpc256 (
      {stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491], stage0_4[492], stage0_4[493]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[118],stage1_6[118],stage1_5[135],stage1_4[247]}
   );
   gpc606_5 gpc257 (
      {stage0_4[494], stage0_4[495], stage0_4[496], stage0_4[497], stage0_4[498], stage0_4[499]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[119],stage1_6[119],stage1_5[136],stage1_4[248]}
   );
   gpc606_5 gpc258 (
      {stage0_4[500], stage0_4[501], stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[120],stage1_6[120],stage1_5[137],stage1_4[249]}
   );
   gpc606_5 gpc259 (
      {stage0_4[506], stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage1_8[77],stage1_7[121],stage1_6[121],stage1_5[138],stage1_4[250]}
   );
   gpc606_5 gpc260 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[78],stage1_7[122],stage1_6[122],stage1_5[139]}
   );
   gpc606_5 gpc261 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[79],stage1_7[123],stage1_6[123],stage1_5[140]}
   );
   gpc606_5 gpc262 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[80],stage1_7[124],stage1_6[124],stage1_5[141]}
   );
   gpc606_5 gpc263 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[81],stage1_7[125],stage1_6[125],stage1_5[142]}
   );
   gpc606_5 gpc264 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[82],stage1_7[126],stage1_6[126],stage1_5[143]}
   );
   gpc606_5 gpc265 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[83],stage1_7[127],stage1_6[127],stage1_5[144]}
   );
   gpc606_5 gpc266 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[84],stage1_7[128],stage1_6[128],stage1_5[145]}
   );
   gpc606_5 gpc267 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[85],stage1_7[129],stage1_6[129],stage1_5[146]}
   );
   gpc606_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[86],stage1_7[130],stage1_6[130],stage1_5[147]}
   );
   gpc606_5 gpc269 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[87],stage1_7[131],stage1_6[131],stage1_5[148]}
   );
   gpc606_5 gpc270 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[88],stage1_7[132],stage1_6[132],stage1_5[149]}
   );
   gpc606_5 gpc271 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[89],stage1_7[133],stage1_6[133],stage1_5[150]}
   );
   gpc606_5 gpc272 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[90],stage1_7[134],stage1_6[134],stage1_5[151]}
   );
   gpc606_5 gpc273 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[91],stage1_7[135],stage1_6[135],stage1_5[152]}
   );
   gpc606_5 gpc274 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[92],stage1_7[136],stage1_6[136],stage1_5[153]}
   );
   gpc606_5 gpc275 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[93],stage1_7[137],stage1_6[137],stage1_5[154]}
   );
   gpc606_5 gpc276 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[94],stage1_7[138],stage1_6[138],stage1_5[155]}
   );
   gpc606_5 gpc277 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[95],stage1_7[139],stage1_6[139],stage1_5[156]}
   );
   gpc606_5 gpc278 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[96],stage1_7[140],stage1_6[140],stage1_5[157]}
   );
   gpc606_5 gpc279 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[97],stage1_7[141],stage1_6[141],stage1_5[158]}
   );
   gpc606_5 gpc280 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[98],stage1_7[142],stage1_6[142],stage1_5[159]}
   );
   gpc606_5 gpc281 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[99],stage1_7[143],stage1_6[143],stage1_5[160]}
   );
   gpc606_5 gpc282 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[100],stage1_7[144],stage1_6[144],stage1_5[161]}
   );
   gpc606_5 gpc283 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[101],stage1_7[145],stage1_6[145],stage1_5[162]}
   );
   gpc606_5 gpc284 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[102],stage1_7[146],stage1_6[146],stage1_5[163]}
   );
   gpc606_5 gpc285 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[103],stage1_7[147],stage1_6[147],stage1_5[164]}
   );
   gpc606_5 gpc286 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[104],stage1_7[148],stage1_6[148],stage1_5[165]}
   );
   gpc606_5 gpc287 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[105],stage1_7[149],stage1_6[149],stage1_5[166]}
   );
   gpc606_5 gpc288 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[106],stage1_7[150],stage1_6[150],stage1_5[167]}
   );
   gpc606_5 gpc289 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[107],stage1_7[151],stage1_6[151],stage1_5[168]}
   );
   gpc606_5 gpc290 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[108],stage1_7[152],stage1_6[152],stage1_5[169]}
   );
   gpc606_5 gpc291 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[109],stage1_7[153],stage1_6[153],stage1_5[170]}
   );
   gpc606_5 gpc292 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[110],stage1_7[154],stage1_6[154],stage1_5[171]}
   );
   gpc606_5 gpc293 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[111],stage1_7[155],stage1_6[155],stage1_5[172]}
   );
   gpc615_5 gpc294 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472]},
      {stage0_7[204]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[34],stage1_8[112],stage1_7[156],stage1_6[156]}
   );
   gpc615_5 gpc295 (
      {stage0_6[473], stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477]},
      {stage0_7[205]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[35],stage1_8[113],stage1_7[157],stage1_6[157]}
   );
   gpc615_5 gpc296 (
      {stage0_6[478], stage0_6[479], stage0_6[480], stage0_6[481], stage0_6[482]},
      {stage0_7[206]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[36],stage1_8[114],stage1_7[158],stage1_6[158]}
   );
   gpc615_5 gpc297 (
      {stage0_6[483], stage0_6[484], stage0_6[485], stage0_6[486], stage0_6[487]},
      {stage0_7[207]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[37],stage1_8[115],stage1_7[159],stage1_6[159]}
   );
   gpc615_5 gpc298 (
      {stage0_6[488], stage0_6[489], stage0_6[490], stage0_6[491], stage0_6[492]},
      {stage0_7[208]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[38],stage1_8[116],stage1_7[160],stage1_6[160]}
   );
   gpc615_5 gpc299 (
      {stage0_7[209], stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[39],stage1_8[117],stage1_7[161]}
   );
   gpc615_5 gpc300 (
      {stage0_7[214], stage0_7[215], stage0_7[216], stage0_7[217], stage0_7[218]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[40],stage1_8[118],stage1_7[162]}
   );
   gpc615_5 gpc301 (
      {stage0_7[219], stage0_7[220], stage0_7[221], stage0_7[222], stage0_7[223]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[41],stage1_8[119],stage1_7[163]}
   );
   gpc615_5 gpc302 (
      {stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227], stage0_7[228]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[42],stage1_8[120],stage1_7[164]}
   );
   gpc615_5 gpc303 (
      {stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[43],stage1_8[121],stage1_7[165]}
   );
   gpc615_5 gpc304 (
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[44],stage1_8[122],stage1_7[166]}
   );
   gpc615_5 gpc305 (
      {stage0_7[239], stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[45],stage1_8[123],stage1_7[167]}
   );
   gpc615_5 gpc306 (
      {stage0_7[244], stage0_7[245], stage0_7[246], stage0_7[247], stage0_7[248]},
      {stage0_8[37]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[12],stage1_9[46],stage1_8[124],stage1_7[168]}
   );
   gpc615_5 gpc307 (
      {stage0_7[249], stage0_7[250], stage0_7[251], stage0_7[252], stage0_7[253]},
      {stage0_8[38]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[13],stage1_9[47],stage1_8[125],stage1_7[169]}
   );
   gpc615_5 gpc308 (
      {stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257], stage0_7[258]},
      {stage0_8[39]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[14],stage1_9[48],stage1_8[126],stage1_7[170]}
   );
   gpc615_5 gpc309 (
      {stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage0_8[40]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[15],stage1_9[49],stage1_8[127],stage1_7[171]}
   );
   gpc615_5 gpc310 (
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268]},
      {stage0_8[41]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[16],stage1_9[50],stage1_8[128],stage1_7[172]}
   );
   gpc615_5 gpc311 (
      {stage0_7[269], stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273]},
      {stage0_8[42]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[17],stage1_9[51],stage1_8[129],stage1_7[173]}
   );
   gpc615_5 gpc312 (
      {stage0_7[274], stage0_7[275], stage0_7[276], stage0_7[277], stage0_7[278]},
      {stage0_8[43]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[18],stage1_9[52],stage1_8[130],stage1_7[174]}
   );
   gpc615_5 gpc313 (
      {stage0_7[279], stage0_7[280], stage0_7[281], stage0_7[282], stage0_7[283]},
      {stage0_8[44]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[19],stage1_9[53],stage1_8[131],stage1_7[175]}
   );
   gpc615_5 gpc314 (
      {stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287], stage0_7[288]},
      {stage0_8[45]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[20],stage1_9[54],stage1_8[132],stage1_7[176]}
   );
   gpc615_5 gpc315 (
      {stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage0_8[46]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[21],stage1_9[55],stage1_8[133],stage1_7[177]}
   );
   gpc615_5 gpc316 (
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298]},
      {stage0_8[47]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[22],stage1_9[56],stage1_8[134],stage1_7[178]}
   );
   gpc615_5 gpc317 (
      {stage0_7[299], stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303]},
      {stage0_8[48]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[23],stage1_9[57],stage1_8[135],stage1_7[179]}
   );
   gpc615_5 gpc318 (
      {stage0_7[304], stage0_7[305], stage0_7[306], stage0_7[307], stage0_7[308]},
      {stage0_8[49]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[24],stage1_9[58],stage1_8[136],stage1_7[180]}
   );
   gpc615_5 gpc319 (
      {stage0_7[309], stage0_7[310], stage0_7[311], stage0_7[312], stage0_7[313]},
      {stage0_8[50]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[25],stage1_9[59],stage1_8[137],stage1_7[181]}
   );
   gpc615_5 gpc320 (
      {stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317], stage0_7[318]},
      {stage0_8[51]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[26],stage1_9[60],stage1_8[138],stage1_7[182]}
   );
   gpc615_5 gpc321 (
      {stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage0_8[52]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[27],stage1_9[61],stage1_8[139],stage1_7[183]}
   );
   gpc615_5 gpc322 (
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328]},
      {stage0_8[53]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[28],stage1_9[62],stage1_8[140],stage1_7[184]}
   );
   gpc615_5 gpc323 (
      {stage0_7[329], stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333]},
      {stage0_8[54]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[29],stage1_9[63],stage1_8[141],stage1_7[185]}
   );
   gpc615_5 gpc324 (
      {stage0_7[334], stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338]},
      {stage0_8[55]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[30],stage1_9[64],stage1_8[142],stage1_7[186]}
   );
   gpc615_5 gpc325 (
      {stage0_7[339], stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343]},
      {stage0_8[56]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[31],stage1_9[65],stage1_8[143],stage1_7[187]}
   );
   gpc615_5 gpc326 (
      {stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348]},
      {stage0_8[57]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[32],stage1_9[66],stage1_8[144],stage1_7[188]}
   );
   gpc615_5 gpc327 (
      {stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage0_8[58]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[33],stage1_9[67],stage1_8[145],stage1_7[189]}
   );
   gpc615_5 gpc328 (
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358]},
      {stage0_8[59]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[34],stage1_9[68],stage1_8[146],stage1_7[190]}
   );
   gpc615_5 gpc329 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363]},
      {stage0_8[60]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[35],stage1_9[69],stage1_8[147],stage1_7[191]}
   );
   gpc606_5 gpc330 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[31],stage1_10[36],stage1_9[70],stage1_8[148]}
   );
   gpc606_5 gpc331 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[32],stage1_10[37],stage1_9[71],stage1_8[149]}
   );
   gpc606_5 gpc332 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[33],stage1_10[38],stage1_9[72],stage1_8[150]}
   );
   gpc606_5 gpc333 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[34],stage1_10[39],stage1_9[73],stage1_8[151]}
   );
   gpc606_5 gpc334 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[35],stage1_10[40],stage1_9[74],stage1_8[152]}
   );
   gpc606_5 gpc335 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[36],stage1_10[41],stage1_9[75],stage1_8[153]}
   );
   gpc606_5 gpc336 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[37],stage1_10[42],stage1_9[76],stage1_8[154]}
   );
   gpc606_5 gpc337 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[38],stage1_10[43],stage1_9[77],stage1_8[155]}
   );
   gpc606_5 gpc338 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[39],stage1_10[44],stage1_9[78],stage1_8[156]}
   );
   gpc606_5 gpc339 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[40],stage1_10[45],stage1_9[79],stage1_8[157]}
   );
   gpc606_5 gpc340 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[41],stage1_10[46],stage1_9[80],stage1_8[158]}
   );
   gpc606_5 gpc341 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[42],stage1_10[47],stage1_9[81],stage1_8[159]}
   );
   gpc606_5 gpc342 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[43],stage1_10[48],stage1_9[82],stage1_8[160]}
   );
   gpc606_5 gpc343 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[44],stage1_10[49],stage1_9[83],stage1_8[161]}
   );
   gpc606_5 gpc344 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[45],stage1_10[50],stage1_9[84],stage1_8[162]}
   );
   gpc606_5 gpc345 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[46],stage1_10[51],stage1_9[85],stage1_8[163]}
   );
   gpc606_5 gpc346 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[47],stage1_10[52],stage1_9[86],stage1_8[164]}
   );
   gpc606_5 gpc347 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[48],stage1_10[53],stage1_9[87],stage1_8[165]}
   );
   gpc606_5 gpc348 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[49],stage1_10[54],stage1_9[88],stage1_8[166]}
   );
   gpc606_5 gpc349 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[50],stage1_10[55],stage1_9[89],stage1_8[167]}
   );
   gpc606_5 gpc350 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[51],stage1_10[56],stage1_9[90],stage1_8[168]}
   );
   gpc606_5 gpc351 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[52],stage1_10[57],stage1_9[91],stage1_8[169]}
   );
   gpc606_5 gpc352 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[53],stage1_10[58],stage1_9[92],stage1_8[170]}
   );
   gpc606_5 gpc353 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[54],stage1_10[59],stage1_9[93],stage1_8[171]}
   );
   gpc606_5 gpc354 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[55],stage1_10[60],stage1_9[94],stage1_8[172]}
   );
   gpc606_5 gpc355 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[56],stage1_10[61],stage1_9[95],stage1_8[173]}
   );
   gpc606_5 gpc356 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[57],stage1_10[62],stage1_9[96],stage1_8[174]}
   );
   gpc606_5 gpc357 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[58],stage1_10[63],stage1_9[97],stage1_8[175]}
   );
   gpc606_5 gpc358 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[59],stage1_10[64],stage1_9[98],stage1_8[176]}
   );
   gpc606_5 gpc359 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[60],stage1_10[65],stage1_9[99],stage1_8[177]}
   );
   gpc606_5 gpc360 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[61],stage1_10[66],stage1_9[100],stage1_8[178]}
   );
   gpc606_5 gpc361 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[62],stage1_10[67],stage1_9[101],stage1_8[179]}
   );
   gpc606_5 gpc362 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[63],stage1_10[68],stage1_9[102],stage1_8[180]}
   );
   gpc606_5 gpc363 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[64],stage1_10[69],stage1_9[103],stage1_8[181]}
   );
   gpc606_5 gpc364 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[65],stage1_10[70],stage1_9[104],stage1_8[182]}
   );
   gpc606_5 gpc365 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[66],stage1_10[71],stage1_9[105],stage1_8[183]}
   );
   gpc606_5 gpc366 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[67],stage1_10[72],stage1_9[106],stage1_8[184]}
   );
   gpc606_5 gpc367 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[68],stage1_10[73],stage1_9[107],stage1_8[185]}
   );
   gpc606_5 gpc368 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[69],stage1_10[74],stage1_9[108],stage1_8[186]}
   );
   gpc606_5 gpc369 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[70],stage1_10[75],stage1_9[109],stage1_8[187]}
   );
   gpc606_5 gpc370 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[71],stage1_10[76],stage1_9[110],stage1_8[188]}
   );
   gpc606_5 gpc371 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[72],stage1_10[77],stage1_9[111],stage1_8[189]}
   );
   gpc606_5 gpc372 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[73],stage1_10[78],stage1_9[112],stage1_8[190]}
   );
   gpc606_5 gpc373 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[74],stage1_10[79],stage1_9[113],stage1_8[191]}
   );
   gpc606_5 gpc374 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[75],stage1_10[80],stage1_9[114],stage1_8[192]}
   );
   gpc606_5 gpc375 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[76],stage1_10[81],stage1_9[115],stage1_8[193]}
   );
   gpc606_5 gpc376 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[77],stage1_10[82],stage1_9[116],stage1_8[194]}
   );
   gpc606_5 gpc377 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[78],stage1_10[83],stage1_9[117],stage1_8[195]}
   );
   gpc606_5 gpc378 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[79],stage1_10[84],stage1_9[118],stage1_8[196]}
   );
   gpc606_5 gpc379 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[80],stage1_10[85],stage1_9[119],stage1_8[197]}
   );
   gpc606_5 gpc380 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[81],stage1_10[86],stage1_9[120],stage1_8[198]}
   );
   gpc606_5 gpc381 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[82],stage1_10[87],stage1_9[121],stage1_8[199]}
   );
   gpc606_5 gpc382 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[83],stage1_10[88],stage1_9[122],stage1_8[200]}
   );
   gpc606_5 gpc383 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[84],stage1_10[89],stage1_9[123],stage1_8[201]}
   );
   gpc606_5 gpc384 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[85],stage1_10[90],stage1_9[124],stage1_8[202]}
   );
   gpc606_5 gpc385 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[86],stage1_10[91],stage1_9[125],stage1_8[203]}
   );
   gpc606_5 gpc386 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[87],stage1_10[92],stage1_9[126],stage1_8[204]}
   );
   gpc606_5 gpc387 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[88],stage1_10[93],stage1_9[127],stage1_8[205]}
   );
   gpc606_5 gpc388 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[89],stage1_10[94],stage1_9[128],stage1_8[206]}
   );
   gpc606_5 gpc389 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[90],stage1_10[95],stage1_9[129],stage1_8[207]}
   );
   gpc606_5 gpc390 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[91],stage1_10[96],stage1_9[130],stage1_8[208]}
   );
   gpc606_5 gpc391 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[92],stage1_10[97],stage1_9[131],stage1_8[209]}
   );
   gpc606_5 gpc392 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[93],stage1_10[98],stage1_9[132],stage1_8[210]}
   );
   gpc606_5 gpc393 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[94],stage1_10[99],stage1_9[133],stage1_8[211]}
   );
   gpc606_5 gpc394 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[95],stage1_10[100],stage1_9[134],stage1_8[212]}
   );
   gpc606_5 gpc395 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[96],stage1_10[101],stage1_9[135],stage1_8[213]}
   );
   gpc606_5 gpc396 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[97],stage1_10[102],stage1_9[136],stage1_8[214]}
   );
   gpc606_5 gpc397 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[98],stage1_10[103],stage1_9[137],stage1_8[215]}
   );
   gpc606_5 gpc398 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[99],stage1_10[104],stage1_9[138],stage1_8[216]}
   );
   gpc606_5 gpc399 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[100],stage1_10[105],stage1_9[139],stage1_8[217]}
   );
   gpc606_5 gpc400 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[101],stage1_10[106],stage1_9[140],stage1_8[218]}
   );
   gpc606_5 gpc401 (
      {stage0_8[487], stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[102],stage1_10[107],stage1_9[141],stage1_8[219]}
   );
   gpc606_5 gpc402 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[72],stage1_11[103],stage1_10[108],stage1_9[142]}
   );
   gpc606_5 gpc403 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[73],stage1_11[104],stage1_10[109],stage1_9[143]}
   );
   gpc606_5 gpc404 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[74],stage1_11[105],stage1_10[110],stage1_9[144]}
   );
   gpc606_5 gpc405 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[75],stage1_11[106],stage1_10[111],stage1_9[145]}
   );
   gpc606_5 gpc406 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[76],stage1_11[107],stage1_10[112],stage1_9[146]}
   );
   gpc606_5 gpc407 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[77],stage1_11[108],stage1_10[113],stage1_9[147]}
   );
   gpc606_5 gpc408 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[78],stage1_11[109],stage1_10[114],stage1_9[148]}
   );
   gpc606_5 gpc409 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[79],stage1_11[110],stage1_10[115],stage1_9[149]}
   );
   gpc606_5 gpc410 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[80],stage1_11[111],stage1_10[116],stage1_9[150]}
   );
   gpc606_5 gpc411 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[81],stage1_11[112],stage1_10[117],stage1_9[151]}
   );
   gpc606_5 gpc412 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[82],stage1_11[113],stage1_10[118],stage1_9[152]}
   );
   gpc606_5 gpc413 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[83],stage1_11[114],stage1_10[119],stage1_9[153]}
   );
   gpc606_5 gpc414 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[84],stage1_11[115],stage1_10[120],stage1_9[154]}
   );
   gpc606_5 gpc415 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[85],stage1_11[116],stage1_10[121],stage1_9[155]}
   );
   gpc606_5 gpc416 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[86],stage1_11[117],stage1_10[122],stage1_9[156]}
   );
   gpc606_5 gpc417 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[87],stage1_11[118],stage1_10[123],stage1_9[157]}
   );
   gpc606_5 gpc418 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[88],stage1_11[119],stage1_10[124],stage1_9[158]}
   );
   gpc606_5 gpc419 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[89],stage1_11[120],stage1_10[125],stage1_9[159]}
   );
   gpc606_5 gpc420 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[90],stage1_11[121],stage1_10[126],stage1_9[160]}
   );
   gpc606_5 gpc421 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[91],stage1_11[122],stage1_10[127],stage1_9[161]}
   );
   gpc606_5 gpc422 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[92],stage1_11[123],stage1_10[128],stage1_9[162]}
   );
   gpc615_5 gpc423 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[126]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[21],stage1_12[93],stage1_11[124],stage1_10[129]}
   );
   gpc615_5 gpc424 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[127]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[22],stage1_12[94],stage1_11[125],stage1_10[130]}
   );
   gpc615_5 gpc425 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[128]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[23],stage1_12[95],stage1_11[126],stage1_10[131]}
   );
   gpc615_5 gpc426 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[129]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[24],stage1_12[96],stage1_11[127],stage1_10[132]}
   );
   gpc615_5 gpc427 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[130]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[25],stage1_12[97],stage1_11[128],stage1_10[133]}
   );
   gpc615_5 gpc428 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[131]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[26],stage1_12[98],stage1_11[129],stage1_10[134]}
   );
   gpc615_5 gpc429 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[132]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[27],stage1_12[99],stage1_11[130],stage1_10[135]}
   );
   gpc615_5 gpc430 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[133]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[28],stage1_12[100],stage1_11[131],stage1_10[136]}
   );
   gpc615_5 gpc431 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[134]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[29],stage1_12[101],stage1_11[132],stage1_10[137]}
   );
   gpc615_5 gpc432 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[135]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[30],stage1_12[102],stage1_11[133],stage1_10[138]}
   );
   gpc615_5 gpc433 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[136]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[31],stage1_12[103],stage1_11[134],stage1_10[139]}
   );
   gpc615_5 gpc434 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[137]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[32],stage1_12[104],stage1_11[135],stage1_10[140]}
   );
   gpc615_5 gpc435 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[138]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[33],stage1_12[105],stage1_11[136],stage1_10[141]}
   );
   gpc615_5 gpc436 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[139]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[34],stage1_12[106],stage1_11[137],stage1_10[142]}
   );
   gpc615_5 gpc437 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[84]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[14],stage1_13[35],stage1_12[107],stage1_11[138]}
   );
   gpc615_5 gpc438 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[85]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[15],stage1_13[36],stage1_12[108],stage1_11[139]}
   );
   gpc615_5 gpc439 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[86]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[16],stage1_13[37],stage1_12[109],stage1_11[140]}
   );
   gpc615_5 gpc440 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[87]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[17],stage1_13[38],stage1_12[110],stage1_11[141]}
   );
   gpc615_5 gpc441 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[88]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[18],stage1_13[39],stage1_12[111],stage1_11[142]}
   );
   gpc615_5 gpc442 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[89]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[19],stage1_13[40],stage1_12[112],stage1_11[143]}
   );
   gpc615_5 gpc443 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[90]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[20],stage1_13[41],stage1_12[113],stage1_11[144]}
   );
   gpc615_5 gpc444 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[91]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[21],stage1_13[42],stage1_12[114],stage1_11[145]}
   );
   gpc615_5 gpc445 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[92]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[22],stage1_13[43],stage1_12[115],stage1_11[146]}
   );
   gpc615_5 gpc446 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[93]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[23],stage1_13[44],stage1_12[116],stage1_11[147]}
   );
   gpc615_5 gpc447 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[94]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[24],stage1_13[45],stage1_12[117],stage1_11[148]}
   );
   gpc615_5 gpc448 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[95]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[25],stage1_13[46],stage1_12[118],stage1_11[149]}
   );
   gpc615_5 gpc449 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[96]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[26],stage1_13[47],stage1_12[119],stage1_11[150]}
   );
   gpc615_5 gpc450 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[97]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[27],stage1_13[48],stage1_12[120],stage1_11[151]}
   );
   gpc615_5 gpc451 (
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214]},
      {stage0_12[98]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[28],stage1_13[49],stage1_12[121],stage1_11[152]}
   );
   gpc615_5 gpc452 (
      {stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage0_12[99]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[29],stage1_13[50],stage1_12[122],stage1_11[153]}
   );
   gpc615_5 gpc453 (
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224]},
      {stage0_12[100]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[30],stage1_13[51],stage1_12[123],stage1_11[154]}
   );
   gpc615_5 gpc454 (
      {stage0_11[225], stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229]},
      {stage0_12[101]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[31],stage1_13[52],stage1_12[124],stage1_11[155]}
   );
   gpc615_5 gpc455 (
      {stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233], stage0_11[234]},
      {stage0_12[102]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[32],stage1_13[53],stage1_12[125],stage1_11[156]}
   );
   gpc615_5 gpc456 (
      {stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage0_12[103]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[33],stage1_13[54],stage1_12[126],stage1_11[157]}
   );
   gpc615_5 gpc457 (
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244]},
      {stage0_12[104]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[34],stage1_13[55],stage1_12[127],stage1_11[158]}
   );
   gpc615_5 gpc458 (
      {stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage0_12[105]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[35],stage1_13[56],stage1_12[128],stage1_11[159]}
   );
   gpc615_5 gpc459 (
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254]},
      {stage0_12[106]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[36],stage1_13[57],stage1_12[129],stage1_11[160]}
   );
   gpc615_5 gpc460 (
      {stage0_11[255], stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259]},
      {stage0_12[107]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[37],stage1_13[58],stage1_12[130],stage1_11[161]}
   );
   gpc615_5 gpc461 (
      {stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263], stage0_11[264]},
      {stage0_12[108]},
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage1_15[24],stage1_14[38],stage1_13[59],stage1_12[131],stage1_11[162]}
   );
   gpc615_5 gpc462 (
      {stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage0_12[109]},
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage1_15[25],stage1_14[39],stage1_13[60],stage1_12[132],stage1_11[163]}
   );
   gpc615_5 gpc463 (
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274]},
      {stage0_12[110]},
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage1_15[26],stage1_14[40],stage1_13[61],stage1_12[133],stage1_11[164]}
   );
   gpc615_5 gpc464 (
      {stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage0_12[111]},
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage1_15[27],stage1_14[41],stage1_13[62],stage1_12[134],stage1_11[165]}
   );
   gpc615_5 gpc465 (
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[112]},
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage1_15[28],stage1_14[42],stage1_13[63],stage1_12[135],stage1_11[166]}
   );
   gpc615_5 gpc466 (
      {stage0_11[285], stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289]},
      {stage0_12[113]},
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage1_15[29],stage1_14[43],stage1_13[64],stage1_12[136],stage1_11[167]}
   );
   gpc615_5 gpc467 (
      {stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293], stage0_11[294]},
      {stage0_12[114]},
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage1_15[30],stage1_14[44],stage1_13[65],stage1_12[137],stage1_11[168]}
   );
   gpc615_5 gpc468 (
      {stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage0_12[115]},
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage1_15[31],stage1_14[45],stage1_13[66],stage1_12[138],stage1_11[169]}
   );
   gpc615_5 gpc469 (
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304]},
      {stage0_12[116]},
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage1_15[32],stage1_14[46],stage1_13[67],stage1_12[139],stage1_11[170]}
   );
   gpc615_5 gpc470 (
      {stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage0_12[117]},
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage1_15[33],stage1_14[47],stage1_13[68],stage1_12[140],stage1_11[171]}
   );
   gpc615_5 gpc471 (
      {stage0_11[310], stage0_11[311], stage0_11[312], stage0_11[313], stage0_11[314]},
      {stage0_12[118]},
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage1_15[34],stage1_14[48],stage1_13[69],stage1_12[141],stage1_11[172]}
   );
   gpc615_5 gpc472 (
      {stage0_11[315], stage0_11[316], stage0_11[317], stage0_11[318], stage0_11[319]},
      {stage0_12[119]},
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage1_15[35],stage1_14[49],stage1_13[70],stage1_12[142],stage1_11[173]}
   );
   gpc615_5 gpc473 (
      {stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323], stage0_11[324]},
      {stage0_12[120]},
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage1_15[36],stage1_14[50],stage1_13[71],stage1_12[143],stage1_11[174]}
   );
   gpc615_5 gpc474 (
      {stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage0_12[121]},
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage1_15[37],stage1_14[51],stage1_13[72],stage1_12[144],stage1_11[175]}
   );
   gpc615_5 gpc475 (
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334]},
      {stage0_12[122]},
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage1_15[38],stage1_14[52],stage1_13[73],stage1_12[145],stage1_11[176]}
   );
   gpc615_5 gpc476 (
      {stage0_11[335], stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339]},
      {stage0_12[123]},
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage1_15[39],stage1_14[53],stage1_13[74],stage1_12[146],stage1_11[177]}
   );
   gpc615_5 gpc477 (
      {stage0_11[340], stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344]},
      {stage0_12[124]},
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage1_15[40],stage1_14[54],stage1_13[75],stage1_12[147],stage1_11[178]}
   );
   gpc615_5 gpc478 (
      {stage0_11[345], stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349]},
      {stage0_12[125]},
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage1_15[41],stage1_14[55],stage1_13[76],stage1_12[148],stage1_11[179]}
   );
   gpc615_5 gpc479 (
      {stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354]},
      {stage0_12[126]},
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage1_15[42],stage1_14[56],stage1_13[77],stage1_12[149],stage1_11[180]}
   );
   gpc615_5 gpc480 (
      {stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage0_12[127]},
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage1_15[43],stage1_14[57],stage1_13[78],stage1_12[150],stage1_11[181]}
   );
   gpc615_5 gpc481 (
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364]},
      {stage0_12[128]},
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage1_15[44],stage1_14[58],stage1_13[79],stage1_12[151],stage1_11[182]}
   );
   gpc615_5 gpc482 (
      {stage0_11[365], stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369]},
      {stage0_12[129]},
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage1_15[45],stage1_14[59],stage1_13[80],stage1_12[152],stage1_11[183]}
   );
   gpc615_5 gpc483 (
      {stage0_11[370], stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374]},
      {stage0_12[130]},
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage1_15[46],stage1_14[60],stage1_13[81],stage1_12[153],stage1_11[184]}
   );
   gpc615_5 gpc484 (
      {stage0_11[375], stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379]},
      {stage0_12[131]},
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage1_15[47],stage1_14[61],stage1_13[82],stage1_12[154],stage1_11[185]}
   );
   gpc606_5 gpc485 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[48],stage1_14[62],stage1_13[83],stage1_12[155]}
   );
   gpc606_5 gpc486 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[49],stage1_14[63],stage1_13[84],stage1_12[156]}
   );
   gpc606_5 gpc487 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[50],stage1_14[64],stage1_13[85],stage1_12[157]}
   );
   gpc606_5 gpc488 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[51],stage1_14[65],stage1_13[86],stage1_12[158]}
   );
   gpc606_5 gpc489 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[52],stage1_14[66],stage1_13[87],stage1_12[159]}
   );
   gpc606_5 gpc490 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[53],stage1_14[67],stage1_13[88],stage1_12[160]}
   );
   gpc606_5 gpc491 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[54],stage1_14[68],stage1_13[89],stage1_12[161]}
   );
   gpc606_5 gpc492 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[55],stage1_14[69],stage1_13[90],stage1_12[162]}
   );
   gpc606_5 gpc493 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[56],stage1_14[70],stage1_13[91],stage1_12[163]}
   );
   gpc606_5 gpc494 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[57],stage1_14[71],stage1_13[92],stage1_12[164]}
   );
   gpc606_5 gpc495 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[58],stage1_14[72],stage1_13[93],stage1_12[165]}
   );
   gpc606_5 gpc496 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[59],stage1_14[73],stage1_13[94],stage1_12[166]}
   );
   gpc606_5 gpc497 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[60],stage1_14[74],stage1_13[95],stage1_12[167]}
   );
   gpc606_5 gpc498 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[61],stage1_14[75],stage1_13[96],stage1_12[168]}
   );
   gpc606_5 gpc499 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[62],stage1_14[76],stage1_13[97],stage1_12[169]}
   );
   gpc606_5 gpc500 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[63],stage1_14[77],stage1_13[98],stage1_12[170]}
   );
   gpc606_5 gpc501 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[64],stage1_14[78],stage1_13[99],stage1_12[171]}
   );
   gpc606_5 gpc502 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[65],stage1_14[79],stage1_13[100],stage1_12[172]}
   );
   gpc606_5 gpc503 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[66],stage1_14[80],stage1_13[101],stage1_12[173]}
   );
   gpc606_5 gpc504 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[67],stage1_14[81],stage1_13[102],stage1_12[174]}
   );
   gpc606_5 gpc505 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[68],stage1_14[82],stage1_13[103],stage1_12[175]}
   );
   gpc606_5 gpc506 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[69],stage1_14[83],stage1_13[104],stage1_12[176]}
   );
   gpc606_5 gpc507 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[70],stage1_14[84],stage1_13[105],stage1_12[177]}
   );
   gpc606_5 gpc508 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[71],stage1_14[85],stage1_13[106],stage1_12[178]}
   );
   gpc606_5 gpc509 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[72],stage1_14[86],stage1_13[107],stage1_12[179]}
   );
   gpc606_5 gpc510 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[73],stage1_14[87],stage1_13[108],stage1_12[180]}
   );
   gpc606_5 gpc511 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[74],stage1_14[88],stage1_13[109],stage1_12[181]}
   );
   gpc606_5 gpc512 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[75],stage1_14[89],stage1_13[110],stage1_12[182]}
   );
   gpc606_5 gpc513 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[76],stage1_14[90],stage1_13[111],stage1_12[183]}
   );
   gpc606_5 gpc514 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[77],stage1_14[91],stage1_13[112],stage1_12[184]}
   );
   gpc606_5 gpc515 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[78],stage1_14[92],stage1_13[113],stage1_12[185]}
   );
   gpc606_5 gpc516 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[79],stage1_14[93],stage1_13[114],stage1_12[186]}
   );
   gpc606_5 gpc517 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[80],stage1_14[94],stage1_13[115],stage1_12[187]}
   );
   gpc606_5 gpc518 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[81],stage1_14[95],stage1_13[116],stage1_12[188]}
   );
   gpc606_5 gpc519 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[82],stage1_14[96],stage1_13[117],stage1_12[189]}
   );
   gpc606_5 gpc520 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[83],stage1_14[97],stage1_13[118],stage1_12[190]}
   );
   gpc606_5 gpc521 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[84],stage1_14[98],stage1_13[119],stage1_12[191]}
   );
   gpc606_5 gpc522 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[85],stage1_14[99],stage1_13[120],stage1_12[192]}
   );
   gpc606_5 gpc523 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[86],stage1_14[100],stage1_13[121],stage1_12[193]}
   );
   gpc606_5 gpc524 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[87],stage1_14[101],stage1_13[122],stage1_12[194]}
   );
   gpc606_5 gpc525 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[88],stage1_14[102],stage1_13[123],stage1_12[195]}
   );
   gpc606_5 gpc526 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[89],stage1_14[103],stage1_13[124],stage1_12[196]}
   );
   gpc606_5 gpc527 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[90],stage1_14[104],stage1_13[125],stage1_12[197]}
   );
   gpc606_5 gpc528 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[91],stage1_14[105],stage1_13[126],stage1_12[198]}
   );
   gpc606_5 gpc529 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[92],stage1_14[106],stage1_13[127],stage1_12[199]}
   );
   gpc606_5 gpc530 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[93],stage1_14[107],stage1_13[128],stage1_12[200]}
   );
   gpc606_5 gpc531 (
      {stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[94],stage1_14[108],stage1_13[129],stage1_12[201]}
   );
   gpc606_5 gpc532 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[95],stage1_14[109],stage1_13[130],stage1_12[202]}
   );
   gpc606_5 gpc533 (
      {stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[96],stage1_14[110],stage1_13[131],stage1_12[203]}
   );
   gpc606_5 gpc534 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[97],stage1_14[111],stage1_13[132],stage1_12[204]}
   );
   gpc606_5 gpc535 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[98],stage1_14[112],stage1_13[133],stage1_12[205]}
   );
   gpc606_5 gpc536 (
      {stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[99],stage1_14[113],stage1_13[134],stage1_12[206]}
   );
   gpc606_5 gpc537 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[100],stage1_14[114],stage1_13[135],stage1_12[207]}
   );
   gpc606_5 gpc538 (
      {stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[101],stage1_14[115],stage1_13[136],stage1_12[208]}
   );
   gpc606_5 gpc539 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[102],stage1_14[116],stage1_13[137],stage1_12[209]}
   );
   gpc606_5 gpc540 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[103],stage1_14[117],stage1_13[138],stage1_12[210]}
   );
   gpc606_5 gpc541 (
      {stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[104],stage1_14[118],stage1_13[139],stage1_12[211]}
   );
   gpc606_5 gpc542 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[105],stage1_14[119],stage1_13[140],stage1_12[212]}
   );
   gpc606_5 gpc543 (
      {stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[106],stage1_14[120],stage1_13[141],stage1_12[213]}
   );
   gpc606_5 gpc544 (
      {stage0_12[486], stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[107],stage1_14[121],stage1_13[142],stage1_12[214]}
   );
   gpc606_5 gpc545 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496], stage0_12[497]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[108],stage1_14[122],stage1_13[143],stage1_12[215]}
   );
   gpc606_5 gpc546 (
      {stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501], stage0_12[502], stage0_12[503]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[109],stage1_14[123],stage1_13[144],stage1_12[216]}
   );
   gpc606_5 gpc547 (
      {stage0_12[504], stage0_12[505], stage0_12[506], stage0_12[507], stage0_12[508], stage0_12[509]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[110],stage1_14[124],stage1_13[145],stage1_12[217]}
   );
   gpc606_5 gpc548 (
      {stage0_12[510], stage0_12[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage1_16[63],stage1_15[111],stage1_14[125],stage1_13[146],stage1_12[218]}
   );
   gpc606_5 gpc549 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[64],stage1_15[112],stage1_14[126],stage1_13[147]}
   );
   gpc606_5 gpc550 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[65],stage1_15[113],stage1_14[127],stage1_13[148]}
   );
   gpc606_5 gpc551 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[66],stage1_15[114],stage1_14[128],stage1_13[149]}
   );
   gpc606_5 gpc552 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[67],stage1_15[115],stage1_14[129],stage1_13[150]}
   );
   gpc606_5 gpc553 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[68],stage1_15[116],stage1_14[130],stage1_13[151]}
   );
   gpc606_5 gpc554 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[69],stage1_15[117],stage1_14[131],stage1_13[152]}
   );
   gpc606_5 gpc555 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[70],stage1_15[118],stage1_14[132],stage1_13[153]}
   );
   gpc606_5 gpc556 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[71],stage1_15[119],stage1_14[133],stage1_13[154]}
   );
   gpc606_5 gpc557 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[72],stage1_15[120],stage1_14[134],stage1_13[155]}
   );
   gpc606_5 gpc558 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[73],stage1_15[121],stage1_14[135],stage1_13[156]}
   );
   gpc606_5 gpc559 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[74],stage1_15[122],stage1_14[136],stage1_13[157]}
   );
   gpc606_5 gpc560 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[75],stage1_15[123],stage1_14[137],stage1_13[158]}
   );
   gpc606_5 gpc561 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[76],stage1_15[124],stage1_14[138],stage1_13[159]}
   );
   gpc606_5 gpc562 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[77],stage1_15[125],stage1_14[139],stage1_13[160]}
   );
   gpc606_5 gpc563 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[78],stage1_15[126],stage1_14[140],stage1_13[161]}
   );
   gpc606_5 gpc564 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[79],stage1_15[127],stage1_14[141],stage1_13[162]}
   );
   gpc606_5 gpc565 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[80],stage1_15[128],stage1_14[142],stage1_13[163]}
   );
   gpc606_5 gpc566 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[81],stage1_15[129],stage1_14[143],stage1_13[164]}
   );
   gpc606_5 gpc567 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[82],stage1_15[130],stage1_14[144],stage1_13[165]}
   );
   gpc606_5 gpc568 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[83],stage1_15[131],stage1_14[145],stage1_13[166]}
   );
   gpc606_5 gpc569 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[84],stage1_15[132],stage1_14[146],stage1_13[167]}
   );
   gpc606_5 gpc570 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[85],stage1_15[133],stage1_14[147],stage1_13[168]}
   );
   gpc606_5 gpc571 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[86],stage1_15[134],stage1_14[148],stage1_13[169]}
   );
   gpc606_5 gpc572 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[87],stage1_15[135],stage1_14[149],stage1_13[170]}
   );
   gpc606_5 gpc573 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[88],stage1_15[136],stage1_14[150],stage1_13[171]}
   );
   gpc606_5 gpc574 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[89],stage1_15[137],stage1_14[151],stage1_13[172]}
   );
   gpc606_5 gpc575 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[90],stage1_15[138],stage1_14[152],stage1_13[173]}
   );
   gpc606_5 gpc576 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[91],stage1_15[139],stage1_14[153],stage1_13[174]}
   );
   gpc606_5 gpc577 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[92],stage1_15[140],stage1_14[154],stage1_13[175]}
   );
   gpc606_5 gpc578 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466], stage0_13[467]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[93],stage1_15[141],stage1_14[155],stage1_13[176]}
   );
   gpc606_5 gpc579 (
      {stage0_13[468], stage0_13[469], stage0_13[470], stage0_13[471], stage0_13[472], stage0_13[473]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[94],stage1_15[142],stage1_14[156],stage1_13[177]}
   );
   gpc606_5 gpc580 (
      {stage0_13[474], stage0_13[475], stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[95],stage1_15[143],stage1_14[157],stage1_13[178]}
   );
   gpc606_5 gpc581 (
      {stage0_13[480], stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[96],stage1_15[144],stage1_14[158],stage1_13[179]}
   );
   gpc606_5 gpc582 (
      {stage0_13[486], stage0_13[487], stage0_13[488], stage0_13[489], stage0_13[490], stage0_13[491]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[97],stage1_15[145],stage1_14[159],stage1_13[180]}
   );
   gpc606_5 gpc583 (
      {stage0_13[492], stage0_13[493], stage0_13[494], stage0_13[495], stage0_13[496], stage0_13[497]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[98],stage1_15[146],stage1_14[160],stage1_13[181]}
   );
   gpc606_5 gpc584 (
      {stage0_13[498], stage0_13[499], stage0_13[500], stage0_13[501], stage0_13[502], stage0_13[503]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[99],stage1_15[147],stage1_14[161],stage1_13[182]}
   );
   gpc606_5 gpc585 (
      {stage0_13[504], stage0_13[505], stage0_13[506], stage0_13[507], stage0_13[508], stage0_13[509]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[100],stage1_15[148],stage1_14[162],stage1_13[183]}
   );
   gpc606_5 gpc586 (
      {stage0_13[510], stage0_13[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[101],stage1_15[149],stage1_14[163],stage1_13[184]}
   );
   gpc615_5 gpc587 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388]},
      {stage0_15[228]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[38],stage1_16[102],stage1_15[150],stage1_14[164]}
   );
   gpc615_5 gpc588 (
      {stage0_14[389], stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393]},
      {stage0_15[229]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[39],stage1_16[103],stage1_15[151],stage1_14[165]}
   );
   gpc615_5 gpc589 (
      {stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397], stage0_14[398]},
      {stage0_15[230]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[40],stage1_16[104],stage1_15[152],stage1_14[166]}
   );
   gpc615_5 gpc590 (
      {stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage0_15[231]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[41],stage1_16[105],stage1_15[153],stage1_14[167]}
   );
   gpc615_5 gpc591 (
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408]},
      {stage0_15[232]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[42],stage1_16[106],stage1_15[154],stage1_14[168]}
   );
   gpc615_5 gpc592 (
      {stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_15[233]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[43],stage1_16[107],stage1_15[155],stage1_14[169]}
   );
   gpc615_5 gpc593 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_15[234]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[44],stage1_16[108],stage1_15[156],stage1_14[170]}
   );
   gpc615_5 gpc594 (
      {stage0_14[419], stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423]},
      {stage0_15[235]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[45],stage1_16[109],stage1_15[157],stage1_14[171]}
   );
   gpc615_5 gpc595 (
      {stage0_14[424], stage0_14[425], stage0_14[426], stage0_14[427], stage0_14[428]},
      {stage0_15[236]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[46],stage1_16[110],stage1_15[158],stage1_14[172]}
   );
   gpc615_5 gpc596 (
      {stage0_15[237], stage0_15[238], stage0_15[239], stage0_15[240], stage0_15[241]},
      {stage0_16[54]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[9],stage1_17[47],stage1_16[111],stage1_15[159]}
   );
   gpc615_5 gpc597 (
      {stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245], stage0_15[246]},
      {stage0_16[55]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[10],stage1_17[48],stage1_16[112],stage1_15[160]}
   );
   gpc615_5 gpc598 (
      {stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage0_16[56]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[11],stage1_17[49],stage1_16[113],stage1_15[161]}
   );
   gpc615_5 gpc599 (
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256]},
      {stage0_16[57]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[12],stage1_17[50],stage1_16[114],stage1_15[162]}
   );
   gpc615_5 gpc600 (
      {stage0_15[257], stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261]},
      {stage0_16[58]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[13],stage1_17[51],stage1_16[115],stage1_15[163]}
   );
   gpc615_5 gpc601 (
      {stage0_15[262], stage0_15[263], stage0_15[264], stage0_15[265], stage0_15[266]},
      {stage0_16[59]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[14],stage1_17[52],stage1_16[116],stage1_15[164]}
   );
   gpc615_5 gpc602 (
      {stage0_15[267], stage0_15[268], stage0_15[269], stage0_15[270], stage0_15[271]},
      {stage0_16[60]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[15],stage1_17[53],stage1_16[117],stage1_15[165]}
   );
   gpc615_5 gpc603 (
      {stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275], stage0_15[276]},
      {stage0_16[61]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[16],stage1_17[54],stage1_16[118],stage1_15[166]}
   );
   gpc615_5 gpc604 (
      {stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage0_16[62]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[17],stage1_17[55],stage1_16[119],stage1_15[167]}
   );
   gpc615_5 gpc605 (
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286]},
      {stage0_16[63]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[18],stage1_17[56],stage1_16[120],stage1_15[168]}
   );
   gpc615_5 gpc606 (
      {stage0_15[287], stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291]},
      {stage0_16[64]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[19],stage1_17[57],stage1_16[121],stage1_15[169]}
   );
   gpc615_5 gpc607 (
      {stage0_15[292], stage0_15[293], stage0_15[294], stage0_15[295], stage0_15[296]},
      {stage0_16[65]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[20],stage1_17[58],stage1_16[122],stage1_15[170]}
   );
   gpc615_5 gpc608 (
      {stage0_15[297], stage0_15[298], stage0_15[299], stage0_15[300], stage0_15[301]},
      {stage0_16[66]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[21],stage1_17[59],stage1_16[123],stage1_15[171]}
   );
   gpc615_5 gpc609 (
      {stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305], stage0_15[306]},
      {stage0_16[67]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[22],stage1_17[60],stage1_16[124],stage1_15[172]}
   );
   gpc615_5 gpc610 (
      {stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage0_16[68]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[23],stage1_17[61],stage1_16[125],stage1_15[173]}
   );
   gpc615_5 gpc611 (
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316]},
      {stage0_16[69]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[24],stage1_17[62],stage1_16[126],stage1_15[174]}
   );
   gpc615_5 gpc612 (
      {stage0_15[317], stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321]},
      {stage0_16[70]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[25],stage1_17[63],stage1_16[127],stage1_15[175]}
   );
   gpc615_5 gpc613 (
      {stage0_15[322], stage0_15[323], stage0_15[324], stage0_15[325], stage0_15[326]},
      {stage0_16[71]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[26],stage1_17[64],stage1_16[128],stage1_15[176]}
   );
   gpc615_5 gpc614 (
      {stage0_15[327], stage0_15[328], stage0_15[329], stage0_15[330], stage0_15[331]},
      {stage0_16[72]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[27],stage1_17[65],stage1_16[129],stage1_15[177]}
   );
   gpc615_5 gpc615 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336]},
      {stage0_16[73]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[28],stage1_17[66],stage1_16[130],stage1_15[178]}
   );
   gpc615_5 gpc616 (
      {stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage0_16[74]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[29],stage1_17[67],stage1_16[131],stage1_15[179]}
   );
   gpc615_5 gpc617 (
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346]},
      {stage0_16[75]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[30],stage1_17[68],stage1_16[132],stage1_15[180]}
   );
   gpc615_5 gpc618 (
      {stage0_15[347], stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351]},
      {stage0_16[76]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[31],stage1_17[69],stage1_16[133],stage1_15[181]}
   );
   gpc615_5 gpc619 (
      {stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355], stage0_15[356]},
      {stage0_16[77]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[32],stage1_17[70],stage1_16[134],stage1_15[182]}
   );
   gpc615_5 gpc620 (
      {stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360], stage0_15[361]},
      {stage0_16[78]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[33],stage1_17[71],stage1_16[135],stage1_15[183]}
   );
   gpc615_5 gpc621 (
      {stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365], stage0_15[366]},
      {stage0_16[79]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[34],stage1_17[72],stage1_16[136],stage1_15[184]}
   );
   gpc615_5 gpc622 (
      {stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage0_16[80]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[35],stage1_17[73],stage1_16[137],stage1_15[185]}
   );
   gpc615_5 gpc623 (
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376]},
      {stage0_16[81]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[36],stage1_17[74],stage1_16[138],stage1_15[186]}
   );
   gpc615_5 gpc624 (
      {stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381]},
      {stage0_16[82]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[37],stage1_17[75],stage1_16[139],stage1_15[187]}
   );
   gpc615_5 gpc625 (
      {stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385], stage0_15[386]},
      {stage0_16[83]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[38],stage1_17[76],stage1_16[140],stage1_15[188]}
   );
   gpc615_5 gpc626 (
      {stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390], stage0_15[391]},
      {stage0_16[84]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[39],stage1_17[77],stage1_16[141],stage1_15[189]}
   );
   gpc615_5 gpc627 (
      {stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395], stage0_15[396]},
      {stage0_16[85]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[40],stage1_17[78],stage1_16[142],stage1_15[190]}
   );
   gpc615_5 gpc628 (
      {stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage0_16[86]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[41],stage1_17[79],stage1_16[143],stage1_15[191]}
   );
   gpc615_5 gpc629 (
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406]},
      {stage0_16[87]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[42],stage1_17[80],stage1_16[144],stage1_15[192]}
   );
   gpc615_5 gpc630 (
      {stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411]},
      {stage0_16[88]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[43],stage1_17[81],stage1_16[145],stage1_15[193]}
   );
   gpc615_5 gpc631 (
      {stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415], stage0_15[416]},
      {stage0_16[89]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[44],stage1_17[82],stage1_16[146],stage1_15[194]}
   );
   gpc615_5 gpc632 (
      {stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420], stage0_15[421]},
      {stage0_16[90]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[45],stage1_17[83],stage1_16[147],stage1_15[195]}
   );
   gpc615_5 gpc633 (
      {stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425], stage0_15[426]},
      {stage0_16[91]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[46],stage1_17[84],stage1_16[148],stage1_15[196]}
   );
   gpc615_5 gpc634 (
      {stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage0_16[92]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[47],stage1_17[85],stage1_16[149],stage1_15[197]}
   );
   gpc615_5 gpc635 (
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436]},
      {stage0_16[93]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[48],stage1_17[86],stage1_16[150],stage1_15[198]}
   );
   gpc615_5 gpc636 (
      {stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441]},
      {stage0_16[94]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[49],stage1_17[87],stage1_16[151],stage1_15[199]}
   );
   gpc615_5 gpc637 (
      {stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445], stage0_15[446]},
      {stage0_16[95]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[50],stage1_17[88],stage1_16[152],stage1_15[200]}
   );
   gpc615_5 gpc638 (
      {stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450], stage0_15[451]},
      {stage0_16[96]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[51],stage1_17[89],stage1_16[153],stage1_15[201]}
   );
   gpc615_5 gpc639 (
      {stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455], stage0_15[456]},
      {stage0_16[97]},
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage1_19[43],stage1_18[52],stage1_17[90],stage1_16[154],stage1_15[202]}
   );
   gpc606_5 gpc640 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[44],stage1_18[53],stage1_17[91],stage1_16[155]}
   );
   gpc606_5 gpc641 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[45],stage1_18[54],stage1_17[92],stage1_16[156]}
   );
   gpc606_5 gpc642 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[46],stage1_18[55],stage1_17[93],stage1_16[157]}
   );
   gpc606_5 gpc643 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[47],stage1_18[56],stage1_17[94],stage1_16[158]}
   );
   gpc606_5 gpc644 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[48],stage1_18[57],stage1_17[95],stage1_16[159]}
   );
   gpc606_5 gpc645 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[49],stage1_18[58],stage1_17[96],stage1_16[160]}
   );
   gpc606_5 gpc646 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[50],stage1_18[59],stage1_17[97],stage1_16[161]}
   );
   gpc606_5 gpc647 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[51],stage1_18[60],stage1_17[98],stage1_16[162]}
   );
   gpc606_5 gpc648 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[52],stage1_18[61],stage1_17[99],stage1_16[163]}
   );
   gpc606_5 gpc649 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[53],stage1_18[62],stage1_17[100],stage1_16[164]}
   );
   gpc606_5 gpc650 (
      {stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[54],stage1_18[63],stage1_17[101],stage1_16[165]}
   );
   gpc606_5 gpc651 (
      {stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[55],stage1_18[64],stage1_17[102],stage1_16[166]}
   );
   gpc606_5 gpc652 (
      {stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[56],stage1_18[65],stage1_17[103],stage1_16[167]}
   );
   gpc606_5 gpc653 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[57],stage1_18[66],stage1_17[104],stage1_16[168]}
   );
   gpc606_5 gpc654 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[58],stage1_18[67],stage1_17[105],stage1_16[169]}
   );
   gpc606_5 gpc655 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[59],stage1_18[68],stage1_17[106],stage1_16[170]}
   );
   gpc606_5 gpc656 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[60],stage1_18[69],stage1_17[107],stage1_16[171]}
   );
   gpc606_5 gpc657 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[61],stage1_18[70],stage1_17[108],stage1_16[172]}
   );
   gpc606_5 gpc658 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[62],stage1_18[71],stage1_17[109],stage1_16[173]}
   );
   gpc606_5 gpc659 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[63],stage1_18[72],stage1_17[110],stage1_16[174]}
   );
   gpc606_5 gpc660 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[64],stage1_18[73],stage1_17[111],stage1_16[175]}
   );
   gpc606_5 gpc661 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[65],stage1_18[74],stage1_17[112],stage1_16[176]}
   );
   gpc606_5 gpc662 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[66],stage1_18[75],stage1_17[113],stage1_16[177]}
   );
   gpc606_5 gpc663 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[67],stage1_18[76],stage1_17[114],stage1_16[178]}
   );
   gpc606_5 gpc664 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[68],stage1_18[77],stage1_17[115],stage1_16[179]}
   );
   gpc606_5 gpc665 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[69],stage1_18[78],stage1_17[116],stage1_16[180]}
   );
   gpc606_5 gpc666 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[70],stage1_18[79],stage1_17[117],stage1_16[181]}
   );
   gpc606_5 gpc667 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[71],stage1_18[80],stage1_17[118],stage1_16[182]}
   );
   gpc606_5 gpc668 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[72],stage1_18[81],stage1_17[119],stage1_16[183]}
   );
   gpc606_5 gpc669 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[73],stage1_18[82],stage1_17[120],stage1_16[184]}
   );
   gpc606_5 gpc670 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[74],stage1_18[83],stage1_17[121],stage1_16[185]}
   );
   gpc606_5 gpc671 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[75],stage1_18[84],stage1_17[122],stage1_16[186]}
   );
   gpc606_5 gpc672 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[76],stage1_18[85],stage1_17[123],stage1_16[187]}
   );
   gpc606_5 gpc673 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[77],stage1_18[86],stage1_17[124],stage1_16[188]}
   );
   gpc606_5 gpc674 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[78],stage1_18[87],stage1_17[125],stage1_16[189]}
   );
   gpc606_5 gpc675 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[79],stage1_18[88],stage1_17[126],stage1_16[190]}
   );
   gpc606_5 gpc676 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[80],stage1_18[89],stage1_17[127],stage1_16[191]}
   );
   gpc606_5 gpc677 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[81],stage1_18[90],stage1_17[128],stage1_16[192]}
   );
   gpc606_5 gpc678 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[82],stage1_18[91],stage1_17[129],stage1_16[193]}
   );
   gpc606_5 gpc679 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[83],stage1_18[92],stage1_17[130],stage1_16[194]}
   );
   gpc606_5 gpc680 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[84],stage1_18[93],stage1_17[131],stage1_16[195]}
   );
   gpc606_5 gpc681 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[85],stage1_18[94],stage1_17[132],stage1_16[196]}
   );
   gpc606_5 gpc682 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[86],stage1_18[95],stage1_17[133],stage1_16[197]}
   );
   gpc606_5 gpc683 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[87],stage1_18[96],stage1_17[134],stage1_16[198]}
   );
   gpc606_5 gpc684 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[88],stage1_18[97],stage1_17[135],stage1_16[199]}
   );
   gpc606_5 gpc685 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[89],stage1_18[98],stage1_17[136],stage1_16[200]}
   );
   gpc606_5 gpc686 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[90],stage1_18[99],stage1_17[137],stage1_16[201]}
   );
   gpc606_5 gpc687 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[91],stage1_18[100],stage1_17[138],stage1_16[202]}
   );
   gpc606_5 gpc688 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[92],stage1_18[101],stage1_17[139],stage1_16[203]}
   );
   gpc606_5 gpc689 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[93],stage1_18[102],stage1_17[140],stage1_16[204]}
   );
   gpc606_5 gpc690 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[94],stage1_18[103],stage1_17[141],stage1_16[205]}
   );
   gpc606_5 gpc691 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[95],stage1_18[104],stage1_17[142],stage1_16[206]}
   );
   gpc606_5 gpc692 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[96],stage1_18[105],stage1_17[143],stage1_16[207]}
   );
   gpc606_5 gpc693 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[97],stage1_18[106],stage1_17[144],stage1_16[208]}
   );
   gpc606_5 gpc694 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[98],stage1_18[107],stage1_17[145],stage1_16[209]}
   );
   gpc606_5 gpc695 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[99],stage1_18[108],stage1_17[146],stage1_16[210]}
   );
   gpc606_5 gpc696 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[100],stage1_18[109],stage1_17[147],stage1_16[211]}
   );
   gpc606_5 gpc697 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[101],stage1_18[110],stage1_17[148],stage1_16[212]}
   );
   gpc606_5 gpc698 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[102],stage1_18[111],stage1_17[149],stage1_16[213]}
   );
   gpc606_5 gpc699 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[103],stage1_18[112],stage1_17[150],stage1_16[214]}
   );
   gpc606_5 gpc700 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[104],stage1_18[113],stage1_17[151],stage1_16[215]}
   );
   gpc606_5 gpc701 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[105],stage1_18[114],stage1_17[152],stage1_16[216]}
   );
   gpc606_5 gpc702 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[106],stage1_18[115],stage1_17[153],stage1_16[217]}
   );
   gpc606_5 gpc703 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[107],stage1_18[116],stage1_17[154],stage1_16[218]}
   );
   gpc606_5 gpc704 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[108],stage1_18[117],stage1_17[155],stage1_16[219]}
   );
   gpc606_5 gpc705 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[109],stage1_18[118],stage1_17[156],stage1_16[220]}
   );
   gpc606_5 gpc706 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[110],stage1_18[119],stage1_17[157],stage1_16[221]}
   );
   gpc606_5 gpc707 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[111],stage1_18[120],stage1_17[158],stage1_16[222]}
   );
   gpc606_5 gpc708 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[112],stage1_18[121],stage1_17[159],stage1_16[223]}
   );
   gpc606_5 gpc709 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[69],stage1_19[113],stage1_18[122],stage1_17[160]}
   );
   gpc606_5 gpc710 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[70],stage1_19[114],stage1_18[123],stage1_17[161]}
   );
   gpc606_5 gpc711 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[71],stage1_19[115],stage1_18[124],stage1_17[162]}
   );
   gpc606_5 gpc712 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[72],stage1_19[116],stage1_18[125],stage1_17[163]}
   );
   gpc606_5 gpc713 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[73],stage1_19[117],stage1_18[126],stage1_17[164]}
   );
   gpc606_5 gpc714 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[74],stage1_19[118],stage1_18[127],stage1_17[165]}
   );
   gpc606_5 gpc715 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[75],stage1_19[119],stage1_18[128],stage1_17[166]}
   );
   gpc606_5 gpc716 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[76],stage1_19[120],stage1_18[129],stage1_17[167]}
   );
   gpc606_5 gpc717 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[77],stage1_19[121],stage1_18[130],stage1_17[168]}
   );
   gpc606_5 gpc718 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[78],stage1_19[122],stage1_18[131],stage1_17[169]}
   );
   gpc606_5 gpc719 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[79],stage1_19[123],stage1_18[132],stage1_17[170]}
   );
   gpc606_5 gpc720 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[80],stage1_19[124],stage1_18[133],stage1_17[171]}
   );
   gpc606_5 gpc721 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[81],stage1_19[125],stage1_18[134],stage1_17[172]}
   );
   gpc606_5 gpc722 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[82],stage1_19[126],stage1_18[135],stage1_17[173]}
   );
   gpc606_5 gpc723 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[83],stage1_19[127],stage1_18[136],stage1_17[174]}
   );
   gpc606_5 gpc724 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[84],stage1_19[128],stage1_18[137],stage1_17[175]}
   );
   gpc606_5 gpc725 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[85],stage1_19[129],stage1_18[138],stage1_17[176]}
   );
   gpc606_5 gpc726 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[86],stage1_19[130],stage1_18[139],stage1_17[177]}
   );
   gpc606_5 gpc727 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[87],stage1_19[131],stage1_18[140],stage1_17[178]}
   );
   gpc606_5 gpc728 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[88],stage1_19[132],stage1_18[141],stage1_17[179]}
   );
   gpc606_5 gpc729 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[89],stage1_19[133],stage1_18[142],stage1_17[180]}
   );
   gpc606_5 gpc730 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[90],stage1_19[134],stage1_18[143],stage1_17[181]}
   );
   gpc606_5 gpc731 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[91],stage1_19[135],stage1_18[144],stage1_17[182]}
   );
   gpc606_5 gpc732 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[92],stage1_19[136],stage1_18[145],stage1_17[183]}
   );
   gpc606_5 gpc733 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[93],stage1_19[137],stage1_18[146],stage1_17[184]}
   );
   gpc606_5 gpc734 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[94],stage1_19[138],stage1_18[147],stage1_17[185]}
   );
   gpc606_5 gpc735 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[95],stage1_19[139],stage1_18[148],stage1_17[186]}
   );
   gpc606_5 gpc736 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[96],stage1_19[140],stage1_18[149],stage1_17[187]}
   );
   gpc606_5 gpc737 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[97],stage1_19[141],stage1_18[150],stage1_17[188]}
   );
   gpc606_5 gpc738 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[98],stage1_19[142],stage1_18[151],stage1_17[189]}
   );
   gpc606_5 gpc739 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[99],stage1_19[143],stage1_18[152],stage1_17[190]}
   );
   gpc606_5 gpc740 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[100],stage1_19[144],stage1_18[153],stage1_17[191]}
   );
   gpc606_5 gpc741 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[101],stage1_19[145],stage1_18[154],stage1_17[192]}
   );
   gpc606_5 gpc742 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[102],stage1_19[146],stage1_18[155],stage1_17[193]}
   );
   gpc606_5 gpc743 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[103],stage1_19[147],stage1_18[156],stage1_17[194]}
   );
   gpc606_5 gpc744 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[104],stage1_19[148],stage1_18[157],stage1_17[195]}
   );
   gpc606_5 gpc745 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[105],stage1_19[149],stage1_18[158],stage1_17[196]}
   );
   gpc606_5 gpc746 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[106],stage1_19[150],stage1_18[159],stage1_17[197]}
   );
   gpc615_5 gpc747 (
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418]},
      {stage0_19[228]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[107],stage1_19[151],stage1_18[160]}
   );
   gpc615_5 gpc748 (
      {stage0_18[419], stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423]},
      {stage0_19[229]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[108],stage1_19[152],stage1_18[161]}
   );
   gpc615_5 gpc749 (
      {stage0_18[424], stage0_18[425], stage0_18[426], stage0_18[427], stage0_18[428]},
      {stage0_19[230]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[109],stage1_19[153],stage1_18[162]}
   );
   gpc615_5 gpc750 (
      {stage0_18[429], stage0_18[430], stage0_18[431], stage0_18[432], stage0_18[433]},
      {stage0_19[231]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[110],stage1_19[154],stage1_18[163]}
   );
   gpc615_5 gpc751 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[24]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[42],stage1_20[111],stage1_19[155]}
   );
   gpc615_5 gpc752 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[25]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[43],stage1_20[112],stage1_19[156]}
   );
   gpc615_5 gpc753 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[26]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[44],stage1_20[113],stage1_19[157]}
   );
   gpc615_5 gpc754 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[27]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[7],stage1_21[45],stage1_20[114],stage1_19[158]}
   );
   gpc615_5 gpc755 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[28]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[8],stage1_21[46],stage1_20[115],stage1_19[159]}
   );
   gpc615_5 gpc756 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[29]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[9],stage1_21[47],stage1_20[116],stage1_19[160]}
   );
   gpc615_5 gpc757 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[30]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[10],stage1_21[48],stage1_20[117],stage1_19[161]}
   );
   gpc615_5 gpc758 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[31]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[11],stage1_21[49],stage1_20[118],stage1_19[162]}
   );
   gpc615_5 gpc759 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[32]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[12],stage1_21[50],stage1_20[119],stage1_19[163]}
   );
   gpc615_5 gpc760 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[33]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[13],stage1_21[51],stage1_20[120],stage1_19[164]}
   );
   gpc615_5 gpc761 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[34]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[14],stage1_21[52],stage1_20[121],stage1_19[165]}
   );
   gpc615_5 gpc762 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[35]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[15],stage1_21[53],stage1_20[122],stage1_19[166]}
   );
   gpc615_5 gpc763 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[36]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[16],stage1_21[54],stage1_20[123],stage1_19[167]}
   );
   gpc615_5 gpc764 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[37]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[17],stage1_21[55],stage1_20[124],stage1_19[168]}
   );
   gpc615_5 gpc765 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[38]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[18],stage1_21[56],stage1_20[125],stage1_19[169]}
   );
   gpc615_5 gpc766 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[39]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[19],stage1_21[57],stage1_20[126],stage1_19[170]}
   );
   gpc615_5 gpc767 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[40]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[20],stage1_21[58],stage1_20[127],stage1_19[171]}
   );
   gpc615_5 gpc768 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[41]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[21],stage1_21[59],stage1_20[128],stage1_19[172]}
   );
   gpc615_5 gpc769 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[42]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[22],stage1_21[60],stage1_20[129],stage1_19[173]}
   );
   gpc615_5 gpc770 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[43]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[23],stage1_21[61],stage1_20[130],stage1_19[174]}
   );
   gpc615_5 gpc771 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[44]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[24],stage1_21[62],stage1_20[131],stage1_19[175]}
   );
   gpc615_5 gpc772 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[45]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[25],stage1_21[63],stage1_20[132],stage1_19[176]}
   );
   gpc615_5 gpc773 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[46]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[26],stage1_21[64],stage1_20[133],stage1_19[177]}
   );
   gpc615_5 gpc774 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[47]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[27],stage1_21[65],stage1_20[134],stage1_19[178]}
   );
   gpc615_5 gpc775 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[48]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[28],stage1_21[66],stage1_20[135],stage1_19[179]}
   );
   gpc615_5 gpc776 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[49]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[29],stage1_21[67],stage1_20[136],stage1_19[180]}
   );
   gpc615_5 gpc777 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[50]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[30],stage1_21[68],stage1_20[137],stage1_19[181]}
   );
   gpc615_5 gpc778 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[51]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[31],stage1_21[69],stage1_20[138],stage1_19[182]}
   );
   gpc615_5 gpc779 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[52]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[32],stage1_21[70],stage1_20[139],stage1_19[183]}
   );
   gpc615_5 gpc780 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[53]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[33],stage1_21[71],stage1_20[140],stage1_19[184]}
   );
   gpc615_5 gpc781 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[54]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[34],stage1_21[72],stage1_20[141],stage1_19[185]}
   );
   gpc615_5 gpc782 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[55]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[35],stage1_21[73],stage1_20[142],stage1_19[186]}
   );
   gpc615_5 gpc783 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[56]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[36],stage1_21[74],stage1_20[143],stage1_19[187]}
   );
   gpc615_5 gpc784 (
      {stage0_19[397], stage0_19[398], stage0_19[399], stage0_19[400], stage0_19[401]},
      {stage0_20[57]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[37],stage1_21[75],stage1_20[144],stage1_19[188]}
   );
   gpc615_5 gpc785 (
      {stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405], stage0_19[406]},
      {stage0_20[58]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[38],stage1_21[76],stage1_20[145],stage1_19[189]}
   );
   gpc615_5 gpc786 (
      {stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410], stage0_19[411]},
      {stage0_20[59]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[39],stage1_21[77],stage1_20[146],stage1_19[190]}
   );
   gpc615_5 gpc787 (
      {stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415], stage0_19[416]},
      {stage0_20[60]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[40],stage1_21[78],stage1_20[147],stage1_19[191]}
   );
   gpc615_5 gpc788 (
      {stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420], stage0_19[421]},
      {stage0_20[61]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[41],stage1_21[79],stage1_20[148],stage1_19[192]}
   );
   gpc615_5 gpc789 (
      {stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425], stage0_19[426]},
      {stage0_20[62]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[42],stage1_21[80],stage1_20[149],stage1_19[193]}
   );
   gpc615_5 gpc790 (
      {stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430], stage0_19[431]},
      {stage0_20[63]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[43],stage1_21[81],stage1_20[150],stage1_19[194]}
   );
   gpc615_5 gpc791 (
      {stage0_19[432], stage0_19[433], stage0_19[434], stage0_19[435], stage0_19[436]},
      {stage0_20[64]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[44],stage1_21[82],stage1_20[151],stage1_19[195]}
   );
   gpc615_5 gpc792 (
      {stage0_19[437], stage0_19[438], stage0_19[439], stage0_19[440], stage0_19[441]},
      {stage0_20[65]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage1_23[41],stage1_22[45],stage1_21[83],stage1_20[152],stage1_19[196]}
   );
   gpc615_5 gpc793 (
      {stage0_19[442], stage0_19[443], stage0_19[444], stage0_19[445], stage0_19[446]},
      {stage0_20[66]},
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage1_23[42],stage1_22[46],stage1_21[84],stage1_20[153],stage1_19[197]}
   );
   gpc615_5 gpc794 (
      {stage0_19[447], stage0_19[448], stage0_19[449], stage0_19[450], stage0_19[451]},
      {stage0_20[67]},
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage1_23[43],stage1_22[47],stage1_21[85],stage1_20[154],stage1_19[198]}
   );
   gpc615_5 gpc795 (
      {stage0_19[452], stage0_19[453], stage0_19[454], stage0_19[455], stage0_19[456]},
      {stage0_20[68]},
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage1_23[44],stage1_22[48],stage1_21[86],stage1_20[155],stage1_19[199]}
   );
   gpc615_5 gpc796 (
      {stage0_19[457], stage0_19[458], stage0_19[459], stage0_19[460], stage0_19[461]},
      {stage0_20[69]},
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage1_23[45],stage1_22[49],stage1_21[87],stage1_20[156],stage1_19[200]}
   );
   gpc615_5 gpc797 (
      {stage0_19[462], stage0_19[463], stage0_19[464], stage0_19[465], stage0_19[466]},
      {stage0_20[70]},
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage1_23[46],stage1_22[50],stage1_21[88],stage1_20[157],stage1_19[201]}
   );
   gpc615_5 gpc798 (
      {stage0_19[467], stage0_19[468], stage0_19[469], stage0_19[470], stage0_19[471]},
      {stage0_20[71]},
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage1_23[47],stage1_22[51],stage1_21[89],stage1_20[158],stage1_19[202]}
   );
   gpc615_5 gpc799 (
      {stage0_19[472], stage0_19[473], stage0_19[474], stage0_19[475], stage0_19[476]},
      {stage0_20[72]},
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage1_23[48],stage1_22[52],stage1_21[90],stage1_20[159],stage1_19[203]}
   );
   gpc615_5 gpc800 (
      {stage0_19[477], stage0_19[478], stage0_19[479], stage0_19[480], stage0_19[481]},
      {stage0_20[73]},
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage1_23[49],stage1_22[53],stage1_21[91],stage1_20[160],stage1_19[204]}
   );
   gpc615_5 gpc801 (
      {stage0_19[482], stage0_19[483], stage0_19[484], stage0_19[485], stage0_19[486]},
      {stage0_20[74]},
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage1_23[50],stage1_22[54],stage1_21[92],stage1_20[161],stage1_19[205]}
   );
   gpc615_5 gpc802 (
      {stage0_19[487], stage0_19[488], stage0_19[489], stage0_19[490], stage0_19[491]},
      {stage0_20[75]},
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage1_23[51],stage1_22[55],stage1_21[93],stage1_20[162],stage1_19[206]}
   );
   gpc615_5 gpc803 (
      {stage0_19[492], stage0_19[493], stage0_19[494], stage0_19[495], stage0_19[496]},
      {stage0_20[76]},
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage1_23[52],stage1_22[56],stage1_21[94],stage1_20[163],stage1_19[207]}
   );
   gpc615_5 gpc804 (
      {stage0_19[497], stage0_19[498], stage0_19[499], stage0_19[500], stage0_19[501]},
      {stage0_20[77]},
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage1_23[53],stage1_22[57],stage1_21[95],stage1_20[164],stage1_19[208]}
   );
   gpc606_5 gpc805 (
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[54],stage1_22[58],stage1_21[96],stage1_20[165]}
   );
   gpc606_5 gpc806 (
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[55],stage1_22[59],stage1_21[97],stage1_20[166]}
   );
   gpc606_5 gpc807 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[56],stage1_22[60],stage1_21[98],stage1_20[167]}
   );
   gpc606_5 gpc808 (
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[57],stage1_22[61],stage1_21[99],stage1_20[168]}
   );
   gpc606_5 gpc809 (
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[58],stage1_22[62],stage1_21[100],stage1_20[169]}
   );
   gpc606_5 gpc810 (
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[59],stage1_22[63],stage1_21[101],stage1_20[170]}
   );
   gpc606_5 gpc811 (
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[60],stage1_22[64],stage1_21[102],stage1_20[171]}
   );
   gpc606_5 gpc812 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[61],stage1_22[65],stage1_21[103],stage1_20[172]}
   );
   gpc606_5 gpc813 (
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[62],stage1_22[66],stage1_21[104],stage1_20[173]}
   );
   gpc606_5 gpc814 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[63],stage1_22[67],stage1_21[105],stage1_20[174]}
   );
   gpc606_5 gpc815 (
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[64],stage1_22[68],stage1_21[106],stage1_20[175]}
   );
   gpc606_5 gpc816 (
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[65],stage1_22[69],stage1_21[107],stage1_20[176]}
   );
   gpc606_5 gpc817 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[66],stage1_22[70],stage1_21[108],stage1_20[177]}
   );
   gpc606_5 gpc818 (
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[67],stage1_22[71],stage1_21[109],stage1_20[178]}
   );
   gpc606_5 gpc819 (
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[68],stage1_22[72],stage1_21[110],stage1_20[179]}
   );
   gpc606_5 gpc820 (
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[69],stage1_22[73],stage1_21[111],stage1_20[180]}
   );
   gpc606_5 gpc821 (
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[70],stage1_22[74],stage1_21[112],stage1_20[181]}
   );
   gpc606_5 gpc822 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[71],stage1_22[75],stage1_21[113],stage1_20[182]}
   );
   gpc606_5 gpc823 (
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[72],stage1_22[76],stage1_21[114],stage1_20[183]}
   );
   gpc606_5 gpc824 (
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[73],stage1_22[77],stage1_21[115],stage1_20[184]}
   );
   gpc606_5 gpc825 (
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[74],stage1_22[78],stage1_21[116],stage1_20[185]}
   );
   gpc606_5 gpc826 (
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[75],stage1_22[79],stage1_21[117],stage1_20[186]}
   );
   gpc606_5 gpc827 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[76],stage1_22[80],stage1_21[118],stage1_20[187]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[77],stage1_22[81],stage1_21[119],stage1_20[188]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[78],stage1_22[82],stage1_21[120],stage1_20[189]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[79],stage1_22[83],stage1_21[121],stage1_20[190]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[80],stage1_22[84],stage1_21[122],stage1_20[191]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[81],stage1_22[85],stage1_21[123],stage1_20[192]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[82],stage1_22[86],stage1_21[124],stage1_20[193]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[83],stage1_22[87],stage1_21[125],stage1_20[194]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[84],stage1_22[88],stage1_21[126],stage1_20[195]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[85],stage1_22[89],stage1_21[127],stage1_20[196]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[86],stage1_22[90],stage1_21[128],stage1_20[197]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[87],stage1_22[91],stage1_21[129],stage1_20[198]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[88],stage1_22[92],stage1_21[130],stage1_20[199]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[89],stage1_22[93],stage1_21[131],stage1_20[200]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[90],stage1_22[94],stage1_21[132],stage1_20[201]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[91],stage1_22[95],stage1_21[133],stage1_20[202]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[92],stage1_22[96],stage1_21[134],stage1_20[203]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[93],stage1_22[97],stage1_21[135],stage1_20[204]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[94],stage1_22[98],stage1_21[136],stage1_20[205]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[95],stage1_22[99],stage1_21[137],stage1_20[206]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[96],stage1_22[100],stage1_21[138],stage1_20[207]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[97],stage1_22[101],stage1_21[139],stage1_20[208]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[98],stage1_22[102],stage1_21[140],stage1_20[209]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[99],stage1_22[103],stage1_21[141],stage1_20[210]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[100],stage1_22[104],stage1_21[142],stage1_20[211]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[101],stage1_22[105],stage1_21[143],stage1_20[212]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291], stage0_22[292], stage0_22[293]},
      {stage1_24[48],stage1_23[102],stage1_22[106],stage1_21[144],stage1_20[213]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[294], stage0_22[295], stage0_22[296], stage0_22[297], stage0_22[298], stage0_22[299]},
      {stage1_24[49],stage1_23[103],stage1_22[107],stage1_21[145],stage1_20[214]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[300], stage0_22[301], stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305]},
      {stage1_24[50],stage1_23[104],stage1_22[108],stage1_21[146],stage1_20[215]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[306], stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage1_24[51],stage1_23[105],stage1_22[109],stage1_21[147],stage1_20[216]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316], stage0_22[317]},
      {stage1_24[52],stage1_23[106],stage1_22[110],stage1_21[148],stage1_20[217]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321], stage0_22[322], stage0_22[323]},
      {stage1_24[53],stage1_23[107],stage1_22[111],stage1_21[149],stage1_20[218]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[324], stage0_22[325], stage0_22[326], stage0_22[327], stage0_22[328], stage0_22[329]},
      {stage1_24[54],stage1_23[108],stage1_22[112],stage1_21[150],stage1_20[219]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[330], stage0_22[331], stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335]},
      {stage1_24[55],stage1_23[109],stage1_22[113],stage1_21[151],stage1_20[220]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[336], stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage1_24[56],stage1_23[110],stage1_22[114],stage1_21[152],stage1_20[221]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346], stage0_22[347]},
      {stage1_24[57],stage1_23[111],stage1_22[115],stage1_21[153],stage1_20[222]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351], stage0_22[352], stage0_22[353]},
      {stage1_24[58],stage1_23[112],stage1_22[116],stage1_21[154],stage1_20[223]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[354], stage0_22[355], stage0_22[356], stage0_22[357], stage0_22[358], stage0_22[359]},
      {stage1_24[59],stage1_23[113],stage1_22[117],stage1_21[155],stage1_20[224]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[360], stage0_22[361], stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365]},
      {stage1_24[60],stage1_23[114],stage1_22[118],stage1_21[156],stage1_20[225]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[366], stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage1_24[61],stage1_23[115],stage1_22[119],stage1_21[157],stage1_20[226]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376], stage0_22[377]},
      {stage1_24[62],stage1_23[116],stage1_22[120],stage1_21[158],stage1_20[227]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381], stage0_22[382], stage0_22[383]},
      {stage1_24[63],stage1_23[117],stage1_22[121],stage1_21[159],stage1_20[228]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[384], stage0_22[385], stage0_22[386], stage0_22[387], stage0_22[388], stage0_22[389]},
      {stage1_24[64],stage1_23[118],stage1_22[122],stage1_21[160],stage1_20[229]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[390], stage0_22[391], stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395]},
      {stage1_24[65],stage1_23[119],stage1_22[123],stage1_21[161],stage1_20[230]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[396], stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage1_24[66],stage1_23[120],stage1_22[124],stage1_21[162],stage1_20[231]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage1_24[67],stage1_23[121],stage1_22[125],stage1_21[163],stage1_20[232]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412], stage0_22[413]},
      {stage1_24[68],stage1_23[122],stage1_22[126],stage1_21[164],stage1_20[233]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417], stage0_22[418], stage0_22[419]},
      {stage1_24[69],stage1_23[123],stage1_22[127],stage1_21[165],stage1_20[234]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[420], stage0_22[421], stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425]},
      {stage1_24[70],stage1_23[124],stage1_22[128],stage1_21[166],stage1_20[235]}
   );
   gpc606_5 gpc876 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[71],stage1_23[125],stage1_22[129],stage1_21[167]}
   );
   gpc606_5 gpc877 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[72],stage1_23[126],stage1_22[130],stage1_21[168]}
   );
   gpc606_5 gpc878 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[73],stage1_23[127],stage1_22[131],stage1_21[169]}
   );
   gpc606_5 gpc879 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[74],stage1_23[128],stage1_22[132],stage1_21[170]}
   );
   gpc606_5 gpc880 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[75],stage1_23[129],stage1_22[133],stage1_21[171]}
   );
   gpc606_5 gpc881 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[76],stage1_23[130],stage1_22[134],stage1_21[172]}
   );
   gpc606_5 gpc882 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[77],stage1_23[131],stage1_22[135],stage1_21[173]}
   );
   gpc606_5 gpc883 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[78],stage1_23[132],stage1_22[136],stage1_21[174]}
   );
   gpc606_5 gpc884 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[79],stage1_23[133],stage1_22[137],stage1_21[175]}
   );
   gpc606_5 gpc885 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[80],stage1_23[134],stage1_22[138],stage1_21[176]}
   );
   gpc606_5 gpc886 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[81],stage1_23[135],stage1_22[139],stage1_21[177]}
   );
   gpc606_5 gpc887 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[82],stage1_23[136],stage1_22[140],stage1_21[178]}
   );
   gpc606_5 gpc888 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[83],stage1_23[137],stage1_22[141],stage1_21[179]}
   );
   gpc606_5 gpc889 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[84],stage1_23[138],stage1_22[142],stage1_21[180]}
   );
   gpc606_5 gpc890 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[85],stage1_23[139],stage1_22[143],stage1_21[181]}
   );
   gpc606_5 gpc891 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[86],stage1_23[140],stage1_22[144],stage1_21[182]}
   );
   gpc606_5 gpc892 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[87],stage1_23[141],stage1_22[145],stage1_21[183]}
   );
   gpc606_5 gpc893 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[88],stage1_23[142],stage1_22[146],stage1_21[184]}
   );
   gpc606_5 gpc894 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[89],stage1_23[143],stage1_22[147],stage1_21[185]}
   );
   gpc606_5 gpc895 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[90],stage1_23[144],stage1_22[148],stage1_21[186]}
   );
   gpc606_5 gpc896 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[91],stage1_23[145],stage1_22[149],stage1_21[187]}
   );
   gpc606_5 gpc897 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[92],stage1_23[146],stage1_22[150],stage1_21[188]}
   );
   gpc606_5 gpc898 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[93],stage1_23[147],stage1_22[151],stage1_21[189]}
   );
   gpc606_5 gpc899 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[94],stage1_23[148],stage1_22[152],stage1_21[190]}
   );
   gpc606_5 gpc900 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[95],stage1_23[149],stage1_22[153],stage1_21[191]}
   );
   gpc606_5 gpc901 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[96],stage1_23[150],stage1_22[154],stage1_21[192]}
   );
   gpc606_5 gpc902 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[97],stage1_23[151],stage1_22[155],stage1_21[193]}
   );
   gpc606_5 gpc903 (
      {stage0_21[486], stage0_21[487], stage0_21[488], stage0_21[489], stage0_21[490], stage0_21[491]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[98],stage1_23[152],stage1_22[156],stage1_21[194]}
   );
   gpc606_5 gpc904 (
      {stage0_21[492], stage0_21[493], stage0_21[494], stage0_21[495], stage0_21[496], stage0_21[497]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[99],stage1_23[153],stage1_22[157],stage1_21[195]}
   );
   gpc606_5 gpc905 (
      {stage0_21[498], stage0_21[499], stage0_21[500], stage0_21[501], stage0_21[502], stage0_21[503]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[100],stage1_23[154],stage1_22[158],stage1_21[196]}
   );
   gpc615_5 gpc906 (
      {stage0_22[426], stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430]},
      {stage0_23[180]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[30],stage1_24[101],stage1_23[155],stage1_22[159]}
   );
   gpc615_5 gpc907 (
      {stage0_22[431], stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435]},
      {stage0_23[181]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[31],stage1_24[102],stage1_23[156],stage1_22[160]}
   );
   gpc615_5 gpc908 (
      {stage0_22[436], stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440]},
      {stage0_23[182]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[32],stage1_24[103],stage1_23[157],stage1_22[161]}
   );
   gpc615_5 gpc909 (
      {stage0_22[441], stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445]},
      {stage0_23[183]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[33],stage1_24[104],stage1_23[158],stage1_22[162]}
   );
   gpc615_5 gpc910 (
      {stage0_22[446], stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450]},
      {stage0_23[184]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[34],stage1_24[105],stage1_23[159],stage1_22[163]}
   );
   gpc615_5 gpc911 (
      {stage0_22[451], stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455]},
      {stage0_23[185]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[35],stage1_24[106],stage1_23[160],stage1_22[164]}
   );
   gpc615_5 gpc912 (
      {stage0_22[456], stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460]},
      {stage0_23[186]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[36],stage1_24[107],stage1_23[161],stage1_22[165]}
   );
   gpc615_5 gpc913 (
      {stage0_22[461], stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465]},
      {stage0_23[187]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[37],stage1_24[108],stage1_23[162],stage1_22[166]}
   );
   gpc615_5 gpc914 (
      {stage0_22[466], stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470]},
      {stage0_23[188]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[38],stage1_24[109],stage1_23[163],stage1_22[167]}
   );
   gpc615_5 gpc915 (
      {stage0_22[471], stage0_22[472], stage0_22[473], stage0_22[474], stage0_22[475]},
      {stage0_23[189]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[39],stage1_24[110],stage1_23[164],stage1_22[168]}
   );
   gpc615_5 gpc916 (
      {stage0_22[476], stage0_22[477], stage0_22[478], stage0_22[479], stage0_22[480]},
      {stage0_23[190]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[40],stage1_24[111],stage1_23[165],stage1_22[169]}
   );
   gpc606_5 gpc917 (
      {stage0_23[191], stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[11],stage1_25[41],stage1_24[112],stage1_23[166]}
   );
   gpc606_5 gpc918 (
      {stage0_23[197], stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[12],stage1_25[42],stage1_24[113],stage1_23[167]}
   );
   gpc606_5 gpc919 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[13],stage1_25[43],stage1_24[114],stage1_23[168]}
   );
   gpc606_5 gpc920 (
      {stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[14],stage1_25[44],stage1_24[115],stage1_23[169]}
   );
   gpc606_5 gpc921 (
      {stage0_23[215], stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[15],stage1_25[45],stage1_24[116],stage1_23[170]}
   );
   gpc606_5 gpc922 (
      {stage0_23[221], stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[16],stage1_25[46],stage1_24[117],stage1_23[171]}
   );
   gpc606_5 gpc923 (
      {stage0_23[227], stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[17],stage1_25[47],stage1_24[118],stage1_23[172]}
   );
   gpc606_5 gpc924 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[18],stage1_25[48],stage1_24[119],stage1_23[173]}
   );
   gpc606_5 gpc925 (
      {stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[19],stage1_25[49],stage1_24[120],stage1_23[174]}
   );
   gpc606_5 gpc926 (
      {stage0_23[245], stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[20],stage1_25[50],stage1_24[121],stage1_23[175]}
   );
   gpc606_5 gpc927 (
      {stage0_23[251], stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[21],stage1_25[51],stage1_24[122],stage1_23[176]}
   );
   gpc606_5 gpc928 (
      {stage0_23[257], stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[22],stage1_25[52],stage1_24[123],stage1_23[177]}
   );
   gpc606_5 gpc929 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[23],stage1_25[53],stage1_24[124],stage1_23[178]}
   );
   gpc606_5 gpc930 (
      {stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[24],stage1_25[54],stage1_24[125],stage1_23[179]}
   );
   gpc606_5 gpc931 (
      {stage0_23[275], stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[25],stage1_25[55],stage1_24[126],stage1_23[180]}
   );
   gpc606_5 gpc932 (
      {stage0_23[281], stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[26],stage1_25[56],stage1_24[127],stage1_23[181]}
   );
   gpc606_5 gpc933 (
      {stage0_23[287], stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[27],stage1_25[57],stage1_24[128],stage1_23[182]}
   );
   gpc606_5 gpc934 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[28],stage1_25[58],stage1_24[129],stage1_23[183]}
   );
   gpc606_5 gpc935 (
      {stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[29],stage1_25[59],stage1_24[130],stage1_23[184]}
   );
   gpc606_5 gpc936 (
      {stage0_23[305], stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[30],stage1_25[60],stage1_24[131],stage1_23[185]}
   );
   gpc606_5 gpc937 (
      {stage0_23[311], stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[31],stage1_25[61],stage1_24[132],stage1_23[186]}
   );
   gpc606_5 gpc938 (
      {stage0_23[317], stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[32],stage1_25[62],stage1_24[133],stage1_23[187]}
   );
   gpc606_5 gpc939 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[33],stage1_25[63],stage1_24[134],stage1_23[188]}
   );
   gpc606_5 gpc940 (
      {stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[34],stage1_25[64],stage1_24[135],stage1_23[189]}
   );
   gpc606_5 gpc941 (
      {stage0_23[335], stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[35],stage1_25[65],stage1_24[136],stage1_23[190]}
   );
   gpc606_5 gpc942 (
      {stage0_23[341], stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[36],stage1_25[66],stage1_24[137],stage1_23[191]}
   );
   gpc606_5 gpc943 (
      {stage0_23[347], stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[37],stage1_25[67],stage1_24[138],stage1_23[192]}
   );
   gpc606_5 gpc944 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[38],stage1_25[68],stage1_24[139],stage1_23[193]}
   );
   gpc606_5 gpc945 (
      {stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[39],stage1_25[69],stage1_24[140],stage1_23[194]}
   );
   gpc606_5 gpc946 (
      {stage0_23[365], stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[40],stage1_25[70],stage1_24[141],stage1_23[195]}
   );
   gpc606_5 gpc947 (
      {stage0_23[371], stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[41],stage1_25[71],stage1_24[142],stage1_23[196]}
   );
   gpc606_5 gpc948 (
      {stage0_23[377], stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[42],stage1_25[72],stage1_24[143],stage1_23[197]}
   );
   gpc615_5 gpc949 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[66]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[43],stage1_25[73],stage1_24[144],stage1_23[198]}
   );
   gpc615_5 gpc950 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[67]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[44],stage1_25[74],stage1_24[145],stage1_23[199]}
   );
   gpc615_5 gpc951 (
      {stage0_23[393], stage0_23[394], stage0_23[395], stage0_23[396], stage0_23[397]},
      {stage0_24[68]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[45],stage1_25[75],stage1_24[146],stage1_23[200]}
   );
   gpc615_5 gpc952 (
      {stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401], stage0_23[402]},
      {stage0_24[69]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[46],stage1_25[76],stage1_24[147],stage1_23[201]}
   );
   gpc615_5 gpc953 (
      {stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage0_24[70]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[47],stage1_25[77],stage1_24[148],stage1_23[202]}
   );
   gpc615_5 gpc954 (
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412]},
      {stage0_24[71]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[48],stage1_25[78],stage1_24[149],stage1_23[203]}
   );
   gpc615_5 gpc955 (
      {stage0_23[413], stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417]},
      {stage0_24[72]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[49],stage1_25[79],stage1_24[150],stage1_23[204]}
   );
   gpc606_5 gpc956 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[39],stage1_26[50],stage1_25[80],stage1_24[151]}
   );
   gpc606_5 gpc957 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[40],stage1_26[51],stage1_25[81],stage1_24[152]}
   );
   gpc606_5 gpc958 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[41],stage1_26[52],stage1_25[82],stage1_24[153]}
   );
   gpc606_5 gpc959 (
      {stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[42],stage1_26[53],stage1_25[83],stage1_24[154]}
   );
   gpc606_5 gpc960 (
      {stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[43],stage1_26[54],stage1_25[84],stage1_24[155]}
   );
   gpc606_5 gpc961 (
      {stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[44],stage1_26[55],stage1_25[85],stage1_24[156]}
   );
   gpc606_5 gpc962 (
      {stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113], stage0_24[114]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[45],stage1_26[56],stage1_25[86],stage1_24[157]}
   );
   gpc606_5 gpc963 (
      {stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119], stage0_24[120]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[46],stage1_26[57],stage1_25[87],stage1_24[158]}
   );
   gpc606_5 gpc964 (
      {stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125], stage0_24[126]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[47],stage1_26[58],stage1_25[88],stage1_24[159]}
   );
   gpc606_5 gpc965 (
      {stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131], stage0_24[132]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[48],stage1_26[59],stage1_25[89],stage1_24[160]}
   );
   gpc606_5 gpc966 (
      {stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137], stage0_24[138]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[49],stage1_26[60],stage1_25[90],stage1_24[161]}
   );
   gpc606_5 gpc967 (
      {stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143], stage0_24[144]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[50],stage1_26[61],stage1_25[91],stage1_24[162]}
   );
   gpc606_5 gpc968 (
      {stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149], stage0_24[150]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[51],stage1_26[62],stage1_25[92],stage1_24[163]}
   );
   gpc606_5 gpc969 (
      {stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155], stage0_24[156]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[52],stage1_26[63],stage1_25[93],stage1_24[164]}
   );
   gpc606_5 gpc970 (
      {stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161], stage0_24[162]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[53],stage1_26[64],stage1_25[94],stage1_24[165]}
   );
   gpc606_5 gpc971 (
      {stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167], stage0_24[168]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[54],stage1_26[65],stage1_25[95],stage1_24[166]}
   );
   gpc606_5 gpc972 (
      {stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172], stage0_24[173], stage0_24[174]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[55],stage1_26[66],stage1_25[96],stage1_24[167]}
   );
   gpc606_5 gpc973 (
      {stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178], stage0_24[179], stage0_24[180]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[56],stage1_26[67],stage1_25[97],stage1_24[168]}
   );
   gpc606_5 gpc974 (
      {stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184], stage0_24[185], stage0_24[186]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[57],stage1_26[68],stage1_25[98],stage1_24[169]}
   );
   gpc606_5 gpc975 (
      {stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190], stage0_24[191], stage0_24[192]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[58],stage1_26[69],stage1_25[99],stage1_24[170]}
   );
   gpc606_5 gpc976 (
      {stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196], stage0_24[197], stage0_24[198]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[59],stage1_26[70],stage1_25[100],stage1_24[171]}
   );
   gpc606_5 gpc977 (
      {stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[60],stage1_26[71],stage1_25[101],stage1_24[172]}
   );
   gpc606_5 gpc978 (
      {stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[61],stage1_26[72],stage1_25[102],stage1_24[173]}
   );
   gpc606_5 gpc979 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215], stage0_24[216]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[62],stage1_26[73],stage1_25[103],stage1_24[174]}
   );
   gpc606_5 gpc980 (
      {stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220], stage0_24[221], stage0_24[222]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[63],stage1_26[74],stage1_25[104],stage1_24[175]}
   );
   gpc606_5 gpc981 (
      {stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226], stage0_24[227], stage0_24[228]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[64],stage1_26[75],stage1_25[105],stage1_24[176]}
   );
   gpc606_5 gpc982 (
      {stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[65],stage1_26[76],stage1_25[106],stage1_24[177]}
   );
   gpc606_5 gpc983 (
      {stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[66],stage1_26[77],stage1_25[107],stage1_24[178]}
   );
   gpc606_5 gpc984 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245], stage0_24[246]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[67],stage1_26[78],stage1_25[108],stage1_24[179]}
   );
   gpc606_5 gpc985 (
      {stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250], stage0_24[251], stage0_24[252]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[68],stage1_26[79],stage1_25[109],stage1_24[180]}
   );
   gpc606_5 gpc986 (
      {stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256], stage0_24[257], stage0_24[258]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[69],stage1_26[80],stage1_25[110],stage1_24[181]}
   );
   gpc606_5 gpc987 (
      {stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[70],stage1_26[81],stage1_25[111],stage1_24[182]}
   );
   gpc606_5 gpc988 (
      {stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[71],stage1_26[82],stage1_25[112],stage1_24[183]}
   );
   gpc606_5 gpc989 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275], stage0_24[276]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[72],stage1_26[83],stage1_25[113],stage1_24[184]}
   );
   gpc606_5 gpc990 (
      {stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280], stage0_24[281], stage0_24[282]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[73],stage1_26[84],stage1_25[114],stage1_24[185]}
   );
   gpc606_5 gpc991 (
      {stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286], stage0_24[287], stage0_24[288]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[74],stage1_26[85],stage1_25[115],stage1_24[186]}
   );
   gpc606_5 gpc992 (
      {stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[75],stage1_26[86],stage1_25[116],stage1_24[187]}
   );
   gpc606_5 gpc993 (
      {stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[76],stage1_26[87],stage1_25[117],stage1_24[188]}
   );
   gpc606_5 gpc994 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305], stage0_24[306]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[77],stage1_26[88],stage1_25[118],stage1_24[189]}
   );
   gpc606_5 gpc995 (
      {stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310], stage0_24[311], stage0_24[312]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[78],stage1_26[89],stage1_25[119],stage1_24[190]}
   );
   gpc606_5 gpc996 (
      {stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316], stage0_24[317], stage0_24[318]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[79],stage1_26[90],stage1_25[120],stage1_24[191]}
   );
   gpc606_5 gpc997 (
      {stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[80],stage1_26[91],stage1_25[121],stage1_24[192]}
   );
   gpc606_5 gpc998 (
      {stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[81],stage1_26[92],stage1_25[122],stage1_24[193]}
   );
   gpc606_5 gpc999 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335], stage0_24[336]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[82],stage1_26[93],stage1_25[123],stage1_24[194]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340], stage0_24[341], stage0_24[342]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[83],stage1_26[94],stage1_25[124],stage1_24[195]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346], stage0_24[347], stage0_24[348]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[84],stage1_26[95],stage1_25[125],stage1_24[196]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[85],stage1_26[96],stage1_25[126],stage1_24[197]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[86],stage1_26[97],stage1_25[127],stage1_24[198]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[87],stage1_26[98],stage1_25[128],stage1_24[199]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371], stage0_24[372]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[88],stage1_26[99],stage1_25[129],stage1_24[200]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376], stage0_24[377], stage0_24[378]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[89],stage1_26[100],stage1_25[130],stage1_24[201]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[90],stage1_26[101],stage1_25[131],stage1_24[202]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[91],stage1_26[102],stage1_25[132],stage1_24[203]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[92],stage1_26[103],stage1_25[133],stage1_24[204]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401], stage0_24[402]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[93],stage1_26[104],stage1_25[134],stage1_24[205]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406], stage0_24[407], stage0_24[408]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[94],stage1_26[105],stage1_25[135],stage1_24[206]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[95],stage1_26[106],stage1_25[136],stage1_24[207]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[96],stage1_26[107],stage1_25[137],stage1_24[208]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[97],stage1_26[108],stage1_25[138],stage1_24[209]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431], stage0_24[432]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[98],stage1_26[109],stage1_25[139],stage1_24[210]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436], stage0_24[437], stage0_24[438]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[99],stage1_26[110],stage1_25[140],stage1_24[211]}
   );
   gpc606_5 gpc1017 (
      {stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[100],stage1_26[111],stage1_25[141],stage1_24[212]}
   );
   gpc606_5 gpc1018 (
      {stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[101],stage1_26[112],stage1_25[142],stage1_24[213]}
   );
   gpc606_5 gpc1019 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[102],stage1_26[113],stage1_25[143],stage1_24[214]}
   );
   gpc606_5 gpc1020 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461], stage0_24[462]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[103],stage1_26[114],stage1_25[144],stage1_24[215]}
   );
   gpc606_5 gpc1021 (
      {stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466], stage0_24[467], stage0_24[468]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[104],stage1_26[115],stage1_25[145],stage1_24[216]}
   );
   gpc606_5 gpc1022 (
      {stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[105],stage1_26[116],stage1_25[146],stage1_24[217]}
   );
   gpc606_5 gpc1023 (
      {stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[106],stage1_26[117],stage1_25[147],stage1_24[218]}
   );
   gpc606_5 gpc1024 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[107],stage1_26[118],stage1_25[148],stage1_24[219]}
   );
   gpc606_5 gpc1025 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491], stage0_24[492]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[108],stage1_26[119],stage1_25[149],stage1_24[220]}
   );
   gpc606_5 gpc1026 (
      {stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496], stage0_24[497], stage0_24[498]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[109],stage1_26[120],stage1_25[150],stage1_24[221]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[71],stage1_27[110],stage1_26[121],stage1_25[151]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[72],stage1_27[111],stage1_26[122],stage1_25[152]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[426]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[73],stage1_27[112],stage1_26[123],stage1_25[153]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[427]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[74],stage1_27[113],stage1_26[124],stage1_25[154]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[428]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[75],stage1_27[114],stage1_26[125],stage1_25[155]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[429]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[76],stage1_27[115],stage1_26[126],stage1_25[156]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[430]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[77],stage1_27[116],stage1_26[127],stage1_25[157]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[431]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[78],stage1_27[117],stage1_26[128],stage1_25[158]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[432]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[79],stage1_27[118],stage1_26[129],stage1_25[159]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[433]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[80],stage1_27[119],stage1_26[130],stage1_25[160]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[434]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[81],stage1_27[120],stage1_26[131],stage1_25[161]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[435]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[82],stage1_27[121],stage1_26[132],stage1_25[162]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[436]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[83],stage1_27[122],stage1_26[133],stage1_25[163]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[437]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[84],stage1_27[123],stage1_26[134],stage1_25[164]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[438]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[85],stage1_27[124],stage1_26[135],stage1_25[165]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[439]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[86],stage1_27[125],stage1_26[136],stage1_25[166]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[440]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[87],stage1_27[126],stage1_26[137],stage1_25[167]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[441]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[88],stage1_27[127],stage1_26[138],stage1_25[168]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[442]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[89],stage1_27[128],stage1_26[139],stage1_25[169]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[443]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[90],stage1_27[129],stage1_26[140],stage1_25[170]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[444]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[91],stage1_27[130],stage1_26[141],stage1_25[171]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[445]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[92],stage1_27[131],stage1_26[142],stage1_25[172]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[446]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[93],stage1_27[132],stage1_26[143],stage1_25[173]}
   );
   gpc615_5 gpc1050 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[447]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[94],stage1_27[133],stage1_26[144],stage1_25[174]}
   );
   gpc615_5 gpc1051 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[448]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[95],stage1_27[134],stage1_26[145],stage1_25[175]}
   );
   gpc615_5 gpc1052 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[449]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[96],stage1_27[135],stage1_26[146],stage1_25[176]}
   );
   gpc615_5 gpc1053 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[450]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[97],stage1_27[136],stage1_26[147],stage1_25[177]}
   );
   gpc615_5 gpc1054 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[451]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[98],stage1_27[137],stage1_26[148],stage1_25[178]}
   );
   gpc615_5 gpc1055 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[452]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[99],stage1_27[138],stage1_26[149],stage1_25[179]}
   );
   gpc615_5 gpc1056 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[453]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[100],stage1_27[139],stage1_26[150],stage1_25[180]}
   );
   gpc615_5 gpc1057 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[454]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[101],stage1_27[140],stage1_26[151],stage1_25[181]}
   );
   gpc615_5 gpc1058 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[455]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[102],stage1_27[141],stage1_26[152],stage1_25[182]}
   );
   gpc615_5 gpc1059 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[456]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[103],stage1_27[142],stage1_26[153],stage1_25[183]}
   );
   gpc615_5 gpc1060 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[457]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[104],stage1_27[143],stage1_26[154],stage1_25[184]}
   );
   gpc615_5 gpc1061 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[458]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[105],stage1_27[144],stage1_26[155],stage1_25[185]}
   );
   gpc615_5 gpc1062 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[459]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[106],stage1_27[145],stage1_26[156],stage1_25[186]}
   );
   gpc615_5 gpc1063 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[460]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[107],stage1_27[146],stage1_26[157],stage1_25[187]}
   );
   gpc615_5 gpc1064 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[461]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[108],stage1_27[147],stage1_26[158],stage1_25[188]}
   );
   gpc615_5 gpc1065 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[462]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[109],stage1_27[148],stage1_26[159],stage1_25[189]}
   );
   gpc615_5 gpc1066 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[463]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[110],stage1_27[149],stage1_26[160],stage1_25[190]}
   );
   gpc615_5 gpc1067 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[464]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[111],stage1_27[150],stage1_26[161],stage1_25[191]}
   );
   gpc615_5 gpc1068 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[465]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[112],stage1_27[151],stage1_26[162],stage1_25[192]}
   );
   gpc615_5 gpc1069 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[466]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[113],stage1_27[152],stage1_26[163],stage1_25[193]}
   );
   gpc615_5 gpc1070 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[467]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[114],stage1_27[153],stage1_26[164],stage1_25[194]}
   );
   gpc615_5 gpc1071 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[468]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[115],stage1_27[154],stage1_26[165],stage1_25[195]}
   );
   gpc615_5 gpc1072 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[469]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[116],stage1_27[155],stage1_26[166],stage1_25[196]}
   );
   gpc615_5 gpc1073 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[470]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[117],stage1_27[156],stage1_26[167],stage1_25[197]}
   );
   gpc615_5 gpc1074 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[471]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[118],stage1_27[157],stage1_26[168],stage1_25[198]}
   );
   gpc615_5 gpc1075 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[472]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[119],stage1_27[158],stage1_26[169],stage1_25[199]}
   );
   gpc615_5 gpc1076 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[473]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[120],stage1_27[159],stage1_26[170],stage1_25[200]}
   );
   gpc615_5 gpc1077 (
      {stage0_25[486], stage0_25[487], stage0_25[488], stage0_25[489], stage0_25[490]},
      {stage0_26[474]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[121],stage1_27[160],stage1_26[171],stage1_25[201]}
   );
   gpc615_5 gpc1078 (
      {stage0_25[491], stage0_25[492], stage0_25[493], stage0_25[494], stage0_25[495]},
      {stage0_26[475]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[122],stage1_27[161],stage1_26[172],stage1_25[202]}
   );
   gpc615_5 gpc1079 (
      {stage0_25[496], stage0_25[497], stage0_25[498], stage0_25[499], stage0_25[500]},
      {stage0_26[476]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[123],stage1_27[162],stage1_26[173],stage1_25[203]}
   );
   gpc615_5 gpc1080 (
      {stage0_25[501], stage0_25[502], stage0_25[503], stage0_25[504], stage0_25[505]},
      {stage0_26[477]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[124],stage1_27[163],stage1_26[174],stage1_25[204]}
   );
   gpc615_5 gpc1081 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[324]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[54],stage1_28[125],stage1_27[164],stage1_26[175]}
   );
   gpc615_5 gpc1082 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[325]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[55],stage1_28[126],stage1_27[165],stage1_26[176]}
   );
   gpc615_5 gpc1083 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[326]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[56],stage1_28[127],stage1_27[166],stage1_26[177]}
   );
   gpc615_5 gpc1084 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[327]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[57],stage1_28[128],stage1_27[167],stage1_26[178]}
   );
   gpc615_5 gpc1085 (
      {stage0_26[498], stage0_26[499], stage0_26[500], stage0_26[501], stage0_26[502]},
      {stage0_27[328]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[58],stage1_28[129],stage1_27[168],stage1_26[179]}
   );
   gpc7_3 gpc1086 (
      {stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[59],stage1_28[130],stage1_27[169]}
   );
   gpc7_3 gpc1087 (
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage1_29[60],stage1_28[131],stage1_27[170]}
   );
   gpc615_5 gpc1088 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[30]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[61],stage1_28[132],stage1_27[171]}
   );
   gpc615_5 gpc1089 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[31]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[62],stage1_28[133],stage1_27[172]}
   );
   gpc615_5 gpc1090 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[32]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[63],stage1_28[134],stage1_27[173]}
   );
   gpc615_5 gpc1091 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[33]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[64],stage1_28[135],stage1_27[174]}
   );
   gpc615_5 gpc1092 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[34]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[65],stage1_28[136],stage1_27[175]}
   );
   gpc615_5 gpc1093 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[35]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[66],stage1_28[137],stage1_27[176]}
   );
   gpc615_5 gpc1094 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[36]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[67],stage1_28[138],stage1_27[177]}
   );
   gpc615_5 gpc1095 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[37]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[68],stage1_28[139],stage1_27[178]}
   );
   gpc615_5 gpc1096 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[38]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[69],stage1_28[140],stage1_27[179]}
   );
   gpc615_5 gpc1097 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[39]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[70],stage1_28[141],stage1_27[180]}
   );
   gpc615_5 gpc1098 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[40]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[15],stage1_29[71],stage1_28[142],stage1_27[181]}
   );
   gpc615_5 gpc1099 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[41]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[16],stage1_29[72],stage1_28[143],stage1_27[182]}
   );
   gpc615_5 gpc1100 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[42]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[17],stage1_29[73],stage1_28[144],stage1_27[183]}
   );
   gpc615_5 gpc1101 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[43]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[18],stage1_29[74],stage1_28[145],stage1_27[184]}
   );
   gpc615_5 gpc1102 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[44]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[19],stage1_29[75],stage1_28[146],stage1_27[185]}
   );
   gpc615_5 gpc1103 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[45]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[20],stage1_29[76],stage1_28[147],stage1_27[186]}
   );
   gpc615_5 gpc1104 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[46]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[21],stage1_29[77],stage1_28[148],stage1_27[187]}
   );
   gpc615_5 gpc1105 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[47]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[22],stage1_29[78],stage1_28[149],stage1_27[188]}
   );
   gpc615_5 gpc1106 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[48]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[23],stage1_29[79],stage1_28[150],stage1_27[189]}
   );
   gpc615_5 gpc1107 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[49]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[24],stage1_29[80],stage1_28[151],stage1_27[190]}
   );
   gpc615_5 gpc1108 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[50]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[25],stage1_29[81],stage1_28[152],stage1_27[191]}
   );
   gpc615_5 gpc1109 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[51]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[26],stage1_29[82],stage1_28[153],stage1_27[192]}
   );
   gpc615_5 gpc1110 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[52]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[27],stage1_29[83],stage1_28[154],stage1_27[193]}
   );
   gpc615_5 gpc1111 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[53]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[28],stage1_29[84],stage1_28[155],stage1_27[194]}
   );
   gpc615_5 gpc1112 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[54]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[29],stage1_29[85],stage1_28[156],stage1_27[195]}
   );
   gpc615_5 gpc1113 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[55]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[30],stage1_29[86],stage1_28[157],stage1_27[196]}
   );
   gpc615_5 gpc1114 (
      {stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477]},
      {stage0_28[56]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[31],stage1_29[87],stage1_28[158],stage1_27[197]}
   );
   gpc615_5 gpc1115 (
      {stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_28[57]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[32],stage1_29[88],stage1_28[159],stage1_27[198]}
   );
   gpc615_5 gpc1116 (
      {stage0_27[483], stage0_27[484], stage0_27[485], stage0_27[486], stage0_27[487]},
      {stage0_28[58]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[33],stage1_29[89],stage1_28[160],stage1_27[199]}
   );
   gpc615_5 gpc1117 (
      {stage0_27[488], stage0_27[489], stage0_27[490], stage0_27[491], stage0_27[492]},
      {stage0_28[59]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[34],stage1_29[90],stage1_28[161],stage1_27[200]}
   );
   gpc615_5 gpc1118 (
      {stage0_27[493], stage0_27[494], stage0_27[495], stage0_27[496], stage0_27[497]},
      {stage0_28[60]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[35],stage1_29[91],stage1_28[162],stage1_27[201]}
   );
   gpc615_5 gpc1119 (
      {stage0_27[498], stage0_27[499], stage0_27[500], stage0_27[501], stage0_27[502]},
      {stage0_28[61]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[36],stage1_29[92],stage1_28[163],stage1_27[202]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65], stage0_28[66], stage0_28[67]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[32],stage1_30[37],stage1_29[93],stage1_28[164]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71], stage0_28[72], stage0_28[73]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[33],stage1_30[38],stage1_29[94],stage1_28[165]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78], stage0_28[79]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[34],stage1_30[39],stage1_29[95],stage1_28[166]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84], stage0_28[85]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[35],stage1_30[40],stage1_29[96],stage1_28[167]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90], stage0_28[91]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[36],stage1_30[41],stage1_29[97],stage1_28[168]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[37],stage1_30[42],stage1_29[98],stage1_28[169]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[38],stage1_30[43],stage1_29[99],stage1_28[170]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[39],stage1_30[44],stage1_29[100],stage1_28[171]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[40],stage1_30[45],stage1_29[101],stage1_28[172]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[41],stage1_30[46],stage1_29[102],stage1_28[173]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[42],stage1_30[47],stage1_29[103],stage1_28[174]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[43],stage1_30[48],stage1_29[104],stage1_28[175]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[44],stage1_30[49],stage1_29[105],stage1_28[176]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144], stage0_28[145]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[45],stage1_30[50],stage1_29[106],stage1_28[177]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150], stage0_28[151]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[46],stage1_30[51],stage1_29[107],stage1_28[178]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156], stage0_28[157]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[47],stage1_30[52],stage1_29[108],stage1_28[179]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162], stage0_28[163]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[48],stage1_30[53],stage1_29[109],stage1_28[180]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168], stage0_28[169]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[49],stage1_30[54],stage1_29[110],stage1_28[181]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174], stage0_28[175]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[50],stage1_30[55],stage1_29[111],stage1_28[182]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180], stage0_28[181]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[51],stage1_30[56],stage1_29[112],stage1_28[183]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186], stage0_28[187]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[52],stage1_30[57],stage1_29[113],stage1_28[184]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192], stage0_28[193]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[53],stage1_30[58],stage1_29[114],stage1_28[185]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198], stage0_28[199]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[54],stage1_30[59],stage1_29[115],stage1_28[186]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204], stage0_28[205]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[55],stage1_30[60],stage1_29[116],stage1_28[187]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210], stage0_28[211]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[56],stage1_30[61],stage1_29[117],stage1_28[188]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216], stage0_28[217]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[57],stage1_30[62],stage1_29[118],stage1_28[189]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222], stage0_28[223]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[58],stage1_30[63],stage1_29[119],stage1_28[190]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228], stage0_28[229]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[59],stage1_30[64],stage1_29[120],stage1_28[191]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234], stage0_28[235]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[60],stage1_30[65],stage1_29[121],stage1_28[192]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240], stage0_28[241]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[61],stage1_30[66],stage1_29[122],stage1_28[193]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246], stage0_28[247]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[62],stage1_30[67],stage1_29[123],stage1_28[194]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252], stage0_28[253]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[63],stage1_30[68],stage1_29[124],stage1_28[195]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258], stage0_28[259]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[64],stage1_30[69],stage1_29[125],stage1_28[196]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264], stage0_28[265]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[65],stage1_30[70],stage1_29[126],stage1_28[197]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270], stage0_28[271]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[66],stage1_30[71],stage1_29[127],stage1_28[198]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276], stage0_28[277]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[67],stage1_30[72],stage1_29[128],stage1_28[199]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282], stage0_28[283]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[68],stage1_30[73],stage1_29[129],stage1_28[200]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288], stage0_28[289]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[69],stage1_30[74],stage1_29[130],stage1_28[201]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294], stage0_28[295]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[70],stage1_30[75],stage1_29[131],stage1_28[202]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300], stage0_28[301]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[71],stage1_30[76],stage1_29[132],stage1_28[203]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306], stage0_28[307]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[72],stage1_30[77],stage1_29[133],stage1_28[204]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312], stage0_28[313]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[73],stage1_30[78],stage1_29[134],stage1_28[205]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[74],stage1_30[79],stage1_29[135],stage1_28[206]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[75],stage1_30[80],stage1_29[136],stage1_28[207]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330], stage0_28[331]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[76],stage1_30[81],stage1_29[137],stage1_28[208]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336], stage0_28[337]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[77],stage1_30[82],stage1_29[138],stage1_28[209]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342], stage0_28[343]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[78],stage1_30[83],stage1_29[139],stage1_28[210]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[79],stage1_30[84],stage1_29[140],stage1_28[211]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[80],stage1_30[85],stage1_29[141],stage1_28[212]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360], stage0_28[361]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[81],stage1_30[86],stage1_29[142],stage1_28[213]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366], stage0_28[367]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[82],stage1_30[87],stage1_29[143],stage1_28[214]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372], stage0_28[373]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[83],stage1_30[88],stage1_29[144],stage1_28[215]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[84],stage1_30[89],stage1_29[145],stage1_28[216]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[85],stage1_30[90],stage1_29[146],stage1_28[217]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390], stage0_28[391]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[86],stage1_30[91],stage1_29[147],stage1_28[218]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396], stage0_28[397]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[87],stage1_30[92],stage1_29[148],stage1_28[219]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402], stage0_28[403]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[88],stage1_30[93],stage1_29[149],stage1_28[220]}
   );
   gpc606_5 gpc1177 (
      {stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[89],stage1_30[94],stage1_29[150],stage1_28[221]}
   );
   gpc606_5 gpc1178 (
      {stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[90],stage1_30[95],stage1_29[151],stage1_28[222]}
   );
   gpc606_5 gpc1179 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420], stage0_28[421]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[91],stage1_30[96],stage1_29[152],stage1_28[223]}
   );
   gpc606_5 gpc1180 (
      {stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426], stage0_28[427]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[92],stage1_30[97],stage1_29[153],stage1_28[224]}
   );
   gpc606_5 gpc1181 (
      {stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432], stage0_28[433]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[93],stage1_30[98],stage1_29[154],stage1_28[225]}
   );
   gpc606_5 gpc1182 (
      {stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[94],stage1_30[99],stage1_29[155],stage1_28[226]}
   );
   gpc606_5 gpc1183 (
      {stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[95],stage1_30[100],stage1_29[156],stage1_28[227]}
   );
   gpc606_5 gpc1184 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450], stage0_28[451]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[96],stage1_30[101],stage1_29[157],stage1_28[228]}
   );
   gpc606_5 gpc1185 (
      {stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456], stage0_28[457]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[97],stage1_30[102],stage1_29[158],stage1_28[229]}
   );
   gpc606_5 gpc1186 (
      {stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462], stage0_28[463]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[98],stage1_30[103],stage1_29[159],stage1_28[230]}
   );
   gpc606_5 gpc1187 (
      {stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[99],stage1_30[104],stage1_29[160],stage1_28[231]}
   );
   gpc606_5 gpc1188 (
      {stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[100],stage1_30[105],stage1_29[161],stage1_28[232]}
   );
   gpc606_5 gpc1189 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480], stage0_28[481]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[101],stage1_30[106],stage1_29[162],stage1_28[233]}
   );
   gpc606_5 gpc1190 (
      {stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485], stage0_28[486], stage0_28[487]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[102],stage1_30[107],stage1_29[163],stage1_28[234]}
   );
   gpc606_5 gpc1191 (
      {stage0_28[488], stage0_28[489], stage0_28[490], stage0_28[491], stage0_28[492], stage0_28[493]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[103],stage1_30[108],stage1_29[164],stage1_28[235]}
   );
   gpc606_5 gpc1192 (
      {stage0_28[494], stage0_28[495], stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[104],stage1_30[109],stage1_29[165],stage1_28[236]}
   );
   gpc606_5 gpc1193 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[73],stage1_31[105],stage1_30[110],stage1_29[166]}
   );
   gpc606_5 gpc1194 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[74],stage1_31[106],stage1_30[111],stage1_29[167]}
   );
   gpc606_5 gpc1195 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[75],stage1_31[107],stage1_30[112],stage1_29[168]}
   );
   gpc606_5 gpc1196 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[76],stage1_31[108],stage1_30[113],stage1_29[169]}
   );
   gpc606_5 gpc1197 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[77],stage1_31[109],stage1_30[114],stage1_29[170]}
   );
   gpc606_5 gpc1198 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[78],stage1_31[110],stage1_30[115],stage1_29[171]}
   );
   gpc606_5 gpc1199 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[79],stage1_31[111],stage1_30[116],stage1_29[172]}
   );
   gpc606_5 gpc1200 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[80],stage1_31[112],stage1_30[117],stage1_29[173]}
   );
   gpc606_5 gpc1201 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[81],stage1_31[113],stage1_30[118],stage1_29[174]}
   );
   gpc606_5 gpc1202 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[82],stage1_31[114],stage1_30[119],stage1_29[175]}
   );
   gpc606_5 gpc1203 (
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[83],stage1_31[115],stage1_30[120],stage1_29[176]}
   );
   gpc606_5 gpc1204 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[84],stage1_31[116],stage1_30[121],stage1_29[177]}
   );
   gpc606_5 gpc1205 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[85],stage1_31[117],stage1_30[122],stage1_29[178]}
   );
   gpc606_5 gpc1206 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[86],stage1_31[118],stage1_30[123],stage1_29[179]}
   );
   gpc606_5 gpc1207 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[87],stage1_31[119],stage1_30[124],stage1_29[180]}
   );
   gpc606_5 gpc1208 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[88],stage1_31[120],stage1_30[125],stage1_29[181]}
   );
   gpc606_5 gpc1209 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[89],stage1_31[121],stage1_30[126],stage1_29[182]}
   );
   gpc606_5 gpc1210 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[90],stage1_31[122],stage1_30[127],stage1_29[183]}
   );
   gpc606_5 gpc1211 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[91],stage1_31[123],stage1_30[128],stage1_29[184]}
   );
   gpc606_5 gpc1212 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[92],stage1_31[124],stage1_30[129],stage1_29[185]}
   );
   gpc606_5 gpc1213 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[93],stage1_31[125],stage1_30[130],stage1_29[186]}
   );
   gpc606_5 gpc1214 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[94],stage1_31[126],stage1_30[131],stage1_29[187]}
   );
   gpc606_5 gpc1215 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[95],stage1_31[127],stage1_30[132],stage1_29[188]}
   );
   gpc606_5 gpc1216 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[96],stage1_31[128],stage1_30[133],stage1_29[189]}
   );
   gpc606_5 gpc1217 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[97],stage1_31[129],stage1_30[134],stage1_29[190]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[98],stage1_31[130],stage1_30[135],stage1_29[191]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[99],stage1_31[131],stage1_30[136],stage1_29[192]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[100],stage1_31[132],stage1_30[137],stage1_29[193]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[101],stage1_31[133],stage1_30[138],stage1_29[194]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[102],stage1_31[134],stage1_30[139],stage1_29[195]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[103],stage1_31[135],stage1_30[140],stage1_29[196]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[104],stage1_31[136],stage1_30[141],stage1_29[197]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[105],stage1_31[137],stage1_30[142],stage1_29[198]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[106],stage1_31[138],stage1_30[143],stage1_29[199]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[107],stage1_31[139],stage1_30[144],stage1_29[200]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[108],stage1_31[140],stage1_30[145],stage1_29[201]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[109],stage1_31[141],stage1_30[146],stage1_29[202]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[110],stage1_31[142],stage1_30[147],stage1_29[203]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[111],stage1_31[143],stage1_30[148],stage1_29[204]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[112],stage1_31[144],stage1_30[149],stage1_29[205]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[113],stage1_31[145],stage1_30[150],stage1_29[206]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[114],stage1_31[146],stage1_30[151],stage1_29[207]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[115],stage1_31[147],stage1_30[152],stage1_29[208]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[116],stage1_31[148],stage1_30[153],stage1_29[209]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460], stage0_29[461]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[117],stage1_31[149],stage1_30[154],stage1_29[210]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466], stage0_29[467]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[118],stage1_31[150],stage1_30[155],stage1_29[211]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472], stage0_29[473]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[119],stage1_31[151],stage1_30[156],stage1_29[212]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[120],stage1_31[152],stage1_30[157],stage1_29[213]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[121],stage1_31[153],stage1_30[158],stage1_29[214]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490], stage0_29[491]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[122],stage1_31[154],stage1_30[159],stage1_29[215]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496], stage0_29[497]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[123],stage1_31[155],stage1_30[160],stage1_29[216]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502], stage0_29[503]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[124],stage1_31[156],stage1_30[161],stage1_29[217]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508], stage0_29[509]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[125],stage1_31[157],stage1_30[162],stage1_29[218]}
   );
   gpc1415_5 gpc1246 (
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442]},
      {stage0_31[318]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[53],stage1_32[126],stage1_31[158],stage1_30[163]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage0_32[4]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[1],stage1_33[54],stage1_32[127],stage1_31[159]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328]},
      {stage0_32[5]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[2],stage1_33[55],stage1_32[128],stage1_31[160]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[329], stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333]},
      {stage0_32[6]},
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage1_35[2],stage1_34[3],stage1_33[56],stage1_32[129],stage1_31[161]}
   );
   gpc615_5 gpc1250 (
      {stage0_31[334], stage0_31[335], stage0_31[336], stage0_31[337], stage0_31[338]},
      {stage0_32[7]},
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage1_35[3],stage1_34[4],stage1_33[57],stage1_32[130],stage1_31[162]}
   );
   gpc615_5 gpc1251 (
      {stage0_31[339], stage0_31[340], stage0_31[341], stage0_31[342], stage0_31[343]},
      {stage0_32[8]},
      {stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29], stage0_33[30]},
      {stage1_35[4],stage1_34[5],stage1_33[58],stage1_32[131],stage1_31[163]}
   );
   gpc615_5 gpc1252 (
      {stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347], stage0_31[348]},
      {stage0_32[9]},
      {stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35], stage0_33[36]},
      {stage1_35[5],stage1_34[6],stage1_33[59],stage1_32[132],stage1_31[164]}
   );
   gpc615_5 gpc1253 (
      {stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage0_32[10]},
      {stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41], stage0_33[42]},
      {stage1_35[6],stage1_34[7],stage1_33[60],stage1_32[133],stage1_31[165]}
   );
   gpc615_5 gpc1254 (
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358]},
      {stage0_32[11]},
      {stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47], stage0_33[48]},
      {stage1_35[7],stage1_34[8],stage1_33[61],stage1_32[134],stage1_31[166]}
   );
   gpc615_5 gpc1255 (
      {stage0_31[359], stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363]},
      {stage0_32[12]},
      {stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53], stage0_33[54]},
      {stage1_35[8],stage1_34[9],stage1_33[62],stage1_32[135],stage1_31[167]}
   );
   gpc615_5 gpc1256 (
      {stage0_31[364], stage0_31[365], stage0_31[366], stage0_31[367], stage0_31[368]},
      {stage0_32[13]},
      {stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59], stage0_33[60]},
      {stage1_35[9],stage1_34[10],stage1_33[63],stage1_32[136],stage1_31[168]}
   );
   gpc615_5 gpc1257 (
      {stage0_31[369], stage0_31[370], stage0_31[371], stage0_31[372], stage0_31[373]},
      {stage0_32[14]},
      {stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65], stage0_33[66]},
      {stage1_35[10],stage1_34[11],stage1_33[64],stage1_32[137],stage1_31[169]}
   );
   gpc615_5 gpc1258 (
      {stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377], stage0_31[378]},
      {stage0_32[15]},
      {stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71], stage0_33[72]},
      {stage1_35[11],stage1_34[12],stage1_33[65],stage1_32[138],stage1_31[170]}
   );
   gpc615_5 gpc1259 (
      {stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage0_32[16]},
      {stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77], stage0_33[78]},
      {stage1_35[12],stage1_34[13],stage1_33[66],stage1_32[139],stage1_31[171]}
   );
   gpc615_5 gpc1260 (
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388]},
      {stage0_32[17]},
      {stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83], stage0_33[84]},
      {stage1_35[13],stage1_34[14],stage1_33[67],stage1_32[140],stage1_31[172]}
   );
   gpc615_5 gpc1261 (
      {stage0_31[389], stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393]},
      {stage0_32[18]},
      {stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89], stage0_33[90]},
      {stage1_35[14],stage1_34[15],stage1_33[68],stage1_32[141],stage1_31[173]}
   );
   gpc615_5 gpc1262 (
      {stage0_31[394], stage0_31[395], stage0_31[396], stage0_31[397], stage0_31[398]},
      {stage0_32[19]},
      {stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95], stage0_33[96]},
      {stage1_35[15],stage1_34[16],stage1_33[69],stage1_32[142],stage1_31[174]}
   );
   gpc615_5 gpc1263 (
      {stage0_31[399], stage0_31[400], stage0_31[401], stage0_31[402], stage0_31[403]},
      {stage0_32[20]},
      {stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101], stage0_33[102]},
      {stage1_35[16],stage1_34[17],stage1_33[70],stage1_32[143],stage1_31[175]}
   );
   gpc615_5 gpc1264 (
      {stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407], stage0_31[408]},
      {stage0_32[21]},
      {stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107], stage0_33[108]},
      {stage1_35[17],stage1_34[18],stage1_33[71],stage1_32[144],stage1_31[176]}
   );
   gpc615_5 gpc1265 (
      {stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage0_32[22]},
      {stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113], stage0_33[114]},
      {stage1_35[18],stage1_34[19],stage1_33[72],stage1_32[145],stage1_31[177]}
   );
   gpc615_5 gpc1266 (
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418]},
      {stage0_32[23]},
      {stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119], stage0_33[120]},
      {stage1_35[19],stage1_34[20],stage1_33[73],stage1_32[146],stage1_31[178]}
   );
   gpc615_5 gpc1267 (
      {stage0_31[419], stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423]},
      {stage0_32[24]},
      {stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125], stage0_33[126]},
      {stage1_35[20],stage1_34[21],stage1_33[74],stage1_32[147],stage1_31[179]}
   );
   gpc615_5 gpc1268 (
      {stage0_31[424], stage0_31[425], stage0_31[426], stage0_31[427], stage0_31[428]},
      {stage0_32[25]},
      {stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131], stage0_33[132]},
      {stage1_35[21],stage1_34[22],stage1_33[75],stage1_32[148],stage1_31[180]}
   );
   gpc615_5 gpc1269 (
      {stage0_31[429], stage0_31[430], stage0_31[431], stage0_31[432], stage0_31[433]},
      {stage0_32[26]},
      {stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137], stage0_33[138]},
      {stage1_35[22],stage1_34[23],stage1_33[76],stage1_32[149],stage1_31[181]}
   );
   gpc615_5 gpc1270 (
      {stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437], stage0_31[438]},
      {stage0_32[27]},
      {stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143], stage0_33[144]},
      {stage1_35[23],stage1_34[24],stage1_33[77],stage1_32[150],stage1_31[182]}
   );
   gpc615_5 gpc1271 (
      {stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage0_32[28]},
      {stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149], stage0_33[150]},
      {stage1_35[24],stage1_34[25],stage1_33[78],stage1_32[151],stage1_31[183]}
   );
   gpc615_5 gpc1272 (
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448]},
      {stage0_32[29]},
      {stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155], stage0_33[156]},
      {stage1_35[25],stage1_34[26],stage1_33[79],stage1_32[152],stage1_31[184]}
   );
   gpc615_5 gpc1273 (
      {stage0_31[449], stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453]},
      {stage0_32[30]},
      {stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161], stage0_33[162]},
      {stage1_35[26],stage1_34[27],stage1_33[80],stage1_32[153],stage1_31[185]}
   );
   gpc615_5 gpc1274 (
      {stage0_31[454], stage0_31[455], stage0_31[456], stage0_31[457], stage0_31[458]},
      {stage0_32[31]},
      {stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167], stage0_33[168]},
      {stage1_35[27],stage1_34[28],stage1_33[81],stage1_32[154],stage1_31[186]}
   );
   gpc615_5 gpc1275 (
      {stage0_31[459], stage0_31[460], stage0_31[461], stage0_31[462], stage0_31[463]},
      {stage0_32[32]},
      {stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173], stage0_33[174]},
      {stage1_35[28],stage1_34[29],stage1_33[82],stage1_32[155],stage1_31[187]}
   );
   gpc615_5 gpc1276 (
      {stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467], stage0_31[468]},
      {stage0_32[33]},
      {stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179], stage0_33[180]},
      {stage1_35[29],stage1_34[30],stage1_33[83],stage1_32[156],stage1_31[188]}
   );
   gpc615_5 gpc1277 (
      {stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage0_32[34]},
      {stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185], stage0_33[186]},
      {stage1_35[30],stage1_34[31],stage1_33[84],stage1_32[157],stage1_31[189]}
   );
   gpc615_5 gpc1278 (
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478]},
      {stage0_32[35]},
      {stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191], stage0_33[192]},
      {stage1_35[31],stage1_34[32],stage1_33[85],stage1_32[158],stage1_31[190]}
   );
   gpc615_5 gpc1279 (
      {stage0_31[479], stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483]},
      {stage0_32[36]},
      {stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197], stage0_33[198]},
      {stage1_35[32],stage1_34[33],stage1_33[86],stage1_32[159],stage1_31[191]}
   );
   gpc615_5 gpc1280 (
      {stage0_31[484], stage0_31[485], stage0_31[486], stage0_31[487], stage0_31[488]},
      {stage0_32[37]},
      {stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203], stage0_33[204]},
      {stage1_35[33],stage1_34[34],stage1_33[87],stage1_32[160],stage1_31[192]}
   );
   gpc615_5 gpc1281 (
      {stage0_31[489], stage0_31[490], stage0_31[491], stage0_31[492], stage0_31[493]},
      {stage0_32[38]},
      {stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209], stage0_33[210]},
      {stage1_35[34],stage1_34[35],stage1_33[88],stage1_32[161],stage1_31[193]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[35],stage1_34[36],stage1_33[89],stage1_32[162]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[36],stage1_34[37],stage1_33[90],stage1_32[163]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[37],stage1_34[38],stage1_33[91],stage1_32[164]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[38],stage1_34[39],stage1_33[92],stage1_32[165]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[63], stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[39],stage1_34[40],stage1_33[93],stage1_32[166]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73], stage0_32[74]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[40],stage1_34[41],stage1_33[94],stage1_32[167]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78], stage0_32[79], stage0_32[80]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[41],stage1_34[42],stage1_33[95],stage1_32[168]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[81], stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[42],stage1_34[43],stage1_33[96],stage1_32[169]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[87], stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[43],stage1_34[44],stage1_33[97],stage1_32[170]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[93], stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[44],stage1_34[45],stage1_33[98],stage1_32[171]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103], stage0_32[104]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[45],stage1_34[46],stage1_33[99],stage1_32[172]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108], stage0_32[109], stage0_32[110]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[46],stage1_34[47],stage1_33[100],stage1_32[173]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[111], stage0_32[112], stage0_32[113], stage0_32[114], stage0_32[115], stage0_32[116]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[47],stage1_34[48],stage1_33[101],stage1_32[174]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[117], stage0_32[118], stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[48],stage1_34[49],stage1_33[102],stage1_32[175]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[123], stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[49],stage1_34[50],stage1_33[103],stage1_32[176]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[129], stage0_32[130], stage0_32[131], stage0_32[132], stage0_32[133], stage0_32[134]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[50],stage1_34[51],stage1_33[104],stage1_32[177]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[135], stage0_32[136], stage0_32[137], stage0_32[138], stage0_32[139], stage0_32[140]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[51],stage1_34[52],stage1_33[105],stage1_32[178]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[141], stage0_32[142], stage0_32[143], stage0_32[144], stage0_32[145], stage0_32[146]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[52],stage1_34[53],stage1_33[106],stage1_32[179]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[147], stage0_32[148], stage0_32[149], stage0_32[150], stage0_32[151], stage0_32[152]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[53],stage1_34[54],stage1_33[107],stage1_32[180]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[153], stage0_32[154], stage0_32[155], stage0_32[156], stage0_32[157], stage0_32[158]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[54],stage1_34[55],stage1_33[108],stage1_32[181]}
   );
   gpc606_5 gpc1302 (
      {stage0_32[159], stage0_32[160], stage0_32[161], stage0_32[162], stage0_32[163], stage0_32[164]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[55],stage1_34[56],stage1_33[109],stage1_32[182]}
   );
   gpc606_5 gpc1303 (
      {stage0_32[165], stage0_32[166], stage0_32[167], stage0_32[168], stage0_32[169], stage0_32[170]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[56],stage1_34[57],stage1_33[110],stage1_32[183]}
   );
   gpc606_5 gpc1304 (
      {stage0_32[171], stage0_32[172], stage0_32[173], stage0_32[174], stage0_32[175], stage0_32[176]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[57],stage1_34[58],stage1_33[111],stage1_32[184]}
   );
   gpc606_5 gpc1305 (
      {stage0_32[177], stage0_32[178], stage0_32[179], stage0_32[180], stage0_32[181], stage0_32[182]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[58],stage1_34[59],stage1_33[112],stage1_32[185]}
   );
   gpc606_5 gpc1306 (
      {stage0_32[183], stage0_32[184], stage0_32[185], stage0_32[186], stage0_32[187], stage0_32[188]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[59],stage1_34[60],stage1_33[113],stage1_32[186]}
   );
   gpc606_5 gpc1307 (
      {stage0_32[189], stage0_32[190], stage0_32[191], stage0_32[192], stage0_32[193], stage0_32[194]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[60],stage1_34[61],stage1_33[114],stage1_32[187]}
   );
   gpc606_5 gpc1308 (
      {stage0_32[195], stage0_32[196], stage0_32[197], stage0_32[198], stage0_32[199], stage0_32[200]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[61],stage1_34[62],stage1_33[115],stage1_32[188]}
   );
   gpc606_5 gpc1309 (
      {stage0_32[201], stage0_32[202], stage0_32[203], stage0_32[204], stage0_32[205], stage0_32[206]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[62],stage1_34[63],stage1_33[116],stage1_32[189]}
   );
   gpc606_5 gpc1310 (
      {stage0_32[207], stage0_32[208], stage0_32[209], stage0_32[210], stage0_32[211], stage0_32[212]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[63],stage1_34[64],stage1_33[117],stage1_32[190]}
   );
   gpc606_5 gpc1311 (
      {stage0_32[213], stage0_32[214], stage0_32[215], stage0_32[216], stage0_32[217], stage0_32[218]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[64],stage1_34[65],stage1_33[118],stage1_32[191]}
   );
   gpc606_5 gpc1312 (
      {stage0_32[219], stage0_32[220], stage0_32[221], stage0_32[222], stage0_32[223], stage0_32[224]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[65],stage1_34[66],stage1_33[119],stage1_32[192]}
   );
   gpc606_5 gpc1313 (
      {stage0_32[225], stage0_32[226], stage0_32[227], stage0_32[228], stage0_32[229], stage0_32[230]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[66],stage1_34[67],stage1_33[120],stage1_32[193]}
   );
   gpc606_5 gpc1314 (
      {stage0_32[231], stage0_32[232], stage0_32[233], stage0_32[234], stage0_32[235], stage0_32[236]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[67],stage1_34[68],stage1_33[121],stage1_32[194]}
   );
   gpc606_5 gpc1315 (
      {stage0_32[237], stage0_32[238], stage0_32[239], stage0_32[240], stage0_32[241], stage0_32[242]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[68],stage1_34[69],stage1_33[122],stage1_32[195]}
   );
   gpc606_5 gpc1316 (
      {stage0_32[243], stage0_32[244], stage0_32[245], stage0_32[246], stage0_32[247], stage0_32[248]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[69],stage1_34[70],stage1_33[123],stage1_32[196]}
   );
   gpc606_5 gpc1317 (
      {stage0_32[249], stage0_32[250], stage0_32[251], stage0_32[252], stage0_32[253], stage0_32[254]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[70],stage1_34[71],stage1_33[124],stage1_32[197]}
   );
   gpc606_5 gpc1318 (
      {stage0_32[255], stage0_32[256], stage0_32[257], stage0_32[258], stage0_32[259], stage0_32[260]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[71],stage1_34[72],stage1_33[125],stage1_32[198]}
   );
   gpc606_5 gpc1319 (
      {stage0_32[261], stage0_32[262], stage0_32[263], stage0_32[264], stage0_32[265], stage0_32[266]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[72],stage1_34[73],stage1_33[126],stage1_32[199]}
   );
   gpc606_5 gpc1320 (
      {stage0_32[267], stage0_32[268], stage0_32[269], stage0_32[270], stage0_32[271], stage0_32[272]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[73],stage1_34[74],stage1_33[127],stage1_32[200]}
   );
   gpc606_5 gpc1321 (
      {stage0_32[273], stage0_32[274], stage0_32[275], stage0_32[276], stage0_32[277], stage0_32[278]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[74],stage1_34[75],stage1_33[128],stage1_32[201]}
   );
   gpc606_5 gpc1322 (
      {stage0_32[279], stage0_32[280], stage0_32[281], stage0_32[282], stage0_32[283], stage0_32[284]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[75],stage1_34[76],stage1_33[129],stage1_32[202]}
   );
   gpc606_5 gpc1323 (
      {stage0_32[285], stage0_32[286], stage0_32[287], stage0_32[288], stage0_32[289], stage0_32[290]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[76],stage1_34[77],stage1_33[130],stage1_32[203]}
   );
   gpc606_5 gpc1324 (
      {stage0_32[291], stage0_32[292], stage0_32[293], stage0_32[294], stage0_32[295], stage0_32[296]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[77],stage1_34[78],stage1_33[131],stage1_32[204]}
   );
   gpc606_5 gpc1325 (
      {stage0_32[297], stage0_32[298], stage0_32[299], stage0_32[300], stage0_32[301], stage0_32[302]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[78],stage1_34[79],stage1_33[132],stage1_32[205]}
   );
   gpc615_5 gpc1326 (
      {stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage0_34[264]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[44],stage1_35[79],stage1_34[80],stage1_33[133]}
   );
   gpc615_5 gpc1327 (
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220]},
      {stage0_34[265]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[45],stage1_35[80],stage1_34[81],stage1_33[134]}
   );
   gpc615_5 gpc1328 (
      {stage0_33[221], stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225]},
      {stage0_34[266]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[46],stage1_35[81],stage1_34[82],stage1_33[135]}
   );
   gpc615_5 gpc1329 (
      {stage0_33[226], stage0_33[227], stage0_33[228], stage0_33[229], stage0_33[230]},
      {stage0_34[267]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[47],stage1_35[82],stage1_34[83],stage1_33[136]}
   );
   gpc615_5 gpc1330 (
      {stage0_33[231], stage0_33[232], stage0_33[233], stage0_33[234], stage0_33[235]},
      {stage0_34[268]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[48],stage1_35[83],stage1_34[84],stage1_33[137]}
   );
   gpc615_5 gpc1331 (
      {stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239], stage0_33[240]},
      {stage0_34[269]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[49],stage1_35[84],stage1_34[85],stage1_33[138]}
   );
   gpc615_5 gpc1332 (
      {stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage0_34[270]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[50],stage1_35[85],stage1_34[86],stage1_33[139]}
   );
   gpc615_5 gpc1333 (
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250]},
      {stage0_34[271]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[51],stage1_35[86],stage1_34[87],stage1_33[140]}
   );
   gpc615_5 gpc1334 (
      {stage0_33[251], stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255]},
      {stage0_34[272]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[52],stage1_35[87],stage1_34[88],stage1_33[141]}
   );
   gpc615_5 gpc1335 (
      {stage0_33[256], stage0_33[257], stage0_33[258], stage0_33[259], stage0_33[260]},
      {stage0_34[273]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[53],stage1_35[88],stage1_34[89],stage1_33[142]}
   );
   gpc615_5 gpc1336 (
      {stage0_33[261], stage0_33[262], stage0_33[263], stage0_33[264], stage0_33[265]},
      {stage0_34[274]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[54],stage1_35[89],stage1_34[90],stage1_33[143]}
   );
   gpc615_5 gpc1337 (
      {stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269], stage0_33[270]},
      {stage0_34[275]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[55],stage1_35[90],stage1_34[91],stage1_33[144]}
   );
   gpc615_5 gpc1338 (
      {stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage0_34[276]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[56],stage1_35[91],stage1_34[92],stage1_33[145]}
   );
   gpc615_5 gpc1339 (
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280]},
      {stage0_34[277]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[57],stage1_35[92],stage1_34[93],stage1_33[146]}
   );
   gpc615_5 gpc1340 (
      {stage0_33[281], stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285]},
      {stage0_34[278]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[58],stage1_35[93],stage1_34[94],stage1_33[147]}
   );
   gpc615_5 gpc1341 (
      {stage0_33[286], stage0_33[287], stage0_33[288], stage0_33[289], stage0_33[290]},
      {stage0_34[279]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[59],stage1_35[94],stage1_34[95],stage1_33[148]}
   );
   gpc615_5 gpc1342 (
      {stage0_33[291], stage0_33[292], stage0_33[293], stage0_33[294], stage0_33[295]},
      {stage0_34[280]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[60],stage1_35[95],stage1_34[96],stage1_33[149]}
   );
   gpc615_5 gpc1343 (
      {stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299], stage0_33[300]},
      {stage0_34[281]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[61],stage1_35[96],stage1_34[97],stage1_33[150]}
   );
   gpc615_5 gpc1344 (
      {stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage0_34[282]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage1_37[18],stage1_36[62],stage1_35[97],stage1_34[98],stage1_33[151]}
   );
   gpc615_5 gpc1345 (
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310]},
      {stage0_34[283]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage1_37[19],stage1_36[63],stage1_35[98],stage1_34[99],stage1_33[152]}
   );
   gpc615_5 gpc1346 (
      {stage0_33[311], stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315]},
      {stage0_34[284]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage1_37[20],stage1_36[64],stage1_35[99],stage1_34[100],stage1_33[153]}
   );
   gpc615_5 gpc1347 (
      {stage0_33[316], stage0_33[317], stage0_33[318], stage0_33[319], stage0_33[320]},
      {stage0_34[285]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage1_37[21],stage1_36[65],stage1_35[100],stage1_34[101],stage1_33[154]}
   );
   gpc615_5 gpc1348 (
      {stage0_33[321], stage0_33[322], stage0_33[323], stage0_33[324], stage0_33[325]},
      {stage0_34[286]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage1_37[22],stage1_36[66],stage1_35[101],stage1_34[102],stage1_33[155]}
   );
   gpc615_5 gpc1349 (
      {stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329], stage0_33[330]},
      {stage0_34[287]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage1_37[23],stage1_36[67],stage1_35[102],stage1_34[103],stage1_33[156]}
   );
   gpc615_5 gpc1350 (
      {stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_34[288]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage1_37[24],stage1_36[68],stage1_35[103],stage1_34[104],stage1_33[157]}
   );
   gpc615_5 gpc1351 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340]},
      {stage0_34[289]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage1_37[25],stage1_36[69],stage1_35[104],stage1_34[105],stage1_33[158]}
   );
   gpc615_5 gpc1352 (
      {stage0_33[341], stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345]},
      {stage0_34[290]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage1_37[26],stage1_36[70],stage1_35[105],stage1_34[106],stage1_33[159]}
   );
   gpc615_5 gpc1353 (
      {stage0_33[346], stage0_33[347], stage0_33[348], stage0_33[349], stage0_33[350]},
      {stage0_34[291]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage1_37[27],stage1_36[71],stage1_35[106],stage1_34[107],stage1_33[160]}
   );
   gpc615_5 gpc1354 (
      {stage0_33[351], stage0_33[352], stage0_33[353], stage0_33[354], stage0_33[355]},
      {stage0_34[292]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage1_37[28],stage1_36[72],stage1_35[107],stage1_34[108],stage1_33[161]}
   );
   gpc615_5 gpc1355 (
      {stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359], stage0_33[360]},
      {stage0_34[293]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage1_37[29],stage1_36[73],stage1_35[108],stage1_34[109],stage1_33[162]}
   );
   gpc615_5 gpc1356 (
      {stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_34[294]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage1_37[30],stage1_36[74],stage1_35[109],stage1_34[110],stage1_33[163]}
   );
   gpc615_5 gpc1357 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370]},
      {stage0_34[295]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage1_37[31],stage1_36[75],stage1_35[110],stage1_34[111],stage1_33[164]}
   );
   gpc615_5 gpc1358 (
      {stage0_33[371], stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375]},
      {stage0_34[296]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage1_37[32],stage1_36[76],stage1_35[111],stage1_34[112],stage1_33[165]}
   );
   gpc615_5 gpc1359 (
      {stage0_33[376], stage0_33[377], stage0_33[378], stage0_33[379], stage0_33[380]},
      {stage0_34[297]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage1_37[33],stage1_36[77],stage1_35[112],stage1_34[113],stage1_33[166]}
   );
   gpc615_5 gpc1360 (
      {stage0_33[381], stage0_33[382], stage0_33[383], stage0_33[384], stage0_33[385]},
      {stage0_34[298]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage1_37[34],stage1_36[78],stage1_35[113],stage1_34[114],stage1_33[167]}
   );
   gpc615_5 gpc1361 (
      {stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389], stage0_33[390]},
      {stage0_34[299]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage1_37[35],stage1_36[79],stage1_35[114],stage1_34[115],stage1_33[168]}
   );
   gpc615_5 gpc1362 (
      {stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_34[300]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage1_37[36],stage1_36[80],stage1_35[115],stage1_34[116],stage1_33[169]}
   );
   gpc615_5 gpc1363 (
      {stage0_33[396], stage0_33[397], stage0_33[398], stage0_33[399], stage0_33[400]},
      {stage0_34[301]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage1_37[37],stage1_36[81],stage1_35[116],stage1_34[117],stage1_33[170]}
   );
   gpc615_5 gpc1364 (
      {stage0_33[401], stage0_33[402], stage0_33[403], stage0_33[404], stage0_33[405]},
      {stage0_34[302]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage1_37[38],stage1_36[82],stage1_35[117],stage1_34[118],stage1_33[171]}
   );
   gpc615_5 gpc1365 (
      {stage0_33[406], stage0_33[407], stage0_33[408], stage0_33[409], stage0_33[410]},
      {stage0_34[303]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage1_37[39],stage1_36[83],stage1_35[118],stage1_34[119],stage1_33[172]}
   );
   gpc615_5 gpc1366 (
      {stage0_33[411], stage0_33[412], stage0_33[413], stage0_33[414], stage0_33[415]},
      {stage0_34[304]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage1_37[40],stage1_36[84],stage1_35[119],stage1_34[120],stage1_33[173]}
   );
   gpc615_5 gpc1367 (
      {stage0_33[416], stage0_33[417], stage0_33[418], stage0_33[419], stage0_33[420]},
      {stage0_34[305]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage1_37[41],stage1_36[85],stage1_35[120],stage1_34[121],stage1_33[174]}
   );
   gpc615_5 gpc1368 (
      {stage0_33[421], stage0_33[422], stage0_33[423], stage0_33[424], stage0_33[425]},
      {stage0_34[306]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage1_37[42],stage1_36[86],stage1_35[121],stage1_34[122],stage1_33[175]}
   );
   gpc615_5 gpc1369 (
      {stage0_33[426], stage0_33[427], stage0_33[428], stage0_33[429], stage0_33[430]},
      {stage0_34[307]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage1_37[43],stage1_36[87],stage1_35[122],stage1_34[123],stage1_33[176]}
   );
   gpc615_5 gpc1370 (
      {stage0_33[431], stage0_33[432], stage0_33[433], stage0_33[434], stage0_33[435]},
      {stage0_34[308]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage1_37[44],stage1_36[88],stage1_35[123],stage1_34[124],stage1_33[177]}
   );
   gpc615_5 gpc1371 (
      {stage0_33[436], stage0_33[437], stage0_33[438], stage0_33[439], stage0_33[440]},
      {stage0_34[309]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage1_37[45],stage1_36[89],stage1_35[124],stage1_34[125],stage1_33[178]}
   );
   gpc615_5 gpc1372 (
      {stage0_33[441], stage0_33[442], stage0_33[443], stage0_33[444], stage0_33[445]},
      {stage0_34[310]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage1_37[46],stage1_36[90],stage1_35[125],stage1_34[126],stage1_33[179]}
   );
   gpc615_5 gpc1373 (
      {stage0_33[446], stage0_33[447], stage0_33[448], stage0_33[449], stage0_33[450]},
      {stage0_34[311]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage1_37[47],stage1_36[91],stage1_35[126],stage1_34[127],stage1_33[180]}
   );
   gpc615_5 gpc1374 (
      {stage0_33[451], stage0_33[452], stage0_33[453], stage0_33[454], stage0_33[455]},
      {stage0_34[312]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage1_37[48],stage1_36[92],stage1_35[127],stage1_34[128],stage1_33[181]}
   );
   gpc615_5 gpc1375 (
      {stage0_33[456], stage0_33[457], stage0_33[458], stage0_33[459], stage0_33[460]},
      {stage0_34[313]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage1_37[49],stage1_36[93],stage1_35[128],stage1_34[129],stage1_33[182]}
   );
   gpc615_5 gpc1376 (
      {stage0_33[461], stage0_33[462], stage0_33[463], stage0_33[464], stage0_33[465]},
      {stage0_34[314]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage1_37[50],stage1_36[94],stage1_35[129],stage1_34[130],stage1_33[183]}
   );
   gpc615_5 gpc1377 (
      {stage0_33[466], stage0_33[467], stage0_33[468], stage0_33[469], stage0_33[470]},
      {stage0_34[315]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage1_37[51],stage1_36[95],stage1_35[130],stage1_34[131],stage1_33[184]}
   );
   gpc615_5 gpc1378 (
      {stage0_33[471], stage0_33[472], stage0_33[473], stage0_33[474], stage0_33[475]},
      {stage0_34[316]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage1_37[52],stage1_36[96],stage1_35[131],stage1_34[132],stage1_33[185]}
   );
   gpc615_5 gpc1379 (
      {stage0_33[476], stage0_33[477], stage0_33[478], stage0_33[479], stage0_33[480]},
      {stage0_34[317]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage1_37[53],stage1_36[97],stage1_35[132],stage1_34[133],stage1_33[186]}
   );
   gpc615_5 gpc1380 (
      {stage0_33[481], stage0_33[482], stage0_33[483], stage0_33[484], stage0_33[485]},
      {stage0_34[318]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage1_37[54],stage1_36[98],stage1_35[133],stage1_34[134],stage1_33[187]}
   );
   gpc615_5 gpc1381 (
      {stage0_33[486], stage0_33[487], stage0_33[488], stage0_33[489], stage0_33[490]},
      {stage0_34[319]},
      {stage0_35[330], stage0_35[331], stage0_35[332], stage0_35[333], stage0_35[334], stage0_35[335]},
      {stage1_37[55],stage1_36[99],stage1_35[134],stage1_34[135],stage1_33[188]}
   );
   gpc1163_5 gpc1382 (
      {stage0_34[320], stage0_34[321], stage0_34[322]},
      {stage0_35[336], stage0_35[337], stage0_35[338], stage0_35[339], stage0_35[340], stage0_35[341]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[56],stage1_36[100],stage1_35[135],stage1_34[136]}
   );
   gpc1163_5 gpc1383 (
      {stage0_34[323], stage0_34[324], stage0_34[325]},
      {stage0_35[342], stage0_35[343], stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[57],stage1_36[101],stage1_35[136],stage1_34[137]}
   );
   gpc615_5 gpc1384 (
      {stage0_34[326], stage0_34[327], stage0_34[328], stage0_34[329], stage0_34[330]},
      {stage0_35[348]},
      {stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5], stage0_36[6], stage0_36[7]},
      {stage1_38[2],stage1_37[58],stage1_36[102],stage1_35[137],stage1_34[138]}
   );
   gpc615_5 gpc1385 (
      {stage0_34[331], stage0_34[332], stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[349]},
      {stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13]},
      {stage1_38[3],stage1_37[59],stage1_36[103],stage1_35[138],stage1_34[139]}
   );
   gpc615_5 gpc1386 (
      {stage0_34[336], stage0_34[337], stage0_34[338], stage0_34[339], stage0_34[340]},
      {stage0_35[350]},
      {stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19]},
      {stage1_38[4],stage1_37[60],stage1_36[104],stage1_35[139],stage1_34[140]}
   );
   gpc615_5 gpc1387 (
      {stage0_34[341], stage0_34[342], stage0_34[343], stage0_34[344], stage0_34[345]},
      {stage0_35[351]},
      {stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25]},
      {stage1_38[5],stage1_37[61],stage1_36[105],stage1_35[140],stage1_34[141]}
   );
   gpc615_5 gpc1388 (
      {stage0_34[346], stage0_34[347], stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[352]},
      {stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31]},
      {stage1_38[6],stage1_37[62],stage1_36[106],stage1_35[141],stage1_34[142]}
   );
   gpc615_5 gpc1389 (
      {stage0_34[351], stage0_34[352], stage0_34[353], stage0_34[354], stage0_34[355]},
      {stage0_35[353]},
      {stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37]},
      {stage1_38[7],stage1_37[63],stage1_36[107],stage1_35[142],stage1_34[143]}
   );
   gpc615_5 gpc1390 (
      {stage0_34[356], stage0_34[357], stage0_34[358], stage0_34[359], stage0_34[360]},
      {stage0_35[354]},
      {stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43]},
      {stage1_38[8],stage1_37[64],stage1_36[108],stage1_35[143],stage1_34[144]}
   );
   gpc615_5 gpc1391 (
      {stage0_34[361], stage0_34[362], stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[355]},
      {stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48], stage0_36[49]},
      {stage1_38[9],stage1_37[65],stage1_36[109],stage1_35[144],stage1_34[145]}
   );
   gpc615_5 gpc1392 (
      {stage0_34[366], stage0_34[367], stage0_34[368], stage0_34[369], stage0_34[370]},
      {stage0_35[356]},
      {stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54], stage0_36[55]},
      {stage1_38[10],stage1_37[66],stage1_36[110],stage1_35[145],stage1_34[146]}
   );
   gpc615_5 gpc1393 (
      {stage0_34[371], stage0_34[372], stage0_34[373], stage0_34[374], stage0_34[375]},
      {stage0_35[357]},
      {stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60], stage0_36[61]},
      {stage1_38[11],stage1_37[67],stage1_36[111],stage1_35[146],stage1_34[147]}
   );
   gpc615_5 gpc1394 (
      {stage0_34[376], stage0_34[377], stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[358]},
      {stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66], stage0_36[67]},
      {stage1_38[12],stage1_37[68],stage1_36[112],stage1_35[147],stage1_34[148]}
   );
   gpc615_5 gpc1395 (
      {stage0_34[381], stage0_34[382], stage0_34[383], stage0_34[384], stage0_34[385]},
      {stage0_35[359]},
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage1_38[13],stage1_37[69],stage1_36[113],stage1_35[148],stage1_34[149]}
   );
   gpc615_5 gpc1396 (
      {stage0_34[386], stage0_34[387], stage0_34[388], stage0_34[389], stage0_34[390]},
      {stage0_35[360]},
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage1_38[14],stage1_37[70],stage1_36[114],stage1_35[149],stage1_34[150]}
   );
   gpc615_5 gpc1397 (
      {stage0_34[391], stage0_34[392], stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[361]},
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage1_38[15],stage1_37[71],stage1_36[115],stage1_35[150],stage1_34[151]}
   );
   gpc606_5 gpc1398 (
      {stage0_35[362], stage0_35[363], stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367]},
      {stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5], stage0_37[6], stage0_37[7]},
      {stage1_39[0],stage1_38[16],stage1_37[72],stage1_36[116],stage1_35[151]}
   );
   gpc606_5 gpc1399 (
      {stage0_35[368], stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12], stage0_37[13]},
      {stage1_39[1],stage1_38[17],stage1_37[73],stage1_36[117],stage1_35[152]}
   );
   gpc606_5 gpc1400 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378], stage0_35[379]},
      {stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17], stage0_37[18], stage0_37[19]},
      {stage1_39[2],stage1_38[18],stage1_37[74],stage1_36[118],stage1_35[153]}
   );
   gpc606_5 gpc1401 (
      {stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383], stage0_35[384], stage0_35[385]},
      {stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23], stage0_37[24], stage0_37[25]},
      {stage1_39[3],stage1_38[19],stage1_37[75],stage1_36[119],stage1_35[154]}
   );
   gpc606_5 gpc1402 (
      {stage0_35[386], stage0_35[387], stage0_35[388], stage0_35[389], stage0_35[390], stage0_35[391]},
      {stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29], stage0_37[30], stage0_37[31]},
      {stage1_39[4],stage1_38[20],stage1_37[76],stage1_36[120],stage1_35[155]}
   );
   gpc606_5 gpc1403 (
      {stage0_35[392], stage0_35[393], stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397]},
      {stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35], stage0_37[36], stage0_37[37]},
      {stage1_39[5],stage1_38[21],stage1_37[77],stage1_36[121],stage1_35[156]}
   );
   gpc606_5 gpc1404 (
      {stage0_35[398], stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41], stage0_37[42], stage0_37[43]},
      {stage1_39[6],stage1_38[22],stage1_37[78],stage1_36[122],stage1_35[157]}
   );
   gpc606_5 gpc1405 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408], stage0_35[409]},
      {stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48], stage0_37[49]},
      {stage1_39[7],stage1_38[23],stage1_37[79],stage1_36[123],stage1_35[158]}
   );
   gpc606_5 gpc1406 (
      {stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413], stage0_35[414], stage0_35[415]},
      {stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54], stage0_37[55]},
      {stage1_39[8],stage1_38[24],stage1_37[80],stage1_36[124],stage1_35[159]}
   );
   gpc606_5 gpc1407 (
      {stage0_35[416], stage0_35[417], stage0_35[418], stage0_35[419], stage0_35[420], stage0_35[421]},
      {stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60], stage0_37[61]},
      {stage1_39[9],stage1_38[25],stage1_37[81],stage1_36[125],stage1_35[160]}
   );
   gpc606_5 gpc1408 (
      {stage0_35[422], stage0_35[423], stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427]},
      {stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66], stage0_37[67]},
      {stage1_39[10],stage1_38[26],stage1_37[82],stage1_36[126],stage1_35[161]}
   );
   gpc606_5 gpc1409 (
      {stage0_35[428], stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72], stage0_37[73]},
      {stage1_39[11],stage1_38[27],stage1_37[83],stage1_36[127],stage1_35[162]}
   );
   gpc606_5 gpc1410 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438], stage0_35[439]},
      {stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78], stage0_37[79]},
      {stage1_39[12],stage1_38[28],stage1_37[84],stage1_36[128],stage1_35[163]}
   );
   gpc606_5 gpc1411 (
      {stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443], stage0_35[444], stage0_35[445]},
      {stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84], stage0_37[85]},
      {stage1_39[13],stage1_38[29],stage1_37[85],stage1_36[129],stage1_35[164]}
   );
   gpc606_5 gpc1412 (
      {stage0_35[446], stage0_35[447], stage0_35[448], stage0_35[449], stage0_35[450], stage0_35[451]},
      {stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90], stage0_37[91]},
      {stage1_39[14],stage1_38[30],stage1_37[86],stage1_36[130],stage1_35[165]}
   );
   gpc606_5 gpc1413 (
      {stage0_35[452], stage0_35[453], stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457]},
      {stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96], stage0_37[97]},
      {stage1_39[15],stage1_38[31],stage1_37[87],stage1_36[131],stage1_35[166]}
   );
   gpc606_5 gpc1414 (
      {stage0_35[458], stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102], stage0_37[103]},
      {stage1_39[16],stage1_38[32],stage1_37[88],stage1_36[132],stage1_35[167]}
   );
   gpc606_5 gpc1415 (
      {stage0_35[464], stage0_35[465], stage0_35[466], stage0_35[467], stage0_35[468], stage0_35[469]},
      {stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108], stage0_37[109]},
      {stage1_39[17],stage1_38[33],stage1_37[89],stage1_36[133],stage1_35[168]}
   );
   gpc615_5 gpc1416 (
      {stage0_35[470], stage0_35[471], stage0_35[472], stage0_35[473], stage0_35[474]},
      {stage0_36[86]},
      {stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114], stage0_37[115]},
      {stage1_39[18],stage1_38[34],stage1_37[90],stage1_36[134],stage1_35[169]}
   );
   gpc615_5 gpc1417 (
      {stage0_35[475], stage0_35[476], stage0_35[477], stage0_35[478], stage0_35[479]},
      {stage0_36[87]},
      {stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120], stage0_37[121]},
      {stage1_39[19],stage1_38[35],stage1_37[91],stage1_36[135],stage1_35[170]}
   );
   gpc615_5 gpc1418 (
      {stage0_35[480], stage0_35[481], stage0_35[482], stage0_35[483], stage0_35[484]},
      {stage0_36[88]},
      {stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126], stage0_37[127]},
      {stage1_39[20],stage1_38[36],stage1_37[92],stage1_36[136],stage1_35[171]}
   );
   gpc615_5 gpc1419 (
      {stage0_35[485], stage0_35[486], stage0_35[487], stage0_35[488], stage0_35[489]},
      {stage0_36[89]},
      {stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132], stage0_37[133]},
      {stage1_39[21],stage1_38[37],stage1_37[93],stage1_36[137],stage1_35[172]}
   );
   gpc615_5 gpc1420 (
      {stage0_35[490], stage0_35[491], stage0_35[492], stage0_35[493], stage0_35[494]},
      {stage0_36[90]},
      {stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138], stage0_37[139]},
      {stage1_39[22],stage1_38[38],stage1_37[94],stage1_36[138],stage1_35[173]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[23],stage1_38[39],stage1_37[95],stage1_36[139]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[97], stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[24],stage1_38[40],stage1_37[96],stage1_36[140]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[25],stage1_38[41],stage1_37[97],stage1_36[141]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[109], stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[26],stage1_38[42],stage1_37[98],stage1_36[142]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[115], stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[27],stage1_38[43],stage1_37[99],stage1_36[143]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[121], stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[28],stage1_38[44],stage1_37[100],stage1_36[144]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[127], stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[29],stage1_38[45],stage1_37[101],stage1_36[145]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[133], stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[30],stage1_38[46],stage1_37[102],stage1_36[146]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[139], stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[31],stage1_38[47],stage1_37[103],stage1_36[147]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[145], stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[32],stage1_38[48],stage1_37[104],stage1_36[148]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[151], stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[33],stage1_38[49],stage1_37[105],stage1_36[149]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[157], stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[34],stage1_38[50],stage1_37[106],stage1_36[150]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[163], stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[35],stage1_38[51],stage1_37[107],stage1_36[151]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[169], stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[36],stage1_38[52],stage1_37[108],stage1_36[152]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[175], stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[37],stage1_38[53],stage1_37[109],stage1_36[153]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[181], stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[38],stage1_38[54],stage1_37[110],stage1_36[154]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[187], stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[39],stage1_38[55],stage1_37[111],stage1_36[155]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[193], stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[40],stage1_38[56],stage1_37[112],stage1_36[156]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[199], stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[41],stage1_38[57],stage1_37[113],stage1_36[157]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[205], stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[42],stage1_38[58],stage1_37[114],stage1_36[158]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[211], stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[43],stage1_38[59],stage1_37[115],stage1_36[159]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[217], stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[44],stage1_38[60],stage1_37[116],stage1_36[160]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[223], stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[45],stage1_38[61],stage1_37[117],stage1_36[161]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[229], stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[46],stage1_38[62],stage1_37[118],stage1_36[162]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[235], stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[47],stage1_38[63],stage1_37[119],stage1_36[163]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[241], stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[48],stage1_38[64],stage1_37[120],stage1_36[164]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[247], stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[49],stage1_38[65],stage1_37[121],stage1_36[165]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[253], stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[50],stage1_38[66],stage1_37[122],stage1_36[166]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[259], stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[51],stage1_38[67],stage1_37[123],stage1_36[167]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[265], stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[52],stage1_38[68],stage1_37[124],stage1_36[168]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[271], stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[53],stage1_38[69],stage1_37[125],stage1_36[169]}
   );
   gpc606_5 gpc1452 (
      {stage0_36[277], stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[54],stage1_38[70],stage1_37[126],stage1_36[170]}
   );
   gpc606_5 gpc1453 (
      {stage0_36[283], stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[55],stage1_38[71],stage1_37[127],stage1_36[171]}
   );
   gpc606_5 gpc1454 (
      {stage0_36[289], stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[56],stage1_38[72],stage1_37[128],stage1_36[172]}
   );
   gpc606_5 gpc1455 (
      {stage0_36[295], stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[57],stage1_38[73],stage1_37[129],stage1_36[173]}
   );
   gpc606_5 gpc1456 (
      {stage0_36[301], stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[58],stage1_38[74],stage1_37[130],stage1_36[174]}
   );
   gpc606_5 gpc1457 (
      {stage0_36[307], stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[59],stage1_38[75],stage1_37[131],stage1_36[175]}
   );
   gpc606_5 gpc1458 (
      {stage0_36[313], stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[60],stage1_38[76],stage1_37[132],stage1_36[176]}
   );
   gpc606_5 gpc1459 (
      {stage0_36[319], stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[61],stage1_38[77],stage1_37[133],stage1_36[177]}
   );
   gpc606_5 gpc1460 (
      {stage0_36[325], stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[62],stage1_38[78],stage1_37[134],stage1_36[178]}
   );
   gpc606_5 gpc1461 (
      {stage0_36[331], stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[63],stage1_38[79],stage1_37[135],stage1_36[179]}
   );
   gpc615_5 gpc1462 (
      {stage0_36[337], stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341]},
      {stage0_37[140]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[64],stage1_38[80],stage1_37[136],stage1_36[180]}
   );
   gpc615_5 gpc1463 (
      {stage0_36[342], stage0_36[343], stage0_36[344], stage0_36[345], stage0_36[346]},
      {stage0_37[141]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[65],stage1_38[81],stage1_37[137],stage1_36[181]}
   );
   gpc615_5 gpc1464 (
      {stage0_36[347], stage0_36[348], stage0_36[349], stage0_36[350], stage0_36[351]},
      {stage0_37[142]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[66],stage1_38[82],stage1_37[138],stage1_36[182]}
   );
   gpc615_5 gpc1465 (
      {stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355], stage0_36[356]},
      {stage0_37[143]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[67],stage1_38[83],stage1_37[139],stage1_36[183]}
   );
   gpc615_5 gpc1466 (
      {stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_37[144]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[68],stage1_38[84],stage1_37[140],stage1_36[184]}
   );
   gpc615_5 gpc1467 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366]},
      {stage0_37[145]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[69],stage1_38[85],stage1_37[141],stage1_36[185]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150], stage0_37[151]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[47],stage1_39[70],stage1_38[86],stage1_37[142]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156], stage0_37[157]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[48],stage1_39[71],stage1_38[87],stage1_37[143]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162], stage0_37[163]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[49],stage1_39[72],stage1_38[88],stage1_37[144]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168], stage0_37[169]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[50],stage1_39[73],stage1_38[89],stage1_37[145]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174], stage0_37[175]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[51],stage1_39[74],stage1_38[90],stage1_37[146]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180], stage0_37[181]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[52],stage1_39[75],stage1_38[91],stage1_37[147]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186], stage0_37[187]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[53],stage1_39[76],stage1_38[92],stage1_37[148]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192], stage0_37[193]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[54],stage1_39[77],stage1_38[93],stage1_37[149]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198], stage0_37[199]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[55],stage1_39[78],stage1_38[94],stage1_37[150]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204], stage0_37[205]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[56],stage1_39[79],stage1_38[95],stage1_37[151]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210], stage0_37[211]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[57],stage1_39[80],stage1_38[96],stage1_37[152]}
   );
   gpc606_5 gpc1479 (
      {stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216], stage0_37[217]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[58],stage1_39[81],stage1_38[97],stage1_37[153]}
   );
   gpc606_5 gpc1480 (
      {stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222], stage0_37[223]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[59],stage1_39[82],stage1_38[98],stage1_37[154]}
   );
   gpc606_5 gpc1481 (
      {stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228], stage0_37[229]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[60],stage1_39[83],stage1_38[99],stage1_37[155]}
   );
   gpc606_5 gpc1482 (
      {stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234], stage0_37[235]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[61],stage1_39[84],stage1_38[100],stage1_37[156]}
   );
   gpc606_5 gpc1483 (
      {stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240], stage0_37[241]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[62],stage1_39[85],stage1_38[101],stage1_37[157]}
   );
   gpc606_5 gpc1484 (
      {stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246], stage0_37[247]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[63],stage1_39[86],stage1_38[102],stage1_37[158]}
   );
   gpc606_5 gpc1485 (
      {stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252], stage0_37[253]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[64],stage1_39[87],stage1_38[103],stage1_37[159]}
   );
   gpc606_5 gpc1486 (
      {stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258], stage0_37[259]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[65],stage1_39[88],stage1_38[104],stage1_37[160]}
   );
   gpc606_5 gpc1487 (
      {stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264], stage0_37[265]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[66],stage1_39[89],stage1_38[105],stage1_37[161]}
   );
   gpc606_5 gpc1488 (
      {stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270], stage0_37[271]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[67],stage1_39[90],stage1_38[106],stage1_37[162]}
   );
   gpc606_5 gpc1489 (
      {stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276], stage0_37[277]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[68],stage1_39[91],stage1_38[107],stage1_37[163]}
   );
   gpc606_5 gpc1490 (
      {stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282], stage0_37[283]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[69],stage1_39[92],stage1_38[108],stage1_37[164]}
   );
   gpc606_5 gpc1491 (
      {stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288], stage0_37[289]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[70],stage1_39[93],stage1_38[109],stage1_37[165]}
   );
   gpc606_5 gpc1492 (
      {stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294], stage0_37[295]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[71],stage1_39[94],stage1_38[110],stage1_37[166]}
   );
   gpc606_5 gpc1493 (
      {stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300], stage0_37[301]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[72],stage1_39[95],stage1_38[111],stage1_37[167]}
   );
   gpc606_5 gpc1494 (
      {stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306], stage0_37[307]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[73],stage1_39[96],stage1_38[112],stage1_37[168]}
   );
   gpc606_5 gpc1495 (
      {stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312], stage0_37[313]},
      {stage0_39[162], stage0_39[163], stage0_39[164], stage0_39[165], stage0_39[166], stage0_39[167]},
      {stage1_41[27],stage1_40[74],stage1_39[97],stage1_38[113],stage1_37[169]}
   );
   gpc606_5 gpc1496 (
      {stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318], stage0_37[319]},
      {stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171], stage0_39[172], stage0_39[173]},
      {stage1_41[28],stage1_40[75],stage1_39[98],stage1_38[114],stage1_37[170]}
   );
   gpc606_5 gpc1497 (
      {stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324], stage0_37[325]},
      {stage0_39[174], stage0_39[175], stage0_39[176], stage0_39[177], stage0_39[178], stage0_39[179]},
      {stage1_41[29],stage1_40[76],stage1_39[99],stage1_38[115],stage1_37[171]}
   );
   gpc606_5 gpc1498 (
      {stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330], stage0_37[331]},
      {stage0_39[180], stage0_39[181], stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185]},
      {stage1_41[30],stage1_40[77],stage1_39[100],stage1_38[116],stage1_37[172]}
   );
   gpc606_5 gpc1499 (
      {stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336], stage0_37[337]},
      {stage0_39[186], stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage1_41[31],stage1_40[78],stage1_39[101],stage1_38[117],stage1_37[173]}
   );
   gpc606_5 gpc1500 (
      {stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342], stage0_37[343]},
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196], stage0_39[197]},
      {stage1_41[32],stage1_40[79],stage1_39[102],stage1_38[118],stage1_37[174]}
   );
   gpc606_5 gpc1501 (
      {stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348], stage0_37[349]},
      {stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201], stage0_39[202], stage0_39[203]},
      {stage1_41[33],stage1_40[80],stage1_39[103],stage1_38[119],stage1_37[175]}
   );
   gpc606_5 gpc1502 (
      {stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354], stage0_37[355]},
      {stage0_39[204], stage0_39[205], stage0_39[206], stage0_39[207], stage0_39[208], stage0_39[209]},
      {stage1_41[34],stage1_40[81],stage1_39[104],stage1_38[120],stage1_37[176]}
   );
   gpc606_5 gpc1503 (
      {stage0_37[356], stage0_37[357], stage0_37[358], stage0_37[359], stage0_37[360], stage0_37[361]},
      {stage0_39[210], stage0_39[211], stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215]},
      {stage1_41[35],stage1_40[82],stage1_39[105],stage1_38[121],stage1_37[177]}
   );
   gpc606_5 gpc1504 (
      {stage0_37[362], stage0_37[363], stage0_37[364], stage0_37[365], stage0_37[366], stage0_37[367]},
      {stage0_39[216], stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage1_41[36],stage1_40[83],stage1_39[106],stage1_38[122],stage1_37[178]}
   );
   gpc606_5 gpc1505 (
      {stage0_37[368], stage0_37[369], stage0_37[370], stage0_37[371], stage0_37[372], stage0_37[373]},
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226], stage0_39[227]},
      {stage1_41[37],stage1_40[84],stage1_39[107],stage1_38[123],stage1_37[179]}
   );
   gpc606_5 gpc1506 (
      {stage0_37[374], stage0_37[375], stage0_37[376], stage0_37[377], stage0_37[378], stage0_37[379]},
      {stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231], stage0_39[232], stage0_39[233]},
      {stage1_41[38],stage1_40[85],stage1_39[108],stage1_38[124],stage1_37[180]}
   );
   gpc606_5 gpc1507 (
      {stage0_37[380], stage0_37[381], stage0_37[382], stage0_37[383], stage0_37[384], stage0_37[385]},
      {stage0_39[234], stage0_39[235], stage0_39[236], stage0_39[237], stage0_39[238], stage0_39[239]},
      {stage1_41[39],stage1_40[86],stage1_39[109],stage1_38[125],stage1_37[181]}
   );
   gpc606_5 gpc1508 (
      {stage0_37[386], stage0_37[387], stage0_37[388], stage0_37[389], stage0_37[390], stage0_37[391]},
      {stage0_39[240], stage0_39[241], stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245]},
      {stage1_41[40],stage1_40[87],stage1_39[110],stage1_38[126],stage1_37[182]}
   );
   gpc615_5 gpc1509 (
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286]},
      {stage0_39[246]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[41],stage1_40[88],stage1_39[111],stage1_38[127]}
   );
   gpc615_5 gpc1510 (
      {stage0_38[287], stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291]},
      {stage0_39[247]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[42],stage1_40[89],stage1_39[112],stage1_38[128]}
   );
   gpc615_5 gpc1511 (
      {stage0_38[292], stage0_38[293], stage0_38[294], stage0_38[295], stage0_38[296]},
      {stage0_39[248]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[43],stage1_40[90],stage1_39[113],stage1_38[129]}
   );
   gpc615_5 gpc1512 (
      {stage0_38[297], stage0_38[298], stage0_38[299], stage0_38[300], stage0_38[301]},
      {stage0_39[249]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[44],stage1_40[91],stage1_39[114],stage1_38[130]}
   );
   gpc615_5 gpc1513 (
      {stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305], stage0_38[306]},
      {stage0_39[250]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[45],stage1_40[92],stage1_39[115],stage1_38[131]}
   );
   gpc615_5 gpc1514 (
      {stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage0_39[251]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[46],stage1_40[93],stage1_39[116],stage1_38[132]}
   );
   gpc615_5 gpc1515 (
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316]},
      {stage0_39[252]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[47],stage1_40[94],stage1_39[117],stage1_38[133]}
   );
   gpc615_5 gpc1516 (
      {stage0_38[317], stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321]},
      {stage0_39[253]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[48],stage1_40[95],stage1_39[118],stage1_38[134]}
   );
   gpc615_5 gpc1517 (
      {stage0_38[322], stage0_38[323], stage0_38[324], stage0_38[325], stage0_38[326]},
      {stage0_39[254]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[49],stage1_40[96],stage1_39[119],stage1_38[135]}
   );
   gpc615_5 gpc1518 (
      {stage0_38[327], stage0_38[328], stage0_38[329], stage0_38[330], stage0_38[331]},
      {stage0_39[255]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[50],stage1_40[97],stage1_39[120],stage1_38[136]}
   );
   gpc615_5 gpc1519 (
      {stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335], stage0_38[336]},
      {stage0_39[256]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[51],stage1_40[98],stage1_39[121],stage1_38[137]}
   );
   gpc615_5 gpc1520 (
      {stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage0_39[257]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[52],stage1_40[99],stage1_39[122],stage1_38[138]}
   );
   gpc615_5 gpc1521 (
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346]},
      {stage0_39[258]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[53],stage1_40[100],stage1_39[123],stage1_38[139]}
   );
   gpc615_5 gpc1522 (
      {stage0_38[347], stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351]},
      {stage0_39[259]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[54],stage1_40[101],stage1_39[124],stage1_38[140]}
   );
   gpc615_5 gpc1523 (
      {stage0_38[352], stage0_38[353], stage0_38[354], stage0_38[355], stage0_38[356]},
      {stage0_39[260]},
      {stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89]},
      {stage1_42[14],stage1_41[55],stage1_40[102],stage1_39[125],stage1_38[141]}
   );
   gpc615_5 gpc1524 (
      {stage0_38[357], stage0_38[358], stage0_38[359], stage0_38[360], stage0_38[361]},
      {stage0_39[261]},
      {stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95]},
      {stage1_42[15],stage1_41[56],stage1_40[103],stage1_39[126],stage1_38[142]}
   );
   gpc615_5 gpc1525 (
      {stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365], stage0_38[366]},
      {stage0_39[262]},
      {stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101]},
      {stage1_42[16],stage1_41[57],stage1_40[104],stage1_39[127],stage1_38[143]}
   );
   gpc615_5 gpc1526 (
      {stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370], stage0_38[371]},
      {stage0_39[263]},
      {stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107]},
      {stage1_42[17],stage1_41[58],stage1_40[105],stage1_39[128],stage1_38[144]}
   );
   gpc615_5 gpc1527 (
      {stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375], stage0_38[376]},
      {stage0_39[264]},
      {stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113]},
      {stage1_42[18],stage1_41[59],stage1_40[106],stage1_39[129],stage1_38[145]}
   );
   gpc615_5 gpc1528 (
      {stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380], stage0_38[381]},
      {stage0_39[265]},
      {stage0_40[114], stage0_40[115], stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119]},
      {stage1_42[19],stage1_41[60],stage1_40[107],stage1_39[130],stage1_38[146]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[266], stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270]},
      {stage0_40[120]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[20],stage1_41[61],stage1_40[108],stage1_39[131]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[271], stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275]},
      {stage0_40[121]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[21],stage1_41[62],stage1_40[109],stage1_39[132]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[276], stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280]},
      {stage0_40[122]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[22],stage1_41[63],stage1_40[110],stage1_39[133]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[281], stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285]},
      {stage0_40[123]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[23],stage1_41[64],stage1_40[111],stage1_39[134]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[286], stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290]},
      {stage0_40[124]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[24],stage1_41[65],stage1_40[112],stage1_39[135]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[291], stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295]},
      {stage0_40[125]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[25],stage1_41[66],stage1_40[113],stage1_39[136]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[296], stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300]},
      {stage0_40[126]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[26],stage1_41[67],stage1_40[114],stage1_39[137]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[301], stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305]},
      {stage0_40[127]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[27],stage1_41[68],stage1_40[115],stage1_39[138]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[306], stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310]},
      {stage0_40[128]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[28],stage1_41[69],stage1_40[116],stage1_39[139]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[311], stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315]},
      {stage0_40[129]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[29],stage1_41[70],stage1_40[117],stage1_39[140]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[316], stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320]},
      {stage0_40[130]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[30],stage1_41[71],stage1_40[118],stage1_39[141]}
   );
   gpc615_5 gpc1540 (
      {stage0_39[321], stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325]},
      {stage0_40[131]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[31],stage1_41[72],stage1_40[119],stage1_39[142]}
   );
   gpc615_5 gpc1541 (
      {stage0_39[326], stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330]},
      {stage0_40[132]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[32],stage1_41[73],stage1_40[120],stage1_39[143]}
   );
   gpc615_5 gpc1542 (
      {stage0_39[331], stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335]},
      {stage0_40[133]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[33],stage1_41[74],stage1_40[121],stage1_39[144]}
   );
   gpc615_5 gpc1543 (
      {stage0_39[336], stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340]},
      {stage0_40[134]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[34],stage1_41[75],stage1_40[122],stage1_39[145]}
   );
   gpc615_5 gpc1544 (
      {stage0_39[341], stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345]},
      {stage0_40[135]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[35],stage1_41[76],stage1_40[123],stage1_39[146]}
   );
   gpc615_5 gpc1545 (
      {stage0_39[346], stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350]},
      {stage0_40[136]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[36],stage1_41[77],stage1_40[124],stage1_39[147]}
   );
   gpc615_5 gpc1546 (
      {stage0_39[351], stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355]},
      {stage0_40[137]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[37],stage1_41[78],stage1_40[125],stage1_39[148]}
   );
   gpc615_5 gpc1547 (
      {stage0_39[356], stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360]},
      {stage0_40[138]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[38],stage1_41[79],stage1_40[126],stage1_39[149]}
   );
   gpc615_5 gpc1548 (
      {stage0_39[361], stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365]},
      {stage0_40[139]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[39],stage1_41[80],stage1_40[127],stage1_39[150]}
   );
   gpc615_5 gpc1549 (
      {stage0_39[366], stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370]},
      {stage0_40[140]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[40],stage1_41[81],stage1_40[128],stage1_39[151]}
   );
   gpc615_5 gpc1550 (
      {stage0_39[371], stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375]},
      {stage0_40[141]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[41],stage1_41[82],stage1_40[129],stage1_39[152]}
   );
   gpc615_5 gpc1551 (
      {stage0_39[376], stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380]},
      {stage0_40[142]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[42],stage1_41[83],stage1_40[130],stage1_39[153]}
   );
   gpc615_5 gpc1552 (
      {stage0_39[381], stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385]},
      {stage0_40[143]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[43],stage1_41[84],stage1_40[131],stage1_39[154]}
   );
   gpc615_5 gpc1553 (
      {stage0_39[386], stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390]},
      {stage0_40[144]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[44],stage1_41[85],stage1_40[132],stage1_39[155]}
   );
   gpc615_5 gpc1554 (
      {stage0_39[391], stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395]},
      {stage0_40[145]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[45],stage1_41[86],stage1_40[133],stage1_39[156]}
   );
   gpc615_5 gpc1555 (
      {stage0_39[396], stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400]},
      {stage0_40[146]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[46],stage1_41[87],stage1_40[134],stage1_39[157]}
   );
   gpc615_5 gpc1556 (
      {stage0_39[401], stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405]},
      {stage0_40[147]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[47],stage1_41[88],stage1_40[135],stage1_39[158]}
   );
   gpc615_5 gpc1557 (
      {stage0_39[406], stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410]},
      {stage0_40[148]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[48],stage1_41[89],stage1_40[136],stage1_39[159]}
   );
   gpc615_5 gpc1558 (
      {stage0_39[411], stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415]},
      {stage0_40[149]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[49],stage1_41[90],stage1_40[137],stage1_39[160]}
   );
   gpc615_5 gpc1559 (
      {stage0_39[416], stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420]},
      {stage0_40[150]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[50],stage1_41[91],stage1_40[138],stage1_39[161]}
   );
   gpc615_5 gpc1560 (
      {stage0_39[421], stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425]},
      {stage0_40[151]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[51],stage1_41[92],stage1_40[139],stage1_39[162]}
   );
   gpc615_5 gpc1561 (
      {stage0_39[426], stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430]},
      {stage0_40[152]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[52],stage1_41[93],stage1_40[140],stage1_39[163]}
   );
   gpc615_5 gpc1562 (
      {stage0_39[431], stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435]},
      {stage0_40[153]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[53],stage1_41[94],stage1_40[141],stage1_39[164]}
   );
   gpc615_5 gpc1563 (
      {stage0_39[436], stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440]},
      {stage0_40[154]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[54],stage1_41[95],stage1_40[142],stage1_39[165]}
   );
   gpc615_5 gpc1564 (
      {stage0_39[441], stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445]},
      {stage0_40[155]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[55],stage1_41[96],stage1_40[143],stage1_39[166]}
   );
   gpc615_5 gpc1565 (
      {stage0_39[446], stage0_39[447], stage0_39[448], stage0_39[449], stage0_39[450]},
      {stage0_40[156]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[56],stage1_41[97],stage1_40[144],stage1_39[167]}
   );
   gpc615_5 gpc1566 (
      {stage0_39[451], stage0_39[452], stage0_39[453], stage0_39[454], stage0_39[455]},
      {stage0_40[157]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[57],stage1_41[98],stage1_40[145],stage1_39[168]}
   );
   gpc615_5 gpc1567 (
      {stage0_39[456], stage0_39[457], stage0_39[458], stage0_39[459], stage0_39[460]},
      {stage0_40[158]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[58],stage1_41[99],stage1_40[146],stage1_39[169]}
   );
   gpc615_5 gpc1568 (
      {stage0_39[461], stage0_39[462], stage0_39[463], stage0_39[464], stage0_39[465]},
      {stage0_40[159]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[59],stage1_41[100],stage1_40[147],stage1_39[170]}
   );
   gpc615_5 gpc1569 (
      {stage0_39[466], stage0_39[467], stage0_39[468], stage0_39[469], stage0_39[470]},
      {stage0_40[160]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[60],stage1_41[101],stage1_40[148],stage1_39[171]}
   );
   gpc615_5 gpc1570 (
      {stage0_39[471], stage0_39[472], stage0_39[473], stage0_39[474], stage0_39[475]},
      {stage0_40[161]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[61],stage1_41[102],stage1_40[149],stage1_39[172]}
   );
   gpc615_5 gpc1571 (
      {stage0_39[476], stage0_39[477], stage0_39[478], stage0_39[479], stage0_39[480]},
      {stage0_40[162]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[62],stage1_41[103],stage1_40[150],stage1_39[173]}
   );
   gpc615_5 gpc1572 (
      {stage0_39[481], stage0_39[482], stage0_39[483], stage0_39[484], stage0_39[485]},
      {stage0_40[163]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[63],stage1_41[104],stage1_40[151],stage1_39[174]}
   );
   gpc615_5 gpc1573 (
      {stage0_39[486], stage0_39[487], stage0_39[488], stage0_39[489], stage0_39[490]},
      {stage0_40[164]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[64],stage1_41[105],stage1_40[152],stage1_39[175]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169], stage0_40[170]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[45],stage1_42[65],stage1_41[106],stage1_40[153]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175], stage0_40[176]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[46],stage1_42[66],stage1_41[107],stage1_40[154]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181], stage0_40[182]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[47],stage1_42[67],stage1_41[108],stage1_40[155]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187], stage0_40[188]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[48],stage1_42[68],stage1_41[109],stage1_40[156]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193], stage0_40[194]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[49],stage1_42[69],stage1_41[110],stage1_40[157]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199], stage0_40[200]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[50],stage1_42[70],stage1_41[111],stage1_40[158]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205], stage0_40[206]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[51],stage1_42[71],stage1_41[112],stage1_40[159]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211], stage0_40[212]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[52],stage1_42[72],stage1_41[113],stage1_40[160]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217], stage0_40[218]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[53],stage1_42[73],stage1_41[114],stage1_40[161]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223], stage0_40[224]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[54],stage1_42[74],stage1_41[115],stage1_40[162]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229], stage0_40[230]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[55],stage1_42[75],stage1_41[116],stage1_40[163]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235], stage0_40[236]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[56],stage1_42[76],stage1_41[117],stage1_40[164]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241], stage0_40[242]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[57],stage1_42[77],stage1_41[118],stage1_40[165]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247], stage0_40[248]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[58],stage1_42[78],stage1_41[119],stage1_40[166]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253], stage0_40[254]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[59],stage1_42[79],stage1_41[120],stage1_40[167]}
   );
   gpc606_5 gpc1589 (
      {stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259], stage0_40[260]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[60],stage1_42[80],stage1_41[121],stage1_40[168]}
   );
   gpc606_5 gpc1590 (
      {stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265], stage0_40[266]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[61],stage1_42[81],stage1_41[122],stage1_40[169]}
   );
   gpc606_5 gpc1591 (
      {stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271], stage0_40[272]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[62],stage1_42[82],stage1_41[123],stage1_40[170]}
   );
   gpc606_5 gpc1592 (
      {stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277], stage0_40[278]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[63],stage1_42[83],stage1_41[124],stage1_40[171]}
   );
   gpc606_5 gpc1593 (
      {stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283], stage0_40[284]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[64],stage1_42[84],stage1_41[125],stage1_40[172]}
   );
   gpc606_5 gpc1594 (
      {stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289], stage0_40[290]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[65],stage1_42[85],stage1_41[126],stage1_40[173]}
   );
   gpc606_5 gpc1595 (
      {stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295], stage0_40[296]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[66],stage1_42[86],stage1_41[127],stage1_40[174]}
   );
   gpc606_5 gpc1596 (
      {stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301], stage0_40[302]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[67],stage1_42[87],stage1_41[128],stage1_40[175]}
   );
   gpc606_5 gpc1597 (
      {stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307], stage0_40[308]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[68],stage1_42[88],stage1_41[129],stage1_40[176]}
   );
   gpc606_5 gpc1598 (
      {stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313], stage0_40[314]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[69],stage1_42[89],stage1_41[130],stage1_40[177]}
   );
   gpc606_5 gpc1599 (
      {stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319], stage0_40[320]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[70],stage1_42[90],stage1_41[131],stage1_40[178]}
   );
   gpc606_5 gpc1600 (
      {stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325], stage0_40[326]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[71],stage1_42[91],stage1_41[132],stage1_40[179]}
   );
   gpc606_5 gpc1601 (
      {stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331], stage0_40[332]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[72],stage1_42[92],stage1_41[133],stage1_40[180]}
   );
   gpc606_5 gpc1602 (
      {stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337], stage0_40[338]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[73],stage1_42[93],stage1_41[134],stage1_40[181]}
   );
   gpc606_5 gpc1603 (
      {stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343], stage0_40[344]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[74],stage1_42[94],stage1_41[135],stage1_40[182]}
   );
   gpc606_5 gpc1604 (
      {stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349], stage0_40[350]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[75],stage1_42[95],stage1_41[136],stage1_40[183]}
   );
   gpc606_5 gpc1605 (
      {stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355], stage0_40[356]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[76],stage1_42[96],stage1_41[137],stage1_40[184]}
   );
   gpc606_5 gpc1606 (
      {stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361], stage0_40[362]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[77],stage1_42[97],stage1_41[138],stage1_40[185]}
   );
   gpc606_5 gpc1607 (
      {stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367], stage0_40[368]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[78],stage1_42[98],stage1_41[139],stage1_40[186]}
   );
   gpc606_5 gpc1608 (
      {stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373], stage0_40[374]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[79],stage1_42[99],stage1_41[140],stage1_40[187]}
   );
   gpc606_5 gpc1609 (
      {stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379], stage0_40[380]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[80],stage1_42[100],stage1_41[141],stage1_40[188]}
   );
   gpc606_5 gpc1610 (
      {stage0_40[381], stage0_40[382], stage0_40[383], stage0_40[384], stage0_40[385], stage0_40[386]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[81],stage1_42[101],stage1_41[142],stage1_40[189]}
   );
   gpc606_5 gpc1611 (
      {stage0_40[387], stage0_40[388], stage0_40[389], stage0_40[390], stage0_40[391], stage0_40[392]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[82],stage1_42[102],stage1_41[143],stage1_40[190]}
   );
   gpc606_5 gpc1612 (
      {stage0_40[393], stage0_40[394], stage0_40[395], stage0_40[396], stage0_40[397], stage0_40[398]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[83],stage1_42[103],stage1_41[144],stage1_40[191]}
   );
   gpc606_5 gpc1613 (
      {stage0_40[399], stage0_40[400], stage0_40[401], stage0_40[402], stage0_40[403], stage0_40[404]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[84],stage1_42[104],stage1_41[145],stage1_40[192]}
   );
   gpc606_5 gpc1614 (
      {stage0_40[405], stage0_40[406], stage0_40[407], stage0_40[408], stage0_40[409], stage0_40[410]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[85],stage1_42[105],stage1_41[146],stage1_40[193]}
   );
   gpc606_5 gpc1615 (
      {stage0_40[411], stage0_40[412], stage0_40[413], stage0_40[414], stage0_40[415], stage0_40[416]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[86],stage1_42[106],stage1_41[147],stage1_40[194]}
   );
   gpc606_5 gpc1616 (
      {stage0_40[417], stage0_40[418], stage0_40[419], stage0_40[420], stage0_40[421], stage0_40[422]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[87],stage1_42[107],stage1_41[148],stage1_40[195]}
   );
   gpc606_5 gpc1617 (
      {stage0_40[423], stage0_40[424], stage0_40[425], stage0_40[426], stage0_40[427], stage0_40[428]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[88],stage1_42[108],stage1_41[149],stage1_40[196]}
   );
   gpc606_5 gpc1618 (
      {stage0_40[429], stage0_40[430], stage0_40[431], stage0_40[432], stage0_40[433], stage0_40[434]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[89],stage1_42[109],stage1_41[150],stage1_40[197]}
   );
   gpc606_5 gpc1619 (
      {stage0_40[435], stage0_40[436], stage0_40[437], stage0_40[438], stage0_40[439], stage0_40[440]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[90],stage1_42[110],stage1_41[151],stage1_40[198]}
   );
   gpc606_5 gpc1620 (
      {stage0_40[441], stage0_40[442], stage0_40[443], stage0_40[444], stage0_40[445], stage0_40[446]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[91],stage1_42[111],stage1_41[152],stage1_40[199]}
   );
   gpc606_5 gpc1621 (
      {stage0_40[447], stage0_40[448], stage0_40[449], stage0_40[450], stage0_40[451], stage0_40[452]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[92],stage1_42[112],stage1_41[153],stage1_40[200]}
   );
   gpc606_5 gpc1622 (
      {stage0_40[453], stage0_40[454], stage0_40[455], stage0_40[456], stage0_40[457], stage0_40[458]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[93],stage1_42[113],stage1_41[154],stage1_40[201]}
   );
   gpc606_5 gpc1623 (
      {stage0_40[459], stage0_40[460], stage0_40[461], stage0_40[462], stage0_40[463], stage0_40[464]},
      {stage0_42[294], stage0_42[295], stage0_42[296], stage0_42[297], stage0_42[298], stage0_42[299]},
      {stage1_44[49],stage1_43[94],stage1_42[114],stage1_41[155],stage1_40[202]}
   );
   gpc606_5 gpc1624 (
      {stage0_40[465], stage0_40[466], stage0_40[467], stage0_40[468], stage0_40[469], stage0_40[470]},
      {stage0_42[300], stage0_42[301], stage0_42[302], stage0_42[303], stage0_42[304], stage0_42[305]},
      {stage1_44[50],stage1_43[95],stage1_42[115],stage1_41[156],stage1_40[203]}
   );
   gpc606_5 gpc1625 (
      {stage0_40[471], stage0_40[472], stage0_40[473], stage0_40[474], stage0_40[475], stage0_40[476]},
      {stage0_42[306], stage0_42[307], stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311]},
      {stage1_44[51],stage1_43[96],stage1_42[116],stage1_41[157],stage1_40[204]}
   );
   gpc606_5 gpc1626 (
      {stage0_40[477], stage0_40[478], stage0_40[479], stage0_40[480], stage0_40[481], stage0_40[482]},
      {stage0_42[312], stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage1_44[52],stage1_43[97],stage1_42[117],stage1_41[158],stage1_40[205]}
   );
   gpc606_5 gpc1627 (
      {stage0_40[483], stage0_40[484], stage0_40[485], stage0_40[486], stage0_40[487], stage0_40[488]},
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322], stage0_42[323]},
      {stage1_44[53],stage1_43[98],stage1_42[118],stage1_41[159],stage1_40[206]}
   );
   gpc606_5 gpc1628 (
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[54],stage1_43[99],stage1_42[119],stage1_41[160]}
   );
   gpc606_5 gpc1629 (
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[55],stage1_43[100],stage1_42[120],stage1_41[161]}
   );
   gpc606_5 gpc1630 (
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[56],stage1_43[101],stage1_42[121],stage1_41[162]}
   );
   gpc606_5 gpc1631 (
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[57],stage1_43[102],stage1_42[122],stage1_41[163]}
   );
   gpc606_5 gpc1632 (
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[58],stage1_43[103],stage1_42[123],stage1_41[164]}
   );
   gpc606_5 gpc1633 (
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[59],stage1_43[104],stage1_42[124],stage1_41[165]}
   );
   gpc606_5 gpc1634 (
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[60],stage1_43[105],stage1_42[125],stage1_41[166]}
   );
   gpc606_5 gpc1635 (
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[61],stage1_43[106],stage1_42[126],stage1_41[167]}
   );
   gpc606_5 gpc1636 (
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[62],stage1_43[107],stage1_42[127],stage1_41[168]}
   );
   gpc606_5 gpc1637 (
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[63],stage1_43[108],stage1_42[128],stage1_41[169]}
   );
   gpc606_5 gpc1638 (
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[64],stage1_43[109],stage1_42[129],stage1_41[170]}
   );
   gpc606_5 gpc1639 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[65],stage1_43[110],stage1_42[130],stage1_41[171]}
   );
   gpc606_5 gpc1640 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[66],stage1_43[111],stage1_42[131],stage1_41[172]}
   );
   gpc606_5 gpc1641 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[67],stage1_43[112],stage1_42[132],stage1_41[173]}
   );
   gpc606_5 gpc1642 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[68],stage1_43[113],stage1_42[133],stage1_41[174]}
   );
   gpc606_5 gpc1643 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[69],stage1_43[114],stage1_42[134],stage1_41[175]}
   );
   gpc606_5 gpc1644 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[70],stage1_43[115],stage1_42[135],stage1_41[176]}
   );
   gpc606_5 gpc1645 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[71],stage1_43[116],stage1_42[136],stage1_41[177]}
   );
   gpc606_5 gpc1646 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[72],stage1_43[117],stage1_42[137],stage1_41[178]}
   );
   gpc606_5 gpc1647 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[73],stage1_43[118],stage1_42[138],stage1_41[179]}
   );
   gpc606_5 gpc1648 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[74],stage1_43[119],stage1_42[139],stage1_41[180]}
   );
   gpc606_5 gpc1649 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[75],stage1_43[120],stage1_42[140],stage1_41[181]}
   );
   gpc606_5 gpc1650 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[76],stage1_43[121],stage1_42[141],stage1_41[182]}
   );
   gpc606_5 gpc1651 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[77],stage1_43[122],stage1_42[142],stage1_41[183]}
   );
   gpc606_5 gpc1652 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[78],stage1_43[123],stage1_42[143],stage1_41[184]}
   );
   gpc606_5 gpc1653 (
      {stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327], stage0_42[328], stage0_42[329]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[79],stage1_43[124],stage1_42[144]}
   );
   gpc606_5 gpc1654 (
      {stage0_42[330], stage0_42[331], stage0_42[332], stage0_42[333], stage0_42[334], stage0_42[335]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[80],stage1_43[125],stage1_42[145]}
   );
   gpc606_5 gpc1655 (
      {stage0_42[336], stage0_42[337], stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[81],stage1_43[126],stage1_42[146]}
   );
   gpc606_5 gpc1656 (
      {stage0_42[342], stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[82],stage1_43[127],stage1_42[147]}
   );
   gpc606_5 gpc1657 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352], stage0_42[353]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[83],stage1_43[128],stage1_42[148]}
   );
   gpc606_5 gpc1658 (
      {stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357], stage0_42[358], stage0_42[359]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[84],stage1_43[129],stage1_42[149]}
   );
   gpc606_5 gpc1659 (
      {stage0_42[360], stage0_42[361], stage0_42[362], stage0_42[363], stage0_42[364], stage0_42[365]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[85],stage1_43[130],stage1_42[150]}
   );
   gpc615_5 gpc1660 (
      {stage0_42[366], stage0_42[367], stage0_42[368], stage0_42[369], stage0_42[370]},
      {stage0_43[150]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[86],stage1_43[131],stage1_42[151]}
   );
   gpc615_5 gpc1661 (
      {stage0_42[371], stage0_42[372], stage0_42[373], stage0_42[374], stage0_42[375]},
      {stage0_43[151]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[87],stage1_43[132],stage1_42[152]}
   );
   gpc615_5 gpc1662 (
      {stage0_42[376], stage0_42[377], stage0_42[378], stage0_42[379], stage0_42[380]},
      {stage0_43[152]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[88],stage1_43[133],stage1_42[153]}
   );
   gpc615_5 gpc1663 (
      {stage0_42[381], stage0_42[382], stage0_42[383], stage0_42[384], stage0_42[385]},
      {stage0_43[153]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[89],stage1_43[134],stage1_42[154]}
   );
   gpc615_5 gpc1664 (
      {stage0_42[386], stage0_42[387], stage0_42[388], stage0_42[389], stage0_42[390]},
      {stage0_43[154]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[90],stage1_43[135],stage1_42[155]}
   );
   gpc615_5 gpc1665 (
      {stage0_42[391], stage0_42[392], stage0_42[393], stage0_42[394], stage0_42[395]},
      {stage0_43[155]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[91],stage1_43[136],stage1_42[156]}
   );
   gpc615_5 gpc1666 (
      {stage0_42[396], stage0_42[397], stage0_42[398], stage0_42[399], stage0_42[400]},
      {stage0_43[156]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[92],stage1_43[137],stage1_42[157]}
   );
   gpc615_5 gpc1667 (
      {stage0_42[401], stage0_42[402], stage0_42[403], stage0_42[404], stage0_42[405]},
      {stage0_43[157]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[93],stage1_43[138],stage1_42[158]}
   );
   gpc615_5 gpc1668 (
      {stage0_42[406], stage0_42[407], stage0_42[408], stage0_42[409], stage0_42[410]},
      {stage0_43[158]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[94],stage1_43[139],stage1_42[159]}
   );
   gpc615_5 gpc1669 (
      {stage0_42[411], stage0_42[412], stage0_42[413], stage0_42[414], stage0_42[415]},
      {stage0_43[159]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[95],stage1_43[140],stage1_42[160]}
   );
   gpc615_5 gpc1670 (
      {stage0_42[416], stage0_42[417], stage0_42[418], stage0_42[419], stage0_42[420]},
      {stage0_43[160]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[96],stage1_43[141],stage1_42[161]}
   );
   gpc615_5 gpc1671 (
      {stage0_42[421], stage0_42[422], stage0_42[423], stage0_42[424], stage0_42[425]},
      {stage0_43[161]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[97],stage1_43[142],stage1_42[162]}
   );
   gpc615_5 gpc1672 (
      {stage0_42[426], stage0_42[427], stage0_42[428], stage0_42[429], stage0_42[430]},
      {stage0_43[162]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[98],stage1_43[143],stage1_42[163]}
   );
   gpc615_5 gpc1673 (
      {stage0_42[431], stage0_42[432], stage0_42[433], stage0_42[434], stage0_42[435]},
      {stage0_43[163]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[99],stage1_43[144],stage1_42[164]}
   );
   gpc615_5 gpc1674 (
      {stage0_42[436], stage0_42[437], stage0_42[438], stage0_42[439], stage0_42[440]},
      {stage0_43[164]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[100],stage1_43[145],stage1_42[165]}
   );
   gpc615_5 gpc1675 (
      {stage0_42[441], stage0_42[442], stage0_42[443], stage0_42[444], stage0_42[445]},
      {stage0_43[165]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[101],stage1_43[146],stage1_42[166]}
   );
   gpc615_5 gpc1676 (
      {stage0_42[446], stage0_42[447], stage0_42[448], stage0_42[449], stage0_42[450]},
      {stage0_43[166]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[102],stage1_43[147],stage1_42[167]}
   );
   gpc606_5 gpc1677 (
      {stage0_43[167], stage0_43[168], stage0_43[169], stage0_43[170], stage0_43[171], stage0_43[172]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[24],stage1_45[49],stage1_44[103],stage1_43[148]}
   );
   gpc606_5 gpc1678 (
      {stage0_43[173], stage0_43[174], stage0_43[175], stage0_43[176], stage0_43[177], stage0_43[178]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[25],stage1_45[50],stage1_44[104],stage1_43[149]}
   );
   gpc606_5 gpc1679 (
      {stage0_43[179], stage0_43[180], stage0_43[181], stage0_43[182], stage0_43[183], stage0_43[184]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[26],stage1_45[51],stage1_44[105],stage1_43[150]}
   );
   gpc606_5 gpc1680 (
      {stage0_43[185], stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[27],stage1_45[52],stage1_44[106],stage1_43[151]}
   );
   gpc606_5 gpc1681 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195], stage0_43[196]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[28],stage1_45[53],stage1_44[107],stage1_43[152]}
   );
   gpc606_5 gpc1682 (
      {stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200], stage0_43[201], stage0_43[202]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[29],stage1_45[54],stage1_44[108],stage1_43[153]}
   );
   gpc606_5 gpc1683 (
      {stage0_43[203], stage0_43[204], stage0_43[205], stage0_43[206], stage0_43[207], stage0_43[208]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[30],stage1_45[55],stage1_44[109],stage1_43[154]}
   );
   gpc606_5 gpc1684 (
      {stage0_43[209], stage0_43[210], stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[31],stage1_45[56],stage1_44[110],stage1_43[155]}
   );
   gpc606_5 gpc1685 (
      {stage0_43[215], stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[32],stage1_45[57],stage1_44[111],stage1_43[156]}
   );
   gpc606_5 gpc1686 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225], stage0_43[226]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[33],stage1_45[58],stage1_44[112],stage1_43[157]}
   );
   gpc606_5 gpc1687 (
      {stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230], stage0_43[231], stage0_43[232]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[34],stage1_45[59],stage1_44[113],stage1_43[158]}
   );
   gpc606_5 gpc1688 (
      {stage0_43[233], stage0_43[234], stage0_43[235], stage0_43[236], stage0_43[237], stage0_43[238]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[35],stage1_45[60],stage1_44[114],stage1_43[159]}
   );
   gpc606_5 gpc1689 (
      {stage0_43[239], stage0_43[240], stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[36],stage1_45[61],stage1_44[115],stage1_43[160]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[245], stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249]},
      {stage0_44[144]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[37],stage1_45[62],stage1_44[116],stage1_43[161]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[250], stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254]},
      {stage0_44[145]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[38],stage1_45[63],stage1_44[117],stage1_43[162]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[255], stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259]},
      {stage0_44[146]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[39],stage1_45[64],stage1_44[118],stage1_43[163]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[260], stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264]},
      {stage0_44[147]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[40],stage1_45[65],stage1_44[119],stage1_43[164]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[265], stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269]},
      {stage0_44[148]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[41],stage1_45[66],stage1_44[120],stage1_43[165]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[270], stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274]},
      {stage0_44[149]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[42],stage1_45[67],stage1_44[121],stage1_43[166]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[275], stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279]},
      {stage0_44[150]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[43],stage1_45[68],stage1_44[122],stage1_43[167]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[280], stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284]},
      {stage0_44[151]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[44],stage1_45[69],stage1_44[123],stage1_43[168]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[285], stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289]},
      {stage0_44[152]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[45],stage1_45[70],stage1_44[124],stage1_43[169]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[290], stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294]},
      {stage0_44[153]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[46],stage1_45[71],stage1_44[125],stage1_43[170]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[295], stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299]},
      {stage0_44[154]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[47],stage1_45[72],stage1_44[126],stage1_43[171]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[300], stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304]},
      {stage0_44[155]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[48],stage1_45[73],stage1_44[127],stage1_43[172]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[305], stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309]},
      {stage0_44[156]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[49],stage1_45[74],stage1_44[128],stage1_43[173]}
   );
   gpc615_5 gpc1703 (
      {stage0_43[310], stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314]},
      {stage0_44[157]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[50],stage1_45[75],stage1_44[129],stage1_43[174]}
   );
   gpc615_5 gpc1704 (
      {stage0_43[315], stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319]},
      {stage0_44[158]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[51],stage1_45[76],stage1_44[130],stage1_43[175]}
   );
   gpc615_5 gpc1705 (
      {stage0_43[320], stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324]},
      {stage0_44[159]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[52],stage1_45[77],stage1_44[131],stage1_43[176]}
   );
   gpc615_5 gpc1706 (
      {stage0_43[325], stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329]},
      {stage0_44[160]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[53],stage1_45[78],stage1_44[132],stage1_43[177]}
   );
   gpc615_5 gpc1707 (
      {stage0_43[330], stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334]},
      {stage0_44[161]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[54],stage1_45[79],stage1_44[133],stage1_43[178]}
   );
   gpc615_5 gpc1708 (
      {stage0_43[335], stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339]},
      {stage0_44[162]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[55],stage1_45[80],stage1_44[134],stage1_43[179]}
   );
   gpc615_5 gpc1709 (
      {stage0_43[340], stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344]},
      {stage0_44[163]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[56],stage1_45[81],stage1_44[135],stage1_43[180]}
   );
   gpc615_5 gpc1710 (
      {stage0_43[345], stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349]},
      {stage0_44[164]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[57],stage1_45[82],stage1_44[136],stage1_43[181]}
   );
   gpc615_5 gpc1711 (
      {stage0_43[350], stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354]},
      {stage0_44[165]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[58],stage1_45[83],stage1_44[137],stage1_43[182]}
   );
   gpc615_5 gpc1712 (
      {stage0_43[355], stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359]},
      {stage0_44[166]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[59],stage1_45[84],stage1_44[138],stage1_43[183]}
   );
   gpc615_5 gpc1713 (
      {stage0_43[360], stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364]},
      {stage0_44[167]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[60],stage1_45[85],stage1_44[139],stage1_43[184]}
   );
   gpc615_5 gpc1714 (
      {stage0_43[365], stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369]},
      {stage0_44[168]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[61],stage1_45[86],stage1_44[140],stage1_43[185]}
   );
   gpc615_5 gpc1715 (
      {stage0_43[370], stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374]},
      {stage0_44[169]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[62],stage1_45[87],stage1_44[141],stage1_43[186]}
   );
   gpc615_5 gpc1716 (
      {stage0_43[375], stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379]},
      {stage0_44[170]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[63],stage1_45[88],stage1_44[142],stage1_43[187]}
   );
   gpc615_5 gpc1717 (
      {stage0_43[380], stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384]},
      {stage0_44[171]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[64],stage1_45[89],stage1_44[143],stage1_43[188]}
   );
   gpc615_5 gpc1718 (
      {stage0_43[385], stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389]},
      {stage0_44[172]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[65],stage1_45[90],stage1_44[144],stage1_43[189]}
   );
   gpc615_5 gpc1719 (
      {stage0_43[390], stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394]},
      {stage0_44[173]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[66],stage1_45[91],stage1_44[145],stage1_43[190]}
   );
   gpc615_5 gpc1720 (
      {stage0_43[395], stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399]},
      {stage0_44[174]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[67],stage1_45[92],stage1_44[146],stage1_43[191]}
   );
   gpc615_5 gpc1721 (
      {stage0_43[400], stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404]},
      {stage0_44[175]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[68],stage1_45[93],stage1_44[147],stage1_43[192]}
   );
   gpc615_5 gpc1722 (
      {stage0_43[405], stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409]},
      {stage0_44[176]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[69],stage1_45[94],stage1_44[148],stage1_43[193]}
   );
   gpc615_5 gpc1723 (
      {stage0_43[410], stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414]},
      {stage0_44[177]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[70],stage1_45[95],stage1_44[149],stage1_43[194]}
   );
   gpc615_5 gpc1724 (
      {stage0_43[415], stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419]},
      {stage0_44[178]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[71],stage1_45[96],stage1_44[150],stage1_43[195]}
   );
   gpc615_5 gpc1725 (
      {stage0_43[420], stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424]},
      {stage0_44[179]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[72],stage1_45[97],stage1_44[151],stage1_43[196]}
   );
   gpc615_5 gpc1726 (
      {stage0_43[425], stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429]},
      {stage0_44[180]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[73],stage1_45[98],stage1_44[152],stage1_43[197]}
   );
   gpc615_5 gpc1727 (
      {stage0_43[430], stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434]},
      {stage0_44[181]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[74],stage1_45[99],stage1_44[153],stage1_43[198]}
   );
   gpc615_5 gpc1728 (
      {stage0_43[435], stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439]},
      {stage0_44[182]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[75],stage1_45[100],stage1_44[154],stage1_43[199]}
   );
   gpc615_5 gpc1729 (
      {stage0_43[440], stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444]},
      {stage0_44[183]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[76],stage1_45[101],stage1_44[155],stage1_43[200]}
   );
   gpc615_5 gpc1730 (
      {stage0_43[445], stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449]},
      {stage0_44[184]},
      {stage0_45[318], stage0_45[319], stage0_45[320], stage0_45[321], stage0_45[322], stage0_45[323]},
      {stage1_47[53],stage1_46[77],stage1_45[102],stage1_44[156],stage1_43[201]}
   );
   gpc615_5 gpc1731 (
      {stage0_43[450], stage0_43[451], stage0_43[452], stage0_43[453], stage0_43[454]},
      {stage0_44[185]},
      {stage0_45[324], stage0_45[325], stage0_45[326], stage0_45[327], stage0_45[328], stage0_45[329]},
      {stage1_47[54],stage1_46[78],stage1_45[103],stage1_44[157],stage1_43[202]}
   );
   gpc615_5 gpc1732 (
      {stage0_43[455], stage0_43[456], stage0_43[457], stage0_43[458], stage0_43[459]},
      {stage0_44[186]},
      {stage0_45[330], stage0_45[331], stage0_45[332], stage0_45[333], stage0_45[334], stage0_45[335]},
      {stage1_47[55],stage1_46[79],stage1_45[104],stage1_44[158],stage1_43[203]}
   );
   gpc615_5 gpc1733 (
      {stage0_43[460], stage0_43[461], stage0_43[462], stage0_43[463], stage0_43[464]},
      {stage0_44[187]},
      {stage0_45[336], stage0_45[337], stage0_45[338], stage0_45[339], stage0_45[340], stage0_45[341]},
      {stage1_47[56],stage1_46[80],stage1_45[105],stage1_44[159],stage1_43[204]}
   );
   gpc615_5 gpc1734 (
      {stage0_43[465], stage0_43[466], stage0_43[467], stage0_43[468], stage0_43[469]},
      {stage0_44[188]},
      {stage0_45[342], stage0_45[343], stage0_45[344], stage0_45[345], stage0_45[346], stage0_45[347]},
      {stage1_47[57],stage1_46[81],stage1_45[106],stage1_44[160],stage1_43[205]}
   );
   gpc615_5 gpc1735 (
      {stage0_43[470], stage0_43[471], stage0_43[472], stage0_43[473], stage0_43[474]},
      {stage0_44[189]},
      {stage0_45[348], stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353]},
      {stage1_47[58],stage1_46[82],stage1_45[107],stage1_44[161],stage1_43[206]}
   );
   gpc606_5 gpc1736 (
      {stage0_44[190], stage0_44[191], stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[59],stage1_46[83],stage1_45[108],stage1_44[162]}
   );
   gpc606_5 gpc1737 (
      {stage0_44[196], stage0_44[197], stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[60],stage1_46[84],stage1_45[109],stage1_44[163]}
   );
   gpc606_5 gpc1738 (
      {stage0_44[202], stage0_44[203], stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[61],stage1_46[85],stage1_45[110],stage1_44[164]}
   );
   gpc606_5 gpc1739 (
      {stage0_44[208], stage0_44[209], stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[62],stage1_46[86],stage1_45[111],stage1_44[165]}
   );
   gpc606_5 gpc1740 (
      {stage0_44[214], stage0_44[215], stage0_44[216], stage0_44[217], stage0_44[218], stage0_44[219]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[63],stage1_46[87],stage1_45[112],stage1_44[166]}
   );
   gpc606_5 gpc1741 (
      {stage0_44[220], stage0_44[221], stage0_44[222], stage0_44[223], stage0_44[224], stage0_44[225]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[64],stage1_46[88],stage1_45[113],stage1_44[167]}
   );
   gpc606_5 gpc1742 (
      {stage0_44[226], stage0_44[227], stage0_44[228], stage0_44[229], stage0_44[230], stage0_44[231]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[65],stage1_46[89],stage1_45[114],stage1_44[168]}
   );
   gpc606_5 gpc1743 (
      {stage0_44[232], stage0_44[233], stage0_44[234], stage0_44[235], stage0_44[236], stage0_44[237]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[66],stage1_46[90],stage1_45[115],stage1_44[169]}
   );
   gpc606_5 gpc1744 (
      {stage0_44[238], stage0_44[239], stage0_44[240], stage0_44[241], stage0_44[242], stage0_44[243]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[67],stage1_46[91],stage1_45[116],stage1_44[170]}
   );
   gpc606_5 gpc1745 (
      {stage0_44[244], stage0_44[245], stage0_44[246], stage0_44[247], stage0_44[248], stage0_44[249]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[68],stage1_46[92],stage1_45[117],stage1_44[171]}
   );
   gpc606_5 gpc1746 (
      {stage0_44[250], stage0_44[251], stage0_44[252], stage0_44[253], stage0_44[254], stage0_44[255]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[69],stage1_46[93],stage1_45[118],stage1_44[172]}
   );
   gpc606_5 gpc1747 (
      {stage0_44[256], stage0_44[257], stage0_44[258], stage0_44[259], stage0_44[260], stage0_44[261]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[70],stage1_46[94],stage1_45[119],stage1_44[173]}
   );
   gpc606_5 gpc1748 (
      {stage0_44[262], stage0_44[263], stage0_44[264], stage0_44[265], stage0_44[266], stage0_44[267]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[71],stage1_46[95],stage1_45[120],stage1_44[174]}
   );
   gpc606_5 gpc1749 (
      {stage0_44[268], stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[72],stage1_46[96],stage1_45[121],stage1_44[175]}
   );
   gpc606_5 gpc1750 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278], stage0_44[279]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[73],stage1_46[97],stage1_45[122],stage1_44[176]}
   );
   gpc606_5 gpc1751 (
      {stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283], stage0_44[284], stage0_44[285]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[74],stage1_46[98],stage1_45[123],stage1_44[177]}
   );
   gpc606_5 gpc1752 (
      {stage0_44[286], stage0_44[287], stage0_44[288], stage0_44[289], stage0_44[290], stage0_44[291]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[75],stage1_46[99],stage1_45[124],stage1_44[178]}
   );
   gpc606_5 gpc1753 (
      {stage0_44[292], stage0_44[293], stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[76],stage1_46[100],stage1_45[125],stage1_44[179]}
   );
   gpc606_5 gpc1754 (
      {stage0_44[298], stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[77],stage1_46[101],stage1_45[126],stage1_44[180]}
   );
   gpc606_5 gpc1755 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308], stage0_44[309]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[78],stage1_46[102],stage1_45[127],stage1_44[181]}
   );
   gpc606_5 gpc1756 (
      {stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313], stage0_44[314], stage0_44[315]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[79],stage1_46[103],stage1_45[128],stage1_44[182]}
   );
   gpc606_5 gpc1757 (
      {stage0_44[316], stage0_44[317], stage0_44[318], stage0_44[319], stage0_44[320], stage0_44[321]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[80],stage1_46[104],stage1_45[129],stage1_44[183]}
   );
   gpc606_5 gpc1758 (
      {stage0_44[322], stage0_44[323], stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[81],stage1_46[105],stage1_45[130],stage1_44[184]}
   );
   gpc606_5 gpc1759 (
      {stage0_44[328], stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[82],stage1_46[106],stage1_45[131],stage1_44[185]}
   );
   gpc606_5 gpc1760 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338], stage0_44[339]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[83],stage1_46[107],stage1_45[132],stage1_44[186]}
   );
   gpc606_5 gpc1761 (
      {stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343], stage0_44[344], stage0_44[345]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[84],stage1_46[108],stage1_45[133],stage1_44[187]}
   );
   gpc606_5 gpc1762 (
      {stage0_44[346], stage0_44[347], stage0_44[348], stage0_44[349], stage0_44[350], stage0_44[351]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[85],stage1_46[109],stage1_45[134],stage1_44[188]}
   );
   gpc606_5 gpc1763 (
      {stage0_44[352], stage0_44[353], stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[86],stage1_46[110],stage1_45[135],stage1_44[189]}
   );
   gpc606_5 gpc1764 (
      {stage0_44[358], stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[87],stage1_46[111],stage1_45[136],stage1_44[190]}
   );
   gpc606_5 gpc1765 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368], stage0_44[369]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[88],stage1_46[112],stage1_45[137],stage1_44[191]}
   );
   gpc606_5 gpc1766 (
      {stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373], stage0_44[374], stage0_44[375]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[89],stage1_46[113],stage1_45[138],stage1_44[192]}
   );
   gpc606_5 gpc1767 (
      {stage0_44[376], stage0_44[377], stage0_44[378], stage0_44[379], stage0_44[380], stage0_44[381]},
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190], stage0_46[191]},
      {stage1_48[31],stage1_47[90],stage1_46[114],stage1_45[139],stage1_44[193]}
   );
   gpc606_5 gpc1768 (
      {stage0_44[382], stage0_44[383], stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387]},
      {stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195], stage0_46[196], stage0_46[197]},
      {stage1_48[32],stage1_47[91],stage1_46[115],stage1_45[140],stage1_44[194]}
   );
   gpc606_5 gpc1769 (
      {stage0_44[388], stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_46[198], stage0_46[199], stage0_46[200], stage0_46[201], stage0_46[202], stage0_46[203]},
      {stage1_48[33],stage1_47[92],stage1_46[116],stage1_45[141],stage1_44[195]}
   );
   gpc606_5 gpc1770 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398], stage0_44[399]},
      {stage0_46[204], stage0_46[205], stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209]},
      {stage1_48[34],stage1_47[93],stage1_46[117],stage1_45[142],stage1_44[196]}
   );
   gpc606_5 gpc1771 (
      {stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403], stage0_44[404], stage0_44[405]},
      {stage0_46[210], stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage1_48[35],stage1_47[94],stage1_46[118],stage1_45[143],stage1_44[197]}
   );
   gpc606_5 gpc1772 (
      {stage0_44[406], stage0_44[407], stage0_44[408], stage0_44[409], stage0_44[410], stage0_44[411]},
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220], stage0_46[221]},
      {stage1_48[36],stage1_47[95],stage1_46[119],stage1_45[144],stage1_44[198]}
   );
   gpc606_5 gpc1773 (
      {stage0_44[412], stage0_44[413], stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417]},
      {stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225], stage0_46[226], stage0_46[227]},
      {stage1_48[37],stage1_47[96],stage1_46[120],stage1_45[145],stage1_44[199]}
   );
   gpc606_5 gpc1774 (
      {stage0_44[418], stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_46[228], stage0_46[229], stage0_46[230], stage0_46[231], stage0_46[232], stage0_46[233]},
      {stage1_48[38],stage1_47[97],stage1_46[121],stage1_45[146],stage1_44[200]}
   );
   gpc606_5 gpc1775 (
      {stage0_44[424], stage0_44[425], stage0_44[426], stage0_44[427], stage0_44[428], stage0_44[429]},
      {stage0_46[234], stage0_46[235], stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239]},
      {stage1_48[39],stage1_47[98],stage1_46[122],stage1_45[147],stage1_44[201]}
   );
   gpc606_5 gpc1776 (
      {stage0_44[430], stage0_44[431], stage0_44[432], stage0_44[433], stage0_44[434], stage0_44[435]},
      {stage0_46[240], stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage1_48[40],stage1_47[99],stage1_46[123],stage1_45[148],stage1_44[202]}
   );
   gpc606_5 gpc1777 (
      {stage0_44[436], stage0_44[437], stage0_44[438], stage0_44[439], stage0_44[440], stage0_44[441]},
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250], stage0_46[251]},
      {stage1_48[41],stage1_47[100],stage1_46[124],stage1_45[149],stage1_44[203]}
   );
   gpc606_5 gpc1778 (
      {stage0_44[442], stage0_44[443], stage0_44[444], stage0_44[445], stage0_44[446], stage0_44[447]},
      {stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255], stage0_46[256], stage0_46[257]},
      {stage1_48[42],stage1_47[101],stage1_46[125],stage1_45[150],stage1_44[204]}
   );
   gpc606_5 gpc1779 (
      {stage0_45[354], stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[43],stage1_47[102],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1780 (
      {stage0_45[360], stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[44],stage1_47[103],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1781 (
      {stage0_45[366], stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[45],stage1_47[104],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1782 (
      {stage0_45[372], stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[46],stage1_47[105],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1783 (
      {stage0_45[378], stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[47],stage1_47[106],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1784 (
      {stage0_45[384], stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[48],stage1_47[107],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1785 (
      {stage0_45[390], stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[49],stage1_47[108],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1786 (
      {stage0_45[396], stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[50],stage1_47[109],stage1_46[133],stage1_45[158]}
   );
   gpc606_5 gpc1787 (
      {stage0_45[402], stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[51],stage1_47[110],stage1_46[134],stage1_45[159]}
   );
   gpc606_5 gpc1788 (
      {stage0_45[408], stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[52],stage1_47[111],stage1_46[135],stage1_45[160]}
   );
   gpc606_5 gpc1789 (
      {stage0_45[414], stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[53],stage1_47[112],stage1_46[136],stage1_45[161]}
   );
   gpc606_5 gpc1790 (
      {stage0_45[420], stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[54],stage1_47[113],stage1_46[137],stage1_45[162]}
   );
   gpc606_5 gpc1791 (
      {stage0_45[426], stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[55],stage1_47[114],stage1_46[138],stage1_45[163]}
   );
   gpc606_5 gpc1792 (
      {stage0_45[432], stage0_45[433], stage0_45[434], stage0_45[435], stage0_45[436], stage0_45[437]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[56],stage1_47[115],stage1_46[139],stage1_45[164]}
   );
   gpc606_5 gpc1793 (
      {stage0_45[438], stage0_45[439], stage0_45[440], stage0_45[441], stage0_45[442], stage0_45[443]},
      {stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage1_49[14],stage1_48[57],stage1_47[116],stage1_46[140],stage1_45[165]}
   );
   gpc606_5 gpc1794 (
      {stage0_45[444], stage0_45[445], stage0_45[446], stage0_45[447], stage0_45[448], stage0_45[449]},
      {stage0_47[90], stage0_47[91], stage0_47[92], stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage1_49[15],stage1_48[58],stage1_47[117],stage1_46[141],stage1_45[166]}
   );
   gpc606_5 gpc1795 (
      {stage0_45[450], stage0_45[451], stage0_45[452], stage0_45[453], stage0_45[454], stage0_45[455]},
      {stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage1_49[16],stage1_48[59],stage1_47[118],stage1_46[142],stage1_45[167]}
   );
   gpc606_5 gpc1796 (
      {stage0_45[456], stage0_45[457], stage0_45[458], stage0_45[459], stage0_45[460], stage0_45[461]},
      {stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage1_49[17],stage1_48[60],stage1_47[119],stage1_46[143],stage1_45[168]}
   );
   gpc606_5 gpc1797 (
      {stage0_45[462], stage0_45[463], stage0_45[464], stage0_45[465], stage0_45[466], stage0_45[467]},
      {stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage1_49[18],stage1_48[61],stage1_47[120],stage1_46[144],stage1_45[169]}
   );
   gpc606_5 gpc1798 (
      {stage0_45[468], stage0_45[469], stage0_45[470], stage0_45[471], stage0_45[472], stage0_45[473]},
      {stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117], stage0_47[118], stage0_47[119]},
      {stage1_49[19],stage1_48[62],stage1_47[121],stage1_46[145],stage1_45[170]}
   );
   gpc606_5 gpc1799 (
      {stage0_45[474], stage0_45[475], stage0_45[476], stage0_45[477], stage0_45[478], stage0_45[479]},
      {stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123], stage0_47[124], stage0_47[125]},
      {stage1_49[20],stage1_48[63],stage1_47[122],stage1_46[146],stage1_45[171]}
   );
   gpc606_5 gpc1800 (
      {stage0_45[480], stage0_45[481], stage0_45[482], stage0_45[483], stage0_45[484], stage0_45[485]},
      {stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129], stage0_47[130], stage0_47[131]},
      {stage1_49[21],stage1_48[64],stage1_47[123],stage1_46[147],stage1_45[172]}
   );
   gpc606_5 gpc1801 (
      {stage0_45[486], stage0_45[487], stage0_45[488], stage0_45[489], stage0_45[490], stage0_45[491]},
      {stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135], stage0_47[136], stage0_47[137]},
      {stage1_49[22],stage1_48[65],stage1_47[124],stage1_46[148],stage1_45[173]}
   );
   gpc606_5 gpc1802 (
      {stage0_45[492], stage0_45[493], stage0_45[494], stage0_45[495], stage0_45[496], stage0_45[497]},
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142], stage0_47[143]},
      {stage1_49[23],stage1_48[66],stage1_47[125],stage1_46[149],stage1_45[174]}
   );
   gpc615_5 gpc1803 (
      {stage0_46[258], stage0_46[259], stage0_46[260], stage0_46[261], stage0_46[262]},
      {stage0_47[144]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[24],stage1_48[67],stage1_47[126],stage1_46[150]}
   );
   gpc615_5 gpc1804 (
      {stage0_46[263], stage0_46[264], stage0_46[265], stage0_46[266], stage0_46[267]},
      {stage0_47[145]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[25],stage1_48[68],stage1_47[127],stage1_46[151]}
   );
   gpc615_5 gpc1805 (
      {stage0_46[268], stage0_46[269], stage0_46[270], stage0_46[271], stage0_46[272]},
      {stage0_47[146]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[26],stage1_48[69],stage1_47[128],stage1_46[152]}
   );
   gpc615_5 gpc1806 (
      {stage0_46[273], stage0_46[274], stage0_46[275], stage0_46[276], stage0_46[277]},
      {stage0_47[147]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[27],stage1_48[70],stage1_47[129],stage1_46[153]}
   );
   gpc615_5 gpc1807 (
      {stage0_46[278], stage0_46[279], stage0_46[280], stage0_46[281], stage0_46[282]},
      {stage0_47[148]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[28],stage1_48[71],stage1_47[130],stage1_46[154]}
   );
   gpc615_5 gpc1808 (
      {stage0_46[283], stage0_46[284], stage0_46[285], stage0_46[286], stage0_46[287]},
      {stage0_47[149]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[29],stage1_48[72],stage1_47[131],stage1_46[155]}
   );
   gpc615_5 gpc1809 (
      {stage0_46[288], stage0_46[289], stage0_46[290], stage0_46[291], stage0_46[292]},
      {stage0_47[150]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[30],stage1_48[73],stage1_47[132],stage1_46[156]}
   );
   gpc615_5 gpc1810 (
      {stage0_46[293], stage0_46[294], stage0_46[295], stage0_46[296], stage0_46[297]},
      {stage0_47[151]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[31],stage1_48[74],stage1_47[133],stage1_46[157]}
   );
   gpc615_5 gpc1811 (
      {stage0_46[298], stage0_46[299], stage0_46[300], stage0_46[301], stage0_46[302]},
      {stage0_47[152]},
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage1_50[8],stage1_49[32],stage1_48[75],stage1_47[134],stage1_46[158]}
   );
   gpc615_5 gpc1812 (
      {stage0_46[303], stage0_46[304], stage0_46[305], stage0_46[306], stage0_46[307]},
      {stage0_47[153]},
      {stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58], stage0_48[59]},
      {stage1_50[9],stage1_49[33],stage1_48[76],stage1_47[135],stage1_46[159]}
   );
   gpc615_5 gpc1813 (
      {stage0_46[308], stage0_46[309], stage0_46[310], stage0_46[311], stage0_46[312]},
      {stage0_47[154]},
      {stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64], stage0_48[65]},
      {stage1_50[10],stage1_49[34],stage1_48[77],stage1_47[136],stage1_46[160]}
   );
   gpc615_5 gpc1814 (
      {stage0_46[313], stage0_46[314], stage0_46[315], stage0_46[316], stage0_46[317]},
      {stage0_47[155]},
      {stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70], stage0_48[71]},
      {stage1_50[11],stage1_49[35],stage1_48[78],stage1_47[137],stage1_46[161]}
   );
   gpc615_5 gpc1815 (
      {stage0_46[318], stage0_46[319], stage0_46[320], stage0_46[321], stage0_46[322]},
      {stage0_47[156]},
      {stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75], stage0_48[76], stage0_48[77]},
      {stage1_50[12],stage1_49[36],stage1_48[79],stage1_47[138],stage1_46[162]}
   );
   gpc615_5 gpc1816 (
      {stage0_46[323], stage0_46[324], stage0_46[325], stage0_46[326], stage0_46[327]},
      {stage0_47[157]},
      {stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81], stage0_48[82], stage0_48[83]},
      {stage1_50[13],stage1_49[37],stage1_48[80],stage1_47[139],stage1_46[163]}
   );
   gpc615_5 gpc1817 (
      {stage0_46[328], stage0_46[329], stage0_46[330], stage0_46[331], stage0_46[332]},
      {stage0_47[158]},
      {stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89]},
      {stage1_50[14],stage1_49[38],stage1_48[81],stage1_47[140],stage1_46[164]}
   );
   gpc615_5 gpc1818 (
      {stage0_46[333], stage0_46[334], stage0_46[335], stage0_46[336], stage0_46[337]},
      {stage0_47[159]},
      {stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage1_50[15],stage1_49[39],stage1_48[82],stage1_47[141],stage1_46[165]}
   );
   gpc615_5 gpc1819 (
      {stage0_46[338], stage0_46[339], stage0_46[340], stage0_46[341], stage0_46[342]},
      {stage0_47[160]},
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100], stage0_48[101]},
      {stage1_50[16],stage1_49[40],stage1_48[83],stage1_47[142],stage1_46[166]}
   );
   gpc615_5 gpc1820 (
      {stage0_46[343], stage0_46[344], stage0_46[345], stage0_46[346], stage0_46[347]},
      {stage0_47[161]},
      {stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105], stage0_48[106], stage0_48[107]},
      {stage1_50[17],stage1_49[41],stage1_48[84],stage1_47[143],stage1_46[167]}
   );
   gpc615_5 gpc1821 (
      {stage0_46[348], stage0_46[349], stage0_46[350], stage0_46[351], stage0_46[352]},
      {stage0_47[162]},
      {stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111], stage0_48[112], stage0_48[113]},
      {stage1_50[18],stage1_49[42],stage1_48[85],stage1_47[144],stage1_46[168]}
   );
   gpc615_5 gpc1822 (
      {stage0_46[353], stage0_46[354], stage0_46[355], stage0_46[356], stage0_46[357]},
      {stage0_47[163]},
      {stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119]},
      {stage1_50[19],stage1_49[43],stage1_48[86],stage1_47[145],stage1_46[169]}
   );
   gpc615_5 gpc1823 (
      {stage0_46[358], stage0_46[359], stage0_46[360], stage0_46[361], stage0_46[362]},
      {stage0_47[164]},
      {stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage1_50[20],stage1_49[44],stage1_48[87],stage1_47[146],stage1_46[170]}
   );
   gpc615_5 gpc1824 (
      {stage0_46[363], stage0_46[364], stage0_46[365], stage0_46[366], stage0_46[367]},
      {stage0_47[165]},
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130], stage0_48[131]},
      {stage1_50[21],stage1_49[45],stage1_48[88],stage1_47[147],stage1_46[171]}
   );
   gpc615_5 gpc1825 (
      {stage0_46[368], stage0_46[369], stage0_46[370], stage0_46[371], stage0_46[372]},
      {stage0_47[166]},
      {stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135], stage0_48[136], stage0_48[137]},
      {stage1_50[22],stage1_49[46],stage1_48[89],stage1_47[148],stage1_46[172]}
   );
   gpc615_5 gpc1826 (
      {stage0_46[373], stage0_46[374], stage0_46[375], stage0_46[376], stage0_46[377]},
      {stage0_47[167]},
      {stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141], stage0_48[142], stage0_48[143]},
      {stage1_50[23],stage1_49[47],stage1_48[90],stage1_47[149],stage1_46[173]}
   );
   gpc615_5 gpc1827 (
      {stage0_46[378], stage0_46[379], stage0_46[380], stage0_46[381], stage0_46[382]},
      {stage0_47[168]},
      {stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149]},
      {stage1_50[24],stage1_49[48],stage1_48[91],stage1_47[150],stage1_46[174]}
   );
   gpc615_5 gpc1828 (
      {stage0_46[383], stage0_46[384], stage0_46[385], stage0_46[386], stage0_46[387]},
      {stage0_47[169]},
      {stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage1_50[25],stage1_49[49],stage1_48[92],stage1_47[151],stage1_46[175]}
   );
   gpc606_5 gpc1829 (
      {stage0_47[170], stage0_47[171], stage0_47[172], stage0_47[173], stage0_47[174], stage0_47[175]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[26],stage1_49[50],stage1_48[93],stage1_47[152]}
   );
   gpc606_5 gpc1830 (
      {stage0_47[176], stage0_47[177], stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[27],stage1_49[51],stage1_48[94],stage1_47[153]}
   );
   gpc606_5 gpc1831 (
      {stage0_47[182], stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[28],stage1_49[52],stage1_48[95],stage1_47[154]}
   );
   gpc606_5 gpc1832 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192], stage0_47[193]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[29],stage1_49[53],stage1_48[96],stage1_47[155]}
   );
   gpc606_5 gpc1833 (
      {stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197], stage0_47[198], stage0_47[199]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[30],stage1_49[54],stage1_48[97],stage1_47[156]}
   );
   gpc606_5 gpc1834 (
      {stage0_47[200], stage0_47[201], stage0_47[202], stage0_47[203], stage0_47[204], stage0_47[205]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[31],stage1_49[55],stage1_48[98],stage1_47[157]}
   );
   gpc606_5 gpc1835 (
      {stage0_47[206], stage0_47[207], stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[32],stage1_49[56],stage1_48[99],stage1_47[158]}
   );
   gpc606_5 gpc1836 (
      {stage0_47[212], stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[33],stage1_49[57],stage1_48[100],stage1_47[159]}
   );
   gpc606_5 gpc1837 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222], stage0_47[223]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[34],stage1_49[58],stage1_48[101],stage1_47[160]}
   );
   gpc606_5 gpc1838 (
      {stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227], stage0_47[228], stage0_47[229]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[35],stage1_49[59],stage1_48[102],stage1_47[161]}
   );
   gpc606_5 gpc1839 (
      {stage0_47[230], stage0_47[231], stage0_47[232], stage0_47[233], stage0_47[234], stage0_47[235]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[36],stage1_49[60],stage1_48[103],stage1_47[162]}
   );
   gpc606_5 gpc1840 (
      {stage0_47[236], stage0_47[237], stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[37],stage1_49[61],stage1_48[104],stage1_47[163]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[242], stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246]},
      {stage0_48[156]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[38],stage1_49[62],stage1_48[105],stage1_47[164]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[247], stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251]},
      {stage0_48[157]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[39],stage1_49[63],stage1_48[106],stage1_47[165]}
   );
   gpc615_5 gpc1843 (
      {stage0_47[252], stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256]},
      {stage0_48[158]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[40],stage1_49[64],stage1_48[107],stage1_47[166]}
   );
   gpc615_5 gpc1844 (
      {stage0_47[257], stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261]},
      {stage0_48[159]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[41],stage1_49[65],stage1_48[108],stage1_47[167]}
   );
   gpc615_5 gpc1845 (
      {stage0_47[262], stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266]},
      {stage0_48[160]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[42],stage1_49[66],stage1_48[109],stage1_47[168]}
   );
   gpc615_5 gpc1846 (
      {stage0_47[267], stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271]},
      {stage0_48[161]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[43],stage1_49[67],stage1_48[110],stage1_47[169]}
   );
   gpc615_5 gpc1847 (
      {stage0_47[272], stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276]},
      {stage0_48[162]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[44],stage1_49[68],stage1_48[111],stage1_47[170]}
   );
   gpc615_5 gpc1848 (
      {stage0_47[277], stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281]},
      {stage0_48[163]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[45],stage1_49[69],stage1_48[112],stage1_47[171]}
   );
   gpc615_5 gpc1849 (
      {stage0_47[282], stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286]},
      {stage0_48[164]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[46],stage1_49[70],stage1_48[113],stage1_47[172]}
   );
   gpc615_5 gpc1850 (
      {stage0_47[287], stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291]},
      {stage0_48[165]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[47],stage1_49[71],stage1_48[114],stage1_47[173]}
   );
   gpc615_5 gpc1851 (
      {stage0_47[292], stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296]},
      {stage0_48[166]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[48],stage1_49[72],stage1_48[115],stage1_47[174]}
   );
   gpc615_5 gpc1852 (
      {stage0_47[297], stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301]},
      {stage0_48[167]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[49],stage1_49[73],stage1_48[116],stage1_47[175]}
   );
   gpc615_5 gpc1853 (
      {stage0_47[302], stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306]},
      {stage0_48[168]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[50],stage1_49[74],stage1_48[117],stage1_47[176]}
   );
   gpc615_5 gpc1854 (
      {stage0_47[307], stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311]},
      {stage0_48[169]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[51],stage1_49[75],stage1_48[118],stage1_47[177]}
   );
   gpc615_5 gpc1855 (
      {stage0_47[312], stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316]},
      {stage0_48[170]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[52],stage1_49[76],stage1_48[119],stage1_47[178]}
   );
   gpc615_5 gpc1856 (
      {stage0_47[317], stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321]},
      {stage0_48[171]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[53],stage1_49[77],stage1_48[120],stage1_47[179]}
   );
   gpc615_5 gpc1857 (
      {stage0_47[322], stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326]},
      {stage0_48[172]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[54],stage1_49[78],stage1_48[121],stage1_47[180]}
   );
   gpc615_5 gpc1858 (
      {stage0_47[327], stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331]},
      {stage0_48[173]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[55],stage1_49[79],stage1_48[122],stage1_47[181]}
   );
   gpc615_5 gpc1859 (
      {stage0_47[332], stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336]},
      {stage0_48[174]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[56],stage1_49[80],stage1_48[123],stage1_47[182]}
   );
   gpc615_5 gpc1860 (
      {stage0_47[337], stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341]},
      {stage0_48[175]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[57],stage1_49[81],stage1_48[124],stage1_47[183]}
   );
   gpc615_5 gpc1861 (
      {stage0_47[342], stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346]},
      {stage0_48[176]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[58],stage1_49[82],stage1_48[125],stage1_47[184]}
   );
   gpc615_5 gpc1862 (
      {stage0_47[347], stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351]},
      {stage0_48[177]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[59],stage1_49[83],stage1_48[126],stage1_47[185]}
   );
   gpc615_5 gpc1863 (
      {stage0_47[352], stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356]},
      {stage0_48[178]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[60],stage1_49[84],stage1_48[127],stage1_47[186]}
   );
   gpc615_5 gpc1864 (
      {stage0_47[357], stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361]},
      {stage0_48[179]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[61],stage1_49[85],stage1_48[128],stage1_47[187]}
   );
   gpc615_5 gpc1865 (
      {stage0_47[362], stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366]},
      {stage0_48[180]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[62],stage1_49[86],stage1_48[129],stage1_47[188]}
   );
   gpc615_5 gpc1866 (
      {stage0_47[367], stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371]},
      {stage0_48[181]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[63],stage1_49[87],stage1_48[130],stage1_47[189]}
   );
   gpc615_5 gpc1867 (
      {stage0_47[372], stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376]},
      {stage0_48[182]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[64],stage1_49[88],stage1_48[131],stage1_47[190]}
   );
   gpc615_5 gpc1868 (
      {stage0_47[377], stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381]},
      {stage0_48[183]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[65],stage1_49[89],stage1_48[132],stage1_47[191]}
   );
   gpc615_5 gpc1869 (
      {stage0_47[382], stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386]},
      {stage0_48[184]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[66],stage1_49[90],stage1_48[133],stage1_47[192]}
   );
   gpc615_5 gpc1870 (
      {stage0_47[387], stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391]},
      {stage0_48[185]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[67],stage1_49[91],stage1_48[134],stage1_47[193]}
   );
   gpc615_5 gpc1871 (
      {stage0_47[392], stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396]},
      {stage0_48[186]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[68],stage1_49[92],stage1_48[135],stage1_47[194]}
   );
   gpc615_5 gpc1872 (
      {stage0_47[397], stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401]},
      {stage0_48[187]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[69],stage1_49[93],stage1_48[136],stage1_47[195]}
   );
   gpc615_5 gpc1873 (
      {stage0_47[402], stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406]},
      {stage0_48[188]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[70],stage1_49[94],stage1_48[137],stage1_47[196]}
   );
   gpc615_5 gpc1874 (
      {stage0_47[407], stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411]},
      {stage0_48[189]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[71],stage1_49[95],stage1_48[138],stage1_47[197]}
   );
   gpc615_5 gpc1875 (
      {stage0_47[412], stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416]},
      {stage0_48[190]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[72],stage1_49[96],stage1_48[139],stage1_47[198]}
   );
   gpc615_5 gpc1876 (
      {stage0_47[417], stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421]},
      {stage0_48[191]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[73],stage1_49[97],stage1_48[140],stage1_47[199]}
   );
   gpc615_5 gpc1877 (
      {stage0_47[422], stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426]},
      {stage0_48[192]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[74],stage1_49[98],stage1_48[141],stage1_47[200]}
   );
   gpc615_5 gpc1878 (
      {stage0_47[427], stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431]},
      {stage0_48[193]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[75],stage1_49[99],stage1_48[142],stage1_47[201]}
   );
   gpc615_5 gpc1879 (
      {stage0_47[432], stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436]},
      {stage0_48[194]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[76],stage1_49[100],stage1_48[143],stage1_47[202]}
   );
   gpc606_5 gpc1880 (
      {stage0_48[195], stage0_48[196], stage0_48[197], stage0_48[198], stage0_48[199], stage0_48[200]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[51],stage1_50[77],stage1_49[101],stage1_48[144]}
   );
   gpc606_5 gpc1881 (
      {stage0_48[201], stage0_48[202], stage0_48[203], stage0_48[204], stage0_48[205], stage0_48[206]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[52],stage1_50[78],stage1_49[102],stage1_48[145]}
   );
   gpc606_5 gpc1882 (
      {stage0_48[207], stage0_48[208], stage0_48[209], stage0_48[210], stage0_48[211], stage0_48[212]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[53],stage1_50[79],stage1_49[103],stage1_48[146]}
   );
   gpc606_5 gpc1883 (
      {stage0_48[213], stage0_48[214], stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[54],stage1_50[80],stage1_49[104],stage1_48[147]}
   );
   gpc606_5 gpc1884 (
      {stage0_48[219], stage0_48[220], stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[55],stage1_50[81],stage1_49[105],stage1_48[148]}
   );
   gpc606_5 gpc1885 (
      {stage0_48[225], stage0_48[226], stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[56],stage1_50[82],stage1_49[106],stage1_48[149]}
   );
   gpc606_5 gpc1886 (
      {stage0_48[231], stage0_48[232], stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[57],stage1_50[83],stage1_49[107],stage1_48[150]}
   );
   gpc606_5 gpc1887 (
      {stage0_48[237], stage0_48[238], stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[58],stage1_50[84],stage1_49[108],stage1_48[151]}
   );
   gpc606_5 gpc1888 (
      {stage0_48[243], stage0_48[244], stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[59],stage1_50[85],stage1_49[109],stage1_48[152]}
   );
   gpc606_5 gpc1889 (
      {stage0_48[249], stage0_48[250], stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[60],stage1_50[86],stage1_49[110],stage1_48[153]}
   );
   gpc606_5 gpc1890 (
      {stage0_48[255], stage0_48[256], stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[61],stage1_50[87],stage1_49[111],stage1_48[154]}
   );
   gpc606_5 gpc1891 (
      {stage0_48[261], stage0_48[262], stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[62],stage1_50[88],stage1_49[112],stage1_48[155]}
   );
   gpc606_5 gpc1892 (
      {stage0_48[267], stage0_48[268], stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[63],stage1_50[89],stage1_49[113],stage1_48[156]}
   );
   gpc606_5 gpc1893 (
      {stage0_48[273], stage0_48[274], stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[64],stage1_50[90],stage1_49[114],stage1_48[157]}
   );
   gpc606_5 gpc1894 (
      {stage0_48[279], stage0_48[280], stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[65],stage1_50[91],stage1_49[115],stage1_48[158]}
   );
   gpc606_5 gpc1895 (
      {stage0_48[285], stage0_48[286], stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[66],stage1_50[92],stage1_49[116],stage1_48[159]}
   );
   gpc606_5 gpc1896 (
      {stage0_48[291], stage0_48[292], stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[67],stage1_50[93],stage1_49[117],stage1_48[160]}
   );
   gpc606_5 gpc1897 (
      {stage0_48[297], stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[68],stage1_50[94],stage1_49[118],stage1_48[161]}
   );
   gpc606_5 gpc1898 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307], stage0_48[308]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[69],stage1_50[95],stage1_49[119],stage1_48[162]}
   );
   gpc606_5 gpc1899 (
      {stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312], stage0_48[313], stage0_48[314]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[70],stage1_50[96],stage1_49[120],stage1_48[163]}
   );
   gpc606_5 gpc1900 (
      {stage0_48[315], stage0_48[316], stage0_48[317], stage0_48[318], stage0_48[319], stage0_48[320]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[71],stage1_50[97],stage1_49[121],stage1_48[164]}
   );
   gpc606_5 gpc1901 (
      {stage0_48[321], stage0_48[322], stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[72],stage1_50[98],stage1_49[122],stage1_48[165]}
   );
   gpc606_5 gpc1902 (
      {stage0_48[327], stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[73],stage1_50[99],stage1_49[123],stage1_48[166]}
   );
   gpc606_5 gpc1903 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337], stage0_48[338]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[74],stage1_50[100],stage1_49[124],stage1_48[167]}
   );
   gpc606_5 gpc1904 (
      {stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342], stage0_48[343], stage0_48[344]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[75],stage1_50[101],stage1_49[125],stage1_48[168]}
   );
   gpc606_5 gpc1905 (
      {stage0_48[345], stage0_48[346], stage0_48[347], stage0_48[348], stage0_48[349], stage0_48[350]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[76],stage1_50[102],stage1_49[126],stage1_48[169]}
   );
   gpc606_5 gpc1906 (
      {stage0_48[351], stage0_48[352], stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[77],stage1_50[103],stage1_49[127],stage1_48[170]}
   );
   gpc606_5 gpc1907 (
      {stage0_48[357], stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[78],stage1_50[104],stage1_49[128],stage1_48[171]}
   );
   gpc606_5 gpc1908 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367], stage0_48[368]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[79],stage1_50[105],stage1_49[129],stage1_48[172]}
   );
   gpc606_5 gpc1909 (
      {stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372], stage0_48[373], stage0_48[374]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[80],stage1_50[106],stage1_49[130],stage1_48[173]}
   );
   gpc606_5 gpc1910 (
      {stage0_48[375], stage0_48[376], stage0_48[377], stage0_48[378], stage0_48[379], stage0_48[380]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[81],stage1_50[107],stage1_49[131],stage1_48[174]}
   );
   gpc606_5 gpc1911 (
      {stage0_48[381], stage0_48[382], stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[82],stage1_50[108],stage1_49[132],stage1_48[175]}
   );
   gpc606_5 gpc1912 (
      {stage0_48[387], stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[83],stage1_50[109],stage1_49[133],stage1_48[176]}
   );
   gpc606_5 gpc1913 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397], stage0_48[398]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[84],stage1_50[110],stage1_49[134],stage1_48[177]}
   );
   gpc606_5 gpc1914 (
      {stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402], stage0_48[403], stage0_48[404]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[85],stage1_50[111],stage1_49[135],stage1_48[178]}
   );
   gpc606_5 gpc1915 (
      {stage0_48[405], stage0_48[406], stage0_48[407], stage0_48[408], stage0_48[409], stage0_48[410]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[86],stage1_50[112],stage1_49[136],stage1_48[179]}
   );
   gpc606_5 gpc1916 (
      {stage0_48[411], stage0_48[412], stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[87],stage1_50[113],stage1_49[137],stage1_48[180]}
   );
   gpc606_5 gpc1917 (
      {stage0_48[417], stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[88],stage1_50[114],stage1_49[138],stage1_48[181]}
   );
   gpc606_5 gpc1918 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427], stage0_48[428]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[89],stage1_50[115],stage1_49[139],stage1_48[182]}
   );
   gpc606_5 gpc1919 (
      {stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432], stage0_48[433], stage0_48[434]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[90],stage1_50[116],stage1_49[140],stage1_48[183]}
   );
   gpc606_5 gpc1920 (
      {stage0_48[435], stage0_48[436], stage0_48[437], stage0_48[438], stage0_48[439], stage0_48[440]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[91],stage1_50[117],stage1_49[141],stage1_48[184]}
   );
   gpc606_5 gpc1921 (
      {stage0_48[441], stage0_48[442], stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[92],stage1_50[118],stage1_49[142],stage1_48[185]}
   );
   gpc606_5 gpc1922 (
      {stage0_48[447], stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[93],stage1_50[119],stage1_49[143],stage1_48[186]}
   );
   gpc606_5 gpc1923 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457], stage0_48[458]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[94],stage1_50[120],stage1_49[144],stage1_48[187]}
   );
   gpc606_5 gpc1924 (
      {stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462], stage0_48[463], stage0_48[464]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[95],stage1_50[121],stage1_49[145],stage1_48[188]}
   );
   gpc606_5 gpc1925 (
      {stage0_48[465], stage0_48[466], stage0_48[467], stage0_48[468], stage0_48[469], stage0_48[470]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[96],stage1_50[122],stage1_49[146],stage1_48[189]}
   );
   gpc606_5 gpc1926 (
      {stage0_48[471], stage0_48[472], stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[97],stage1_50[123],stage1_49[147],stage1_48[190]}
   );
   gpc606_5 gpc1927 (
      {stage0_48[477], stage0_48[478], stage0_48[479], stage0_48[480], stage0_48[481], stage0_48[482]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[98],stage1_50[124],stage1_49[148],stage1_48[191]}
   );
   gpc606_5 gpc1928 (
      {stage0_48[483], stage0_48[484], stage0_48[485], stage0_48[486], stage0_48[487], stage0_48[488]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[99],stage1_50[125],stage1_49[149],stage1_48[192]}
   );
   gpc606_5 gpc1929 (
      {stage0_48[489], stage0_48[490], stage0_48[491], stage0_48[492], stage0_48[493], stage0_48[494]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[100],stage1_50[126],stage1_49[150],stage1_48[193]}
   );
   gpc606_5 gpc1930 (
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[101],stage1_50[127],stage1_49[151]}
   );
   gpc606_5 gpc1931 (
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[102],stage1_50[128],stage1_49[152]}
   );
   gpc606_5 gpc1932 (
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[103],stage1_50[129],stage1_49[153]}
   );
   gpc606_5 gpc1933 (
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[104],stage1_50[130],stage1_49[154]}
   );
   gpc606_5 gpc1934 (
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[105],stage1_50[131],stage1_49[155]}
   );
   gpc606_5 gpc1935 (
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[106],stage1_50[132],stage1_49[156]}
   );
   gpc606_5 gpc1936 (
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[107],stage1_50[133],stage1_49[157]}
   );
   gpc606_5 gpc1937 (
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[108],stage1_50[134],stage1_49[158]}
   );
   gpc606_5 gpc1938 (
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[109],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1939 (
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[110],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1940 (
      {stage0_49[366], stage0_49[367], stage0_49[368], stage0_49[369], stage0_49[370], stage0_49[371]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[111],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1941 (
      {stage0_49[372], stage0_49[373], stage0_49[374], stage0_49[375], stage0_49[376], stage0_49[377]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[112],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1942 (
      {stage0_49[378], stage0_49[379], stage0_49[380], stage0_49[381], stage0_49[382], stage0_49[383]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[113],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1943 (
      {stage0_49[384], stage0_49[385], stage0_49[386], stage0_49[387], stage0_49[388], stage0_49[389]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[114],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1944 (
      {stage0_49[390], stage0_49[391], stage0_49[392], stage0_49[393], stage0_49[394], stage0_49[395]},
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage1_53[14],stage1_52[64],stage1_51[115],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1945 (
      {stage0_49[396], stage0_49[397], stage0_49[398], stage0_49[399], stage0_49[400], stage0_49[401]},
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage1_53[15],stage1_52[65],stage1_51[116],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1946 (
      {stage0_49[402], stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407]},
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage1_53[16],stage1_52[66],stage1_51[117],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1947 (
      {stage0_49[408], stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413]},
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage1_53[17],stage1_52[67],stage1_51[118],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1948 (
      {stage0_49[414], stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419]},
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage1_53[18],stage1_52[68],stage1_51[119],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1949 (
      {stage0_49[420], stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425]},
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage1_53[19],stage1_52[69],stage1_51[120],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1950 (
      {stage0_49[426], stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431]},
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage1_53[20],stage1_52[70],stage1_51[121],stage1_50[147],stage1_49[171]}
   );
   gpc606_5 gpc1951 (
      {stage0_49[432], stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437]},
      {stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129], stage0_51[130], stage0_51[131]},
      {stage1_53[21],stage1_52[71],stage1_51[122],stage1_50[148],stage1_49[172]}
   );
   gpc606_5 gpc1952 (
      {stage0_49[438], stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443]},
      {stage0_51[132], stage0_51[133], stage0_51[134], stage0_51[135], stage0_51[136], stage0_51[137]},
      {stage1_53[22],stage1_52[72],stage1_51[123],stage1_50[149],stage1_49[173]}
   );
   gpc606_5 gpc1953 (
      {stage0_50[300], stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[23],stage1_52[73],stage1_51[124],stage1_50[150]}
   );
   gpc606_5 gpc1954 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310], stage0_50[311]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[24],stage1_52[74],stage1_51[125],stage1_50[151]}
   );
   gpc606_5 gpc1955 (
      {stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315], stage0_50[316], stage0_50[317]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[25],stage1_52[75],stage1_51[126],stage1_50[152]}
   );
   gpc606_5 gpc1956 (
      {stage0_50[318], stage0_50[319], stage0_50[320], stage0_50[321], stage0_50[322], stage0_50[323]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[26],stage1_52[76],stage1_51[127],stage1_50[153]}
   );
   gpc606_5 gpc1957 (
      {stage0_50[324], stage0_50[325], stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[27],stage1_52[77],stage1_51[128],stage1_50[154]}
   );
   gpc606_5 gpc1958 (
      {stage0_50[330], stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[28],stage1_52[78],stage1_51[129],stage1_50[155]}
   );
   gpc606_5 gpc1959 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340], stage0_50[341]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[29],stage1_52[79],stage1_51[130],stage1_50[156]}
   );
   gpc606_5 gpc1960 (
      {stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345], stage0_50[346], stage0_50[347]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[30],stage1_52[80],stage1_51[131],stage1_50[157]}
   );
   gpc606_5 gpc1961 (
      {stage0_50[348], stage0_50[349], stage0_50[350], stage0_50[351], stage0_50[352], stage0_50[353]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[31],stage1_52[81],stage1_51[132],stage1_50[158]}
   );
   gpc606_5 gpc1962 (
      {stage0_50[354], stage0_50[355], stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[32],stage1_52[82],stage1_51[133],stage1_50[159]}
   );
   gpc606_5 gpc1963 (
      {stage0_50[360], stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[33],stage1_52[83],stage1_51[134],stage1_50[160]}
   );
   gpc606_5 gpc1964 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370], stage0_50[371]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[34],stage1_52[84],stage1_51[135],stage1_50[161]}
   );
   gpc606_5 gpc1965 (
      {stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375], stage0_50[376], stage0_50[377]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[35],stage1_52[85],stage1_51[136],stage1_50[162]}
   );
   gpc606_5 gpc1966 (
      {stage0_50[378], stage0_50[379], stage0_50[380], stage0_50[381], stage0_50[382], stage0_50[383]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[36],stage1_52[86],stage1_51[137],stage1_50[163]}
   );
   gpc606_5 gpc1967 (
      {stage0_50[384], stage0_50[385], stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[37],stage1_52[87],stage1_51[138],stage1_50[164]}
   );
   gpc606_5 gpc1968 (
      {stage0_50[390], stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[38],stage1_52[88],stage1_51[139],stage1_50[165]}
   );
   gpc606_5 gpc1969 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400], stage0_50[401]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[39],stage1_52[89],stage1_51[140],stage1_50[166]}
   );
   gpc606_5 gpc1970 (
      {stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405], stage0_50[406], stage0_50[407]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[40],stage1_52[90],stage1_51[141],stage1_50[167]}
   );
   gpc606_5 gpc1971 (
      {stage0_50[408], stage0_50[409], stage0_50[410], stage0_50[411], stage0_50[412], stage0_50[413]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[41],stage1_52[91],stage1_51[142],stage1_50[168]}
   );
   gpc606_5 gpc1972 (
      {stage0_50[414], stage0_50[415], stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[42],stage1_52[92],stage1_51[143],stage1_50[169]}
   );
   gpc606_5 gpc1973 (
      {stage0_50[420], stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[43],stage1_52[93],stage1_51[144],stage1_50[170]}
   );
   gpc606_5 gpc1974 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430], stage0_50[431]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[44],stage1_52[94],stage1_51[145],stage1_50[171]}
   );
   gpc606_5 gpc1975 (
      {stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435], stage0_50[436], stage0_50[437]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[45],stage1_52[95],stage1_51[146],stage1_50[172]}
   );
   gpc606_5 gpc1976 (
      {stage0_50[438], stage0_50[439], stage0_50[440], stage0_50[441], stage0_50[442], stage0_50[443]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[46],stage1_52[96],stage1_51[147],stage1_50[173]}
   );
   gpc606_5 gpc1977 (
      {stage0_50[444], stage0_50[445], stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[47],stage1_52[97],stage1_51[148],stage1_50[174]}
   );
   gpc606_5 gpc1978 (
      {stage0_50[450], stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[48],stage1_52[98],stage1_51[149],stage1_50[175]}
   );
   gpc606_5 gpc1979 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460], stage0_50[461]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[49],stage1_52[99],stage1_51[150],stage1_50[176]}
   );
   gpc606_5 gpc1980 (
      {stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465], stage0_50[466], stage0_50[467]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[50],stage1_52[100],stage1_51[151],stage1_50[177]}
   );
   gpc606_5 gpc1981 (
      {stage0_50[468], stage0_50[469], stage0_50[470], stage0_50[471], stage0_50[472], stage0_50[473]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[51],stage1_52[101],stage1_51[152],stage1_50[178]}
   );
   gpc606_5 gpc1982 (
      {stage0_51[138], stage0_51[139], stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[29],stage1_53[52],stage1_52[102],stage1_51[153]}
   );
   gpc606_5 gpc1983 (
      {stage0_51[144], stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[30],stage1_53[53],stage1_52[103],stage1_51[154]}
   );
   gpc606_5 gpc1984 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154], stage0_51[155]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[31],stage1_53[54],stage1_52[104],stage1_51[155]}
   );
   gpc606_5 gpc1985 (
      {stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159], stage0_51[160], stage0_51[161]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[32],stage1_53[55],stage1_52[105],stage1_51[156]}
   );
   gpc606_5 gpc1986 (
      {stage0_51[162], stage0_51[163], stage0_51[164], stage0_51[165], stage0_51[166], stage0_51[167]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[33],stage1_53[56],stage1_52[106],stage1_51[157]}
   );
   gpc606_5 gpc1987 (
      {stage0_51[168], stage0_51[169], stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[34],stage1_53[57],stage1_52[107],stage1_51[158]}
   );
   gpc606_5 gpc1988 (
      {stage0_51[174], stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[35],stage1_53[58],stage1_52[108],stage1_51[159]}
   );
   gpc606_5 gpc1989 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184], stage0_51[185]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[36],stage1_53[59],stage1_52[109],stage1_51[160]}
   );
   gpc606_5 gpc1990 (
      {stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189], stage0_51[190], stage0_51[191]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[37],stage1_53[60],stage1_52[110],stage1_51[161]}
   );
   gpc606_5 gpc1991 (
      {stage0_51[192], stage0_51[193], stage0_51[194], stage0_51[195], stage0_51[196], stage0_51[197]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[38],stage1_53[61],stage1_52[111],stage1_51[162]}
   );
   gpc606_5 gpc1992 (
      {stage0_51[198], stage0_51[199], stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[39],stage1_53[62],stage1_52[112],stage1_51[163]}
   );
   gpc606_5 gpc1993 (
      {stage0_51[204], stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[40],stage1_53[63],stage1_52[113],stage1_51[164]}
   );
   gpc606_5 gpc1994 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214], stage0_51[215]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[41],stage1_53[64],stage1_52[114],stage1_51[165]}
   );
   gpc606_5 gpc1995 (
      {stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219], stage0_51[220], stage0_51[221]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[42],stage1_53[65],stage1_52[115],stage1_51[166]}
   );
   gpc606_5 gpc1996 (
      {stage0_51[222], stage0_51[223], stage0_51[224], stage0_51[225], stage0_51[226], stage0_51[227]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[43],stage1_53[66],stage1_52[116],stage1_51[167]}
   );
   gpc606_5 gpc1997 (
      {stage0_51[228], stage0_51[229], stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[44],stage1_53[67],stage1_52[117],stage1_51[168]}
   );
   gpc606_5 gpc1998 (
      {stage0_51[234], stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[45],stage1_53[68],stage1_52[118],stage1_51[169]}
   );
   gpc606_5 gpc1999 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244], stage0_51[245]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[46],stage1_53[69],stage1_52[119],stage1_51[170]}
   );
   gpc606_5 gpc2000 (
      {stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249], stage0_51[250], stage0_51[251]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[47],stage1_53[70],stage1_52[120],stage1_51[171]}
   );
   gpc606_5 gpc2001 (
      {stage0_51[252], stage0_51[253], stage0_51[254], stage0_51[255], stage0_51[256], stage0_51[257]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[48],stage1_53[71],stage1_52[121],stage1_51[172]}
   );
   gpc606_5 gpc2002 (
      {stage0_51[258], stage0_51[259], stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[49],stage1_53[72],stage1_52[122],stage1_51[173]}
   );
   gpc606_5 gpc2003 (
      {stage0_51[264], stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[50],stage1_53[73],stage1_52[123],stage1_51[174]}
   );
   gpc606_5 gpc2004 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274], stage0_51[275]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[51],stage1_53[74],stage1_52[124],stage1_51[175]}
   );
   gpc606_5 gpc2005 (
      {stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279], stage0_51[280], stage0_51[281]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[52],stage1_53[75],stage1_52[125],stage1_51[176]}
   );
   gpc606_5 gpc2006 (
      {stage0_51[282], stage0_51[283], stage0_51[284], stage0_51[285], stage0_51[286], stage0_51[287]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[53],stage1_53[76],stage1_52[126],stage1_51[177]}
   );
   gpc606_5 gpc2007 (
      {stage0_51[288], stage0_51[289], stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[54],stage1_53[77],stage1_52[127],stage1_51[178]}
   );
   gpc606_5 gpc2008 (
      {stage0_51[294], stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[55],stage1_53[78],stage1_52[128],stage1_51[179]}
   );
   gpc606_5 gpc2009 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304], stage0_51[305]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[56],stage1_53[79],stage1_52[129],stage1_51[180]}
   );
   gpc606_5 gpc2010 (
      {stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309], stage0_51[310], stage0_51[311]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[57],stage1_53[80],stage1_52[130],stage1_51[181]}
   );
   gpc606_5 gpc2011 (
      {stage0_51[312], stage0_51[313], stage0_51[314], stage0_51[315], stage0_51[316], stage0_51[317]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[58],stage1_53[81],stage1_52[131],stage1_51[182]}
   );
   gpc606_5 gpc2012 (
      {stage0_51[318], stage0_51[319], stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[59],stage1_53[82],stage1_52[132],stage1_51[183]}
   );
   gpc606_5 gpc2013 (
      {stage0_51[324], stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[60],stage1_53[83],stage1_52[133],stage1_51[184]}
   );
   gpc606_5 gpc2014 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334], stage0_51[335]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[61],stage1_53[84],stage1_52[134],stage1_51[185]}
   );
   gpc606_5 gpc2015 (
      {stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339], stage0_51[340], stage0_51[341]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[62],stage1_53[85],stage1_52[135],stage1_51[186]}
   );
   gpc606_5 gpc2016 (
      {stage0_51[342], stage0_51[343], stage0_51[344], stage0_51[345], stage0_51[346], stage0_51[347]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[63],stage1_53[86],stage1_52[136],stage1_51[187]}
   );
   gpc606_5 gpc2017 (
      {stage0_51[348], stage0_51[349], stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[64],stage1_53[87],stage1_52[137],stage1_51[188]}
   );
   gpc606_5 gpc2018 (
      {stage0_51[354], stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[65],stage1_53[88],stage1_52[138],stage1_51[189]}
   );
   gpc606_5 gpc2019 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364], stage0_51[365]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[66],stage1_53[89],stage1_52[139],stage1_51[190]}
   );
   gpc606_5 gpc2020 (
      {stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369], stage0_51[370], stage0_51[371]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[67],stage1_53[90],stage1_52[140],stage1_51[191]}
   );
   gpc606_5 gpc2021 (
      {stage0_51[372], stage0_51[373], stage0_51[374], stage0_51[375], stage0_51[376], stage0_51[377]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[68],stage1_53[91],stage1_52[141],stage1_51[192]}
   );
   gpc606_5 gpc2022 (
      {stage0_51[378], stage0_51[379], stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[69],stage1_53[92],stage1_52[142],stage1_51[193]}
   );
   gpc606_5 gpc2023 (
      {stage0_51[384], stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[70],stage1_53[93],stage1_52[143],stage1_51[194]}
   );
   gpc606_5 gpc2024 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394], stage0_51[395]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[71],stage1_53[94],stage1_52[144],stage1_51[195]}
   );
   gpc606_5 gpc2025 (
      {stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399], stage0_51[400], stage0_51[401]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[72],stage1_53[95],stage1_52[145],stage1_51[196]}
   );
   gpc606_5 gpc2026 (
      {stage0_51[402], stage0_51[403], stage0_51[404], stage0_51[405], stage0_51[406], stage0_51[407]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[73],stage1_53[96],stage1_52[146],stage1_51[197]}
   );
   gpc606_5 gpc2027 (
      {stage0_51[408], stage0_51[409], stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[74],stage1_53[97],stage1_52[147],stage1_51[198]}
   );
   gpc606_5 gpc2028 (
      {stage0_51[414], stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[75],stage1_53[98],stage1_52[148],stage1_51[199]}
   );
   gpc606_5 gpc2029 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424], stage0_51[425]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[76],stage1_53[99],stage1_52[149],stage1_51[200]}
   );
   gpc606_5 gpc2030 (
      {stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429], stage0_51[430], stage0_51[431]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[77],stage1_53[100],stage1_52[150],stage1_51[201]}
   );
   gpc606_5 gpc2031 (
      {stage0_51[432], stage0_51[433], stage0_51[434], stage0_51[435], stage0_51[436], stage0_51[437]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[78],stage1_53[101],stage1_52[151],stage1_51[202]}
   );
   gpc615_5 gpc2032 (
      {stage0_51[438], stage0_51[439], stage0_51[440], stage0_51[441], stage0_51[442]},
      {stage0_52[174]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[79],stage1_53[102],stage1_52[152],stage1_51[203]}
   );
   gpc615_5 gpc2033 (
      {stage0_51[443], stage0_51[444], stage0_51[445], stage0_51[446], stage0_51[447]},
      {stage0_52[175]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[80],stage1_53[103],stage1_52[153],stage1_51[204]}
   );
   gpc615_5 gpc2034 (
      {stage0_51[448], stage0_51[449], stage0_51[450], stage0_51[451], stage0_51[452]},
      {stage0_52[176]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[81],stage1_53[104],stage1_52[154],stage1_51[205]}
   );
   gpc615_5 gpc2035 (
      {stage0_51[453], stage0_51[454], stage0_51[455], stage0_51[456], stage0_51[457]},
      {stage0_52[177]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[82],stage1_53[105],stage1_52[155],stage1_51[206]}
   );
   gpc615_5 gpc2036 (
      {stage0_51[458], stage0_51[459], stage0_51[460], stage0_51[461], stage0_51[462]},
      {stage0_52[178]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[83],stage1_53[106],stage1_52[156],stage1_51[207]}
   );
   gpc615_5 gpc2037 (
      {stage0_51[463], stage0_51[464], stage0_51[465], stage0_51[466], stage0_51[467]},
      {stage0_52[179]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[84],stage1_53[107],stage1_52[157],stage1_51[208]}
   );
   gpc615_5 gpc2038 (
      {stage0_51[468], stage0_51[469], stage0_51[470], stage0_51[471], stage0_51[472]},
      {stage0_52[180]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[85],stage1_53[108],stage1_52[158],stage1_51[209]}
   );
   gpc615_5 gpc2039 (
      {stage0_51[473], stage0_51[474], stage0_51[475], stage0_51[476], stage0_51[477]},
      {stage0_52[181]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[86],stage1_53[109],stage1_52[159],stage1_51[210]}
   );
   gpc615_5 gpc2040 (
      {stage0_51[478], stage0_51[479], stage0_51[480], stage0_51[481], stage0_51[482]},
      {stage0_52[182]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[87],stage1_53[110],stage1_52[160],stage1_51[211]}
   );
   gpc615_5 gpc2041 (
      {stage0_51[483], stage0_51[484], stage0_51[485], stage0_51[486], stage0_51[487]},
      {stage0_52[183]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[88],stage1_53[111],stage1_52[161],stage1_51[212]}
   );
   gpc615_5 gpc2042 (
      {stage0_51[488], stage0_51[489], stage0_51[490], stage0_51[491], stage0_51[492]},
      {stage0_52[184]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[89],stage1_53[112],stage1_52[162],stage1_51[213]}
   );
   gpc615_5 gpc2043 (
      {stage0_51[493], stage0_51[494], stage0_51[495], stage0_51[496], stage0_51[497]},
      {stage0_52[185]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[90],stage1_53[113],stage1_52[163],stage1_51[214]}
   );
   gpc623_5 gpc2044 (
      {stage0_51[498], stage0_51[499], stage0_51[500]},
      {stage0_52[186], stage0_52[187]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[91],stage1_53[114],stage1_52[164],stage1_51[215]}
   );
   gpc606_5 gpc2045 (
      {stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191], stage0_52[192], stage0_52[193]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[92],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2046 (
      {stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197], stage0_52[198], stage0_52[199]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[93],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2047 (
      {stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203], stage0_52[204], stage0_52[205]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[94],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2048 (
      {stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209], stage0_52[210], stage0_52[211]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[95],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2049 (
      {stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215], stage0_52[216], stage0_52[217]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[96],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2050 (
      {stage0_52[218], stage0_52[219], stage0_52[220], stage0_52[221], stage0_52[222], stage0_52[223]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[97],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2051 (
      {stage0_52[224], stage0_52[225], stage0_52[226], stage0_52[227], stage0_52[228], stage0_52[229]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[98],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2052 (
      {stage0_52[230], stage0_52[231], stage0_52[232], stage0_52[233], stage0_52[234], stage0_52[235]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[99],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2053 (
      {stage0_52[236], stage0_52[237], stage0_52[238], stage0_52[239], stage0_52[240], stage0_52[241]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[100],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2054 (
      {stage0_52[242], stage0_52[243], stage0_52[244], stage0_52[245], stage0_52[246], stage0_52[247]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[101],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2055 (
      {stage0_52[248], stage0_52[249], stage0_52[250], stage0_52[251], stage0_52[252], stage0_52[253]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[102],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2056 (
      {stage0_52[254], stage0_52[255], stage0_52[256], stage0_52[257], stage0_52[258], stage0_52[259]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[103],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2057 (
      {stage0_52[260], stage0_52[261], stage0_52[262], stage0_52[263], stage0_52[264], stage0_52[265]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[104],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2058 (
      {stage0_52[266], stage0_52[267], stage0_52[268], stage0_52[269], stage0_52[270], stage0_52[271]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[105],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2059 (
      {stage0_52[272], stage0_52[273], stage0_52[274], stage0_52[275], stage0_52[276], stage0_52[277]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[106],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2060 (
      {stage0_52[278], stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[107],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2061 (
      {stage0_52[284], stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[108],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2062 (
      {stage0_52[290], stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[109],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2063 (
      {stage0_52[296], stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[110],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2064 (
      {stage0_52[302], stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[111],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2065 (
      {stage0_52[308], stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[112],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2066 (
      {stage0_52[314], stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[113],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2067 (
      {stage0_52[320], stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[114],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2068 (
      {stage0_52[326], stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[115],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2069 (
      {stage0_52[332], stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[116],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2070 (
      {stage0_52[338], stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[117],stage1_53[140],stage1_52[190]}
   );
   gpc606_5 gpc2071 (
      {stage0_52[344], stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[118],stage1_53[141],stage1_52[191]}
   );
   gpc606_5 gpc2072 (
      {stage0_52[350], stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[119],stage1_53[142],stage1_52[192]}
   );
   gpc606_5 gpc2073 (
      {stage0_52[356], stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[120],stage1_53[143],stage1_52[193]}
   );
   gpc606_5 gpc2074 (
      {stage0_52[362], stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[121],stage1_53[144],stage1_52[194]}
   );
   gpc606_5 gpc2075 (
      {stage0_52[368], stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[122],stage1_53[145],stage1_52[195]}
   );
   gpc606_5 gpc2076 (
      {stage0_52[374], stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[123],stage1_53[146],stage1_52[196]}
   );
   gpc606_5 gpc2077 (
      {stage0_52[380], stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[124],stage1_53[147],stage1_52[197]}
   );
   gpc606_5 gpc2078 (
      {stage0_52[386], stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[125],stage1_53[148],stage1_52[198]}
   );
   gpc606_5 gpc2079 (
      {stage0_52[392], stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[126],stage1_53[149],stage1_52[199]}
   );
   gpc606_5 gpc2080 (
      {stage0_52[398], stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[127],stage1_53[150],stage1_52[200]}
   );
   gpc606_5 gpc2081 (
      {stage0_52[404], stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409]},
      {stage0_54[216], stage0_54[217], stage0_54[218], stage0_54[219], stage0_54[220], stage0_54[221]},
      {stage1_56[36],stage1_55[99],stage1_54[128],stage1_53[151],stage1_52[201]}
   );
   gpc606_5 gpc2082 (
      {stage0_53[378], stage0_53[379], stage0_53[380], stage0_53[381], stage0_53[382], stage0_53[383]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[37],stage1_55[100],stage1_54[129],stage1_53[152]}
   );
   gpc606_5 gpc2083 (
      {stage0_53[384], stage0_53[385], stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[38],stage1_55[101],stage1_54[130],stage1_53[153]}
   );
   gpc606_5 gpc2084 (
      {stage0_53[390], stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[39],stage1_55[102],stage1_54[131],stage1_53[154]}
   );
   gpc606_5 gpc2085 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400], stage0_53[401]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[40],stage1_55[103],stage1_54[132],stage1_53[155]}
   );
   gpc606_5 gpc2086 (
      {stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405], stage0_53[406], stage0_53[407]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[41],stage1_55[104],stage1_54[133],stage1_53[156]}
   );
   gpc606_5 gpc2087 (
      {stage0_53[408], stage0_53[409], stage0_53[410], stage0_53[411], stage0_53[412], stage0_53[413]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[42],stage1_55[105],stage1_54[134],stage1_53[157]}
   );
   gpc606_5 gpc2088 (
      {stage0_53[414], stage0_53[415], stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[43],stage1_55[106],stage1_54[135],stage1_53[158]}
   );
   gpc606_5 gpc2089 (
      {stage0_53[420], stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[44],stage1_55[107],stage1_54[136],stage1_53[159]}
   );
   gpc606_5 gpc2090 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430], stage0_53[431]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[45],stage1_55[108],stage1_54[137],stage1_53[160]}
   );
   gpc606_5 gpc2091 (
      {stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435], stage0_53[436], stage0_53[437]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[46],stage1_55[109],stage1_54[138],stage1_53[161]}
   );
   gpc606_5 gpc2092 (
      {stage0_53[438], stage0_53[439], stage0_53[440], stage0_53[441], stage0_53[442], stage0_53[443]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[47],stage1_55[110],stage1_54[139],stage1_53[162]}
   );
   gpc606_5 gpc2093 (
      {stage0_53[444], stage0_53[445], stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[48],stage1_55[111],stage1_54[140],stage1_53[163]}
   );
   gpc606_5 gpc2094 (
      {stage0_53[450], stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[49],stage1_55[112],stage1_54[141],stage1_53[164]}
   );
   gpc606_5 gpc2095 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460], stage0_53[461]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[50],stage1_55[113],stage1_54[142],stage1_53[165]}
   );
   gpc606_5 gpc2096 (
      {stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465], stage0_53[466], stage0_53[467]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[51],stage1_55[114],stage1_54[143],stage1_53[166]}
   );
   gpc606_5 gpc2097 (
      {stage0_53[468], stage0_53[469], stage0_53[470], stage0_53[471], stage0_53[472], stage0_53[473]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[52],stage1_55[115],stage1_54[144],stage1_53[167]}
   );
   gpc606_5 gpc2098 (
      {stage0_53[474], stage0_53[475], stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[53],stage1_55[116],stage1_54[145],stage1_53[168]}
   );
   gpc606_5 gpc2099 (
      {stage0_53[480], stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[54],stage1_55[117],stage1_54[146],stage1_53[169]}
   );
   gpc606_5 gpc2100 (
      {stage0_53[486], stage0_53[487], stage0_53[488], stage0_53[489], stage0_53[490], stage0_53[491]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[55],stage1_55[118],stage1_54[147],stage1_53[170]}
   );
   gpc615_5 gpc2101 (
      {stage0_53[492], stage0_53[493], stage0_53[494], stage0_53[495], stage0_53[496]},
      {stage0_54[222]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[56],stage1_55[119],stage1_54[148],stage1_53[171]}
   );
   gpc606_5 gpc2102 (
      {stage0_54[223], stage0_54[224], stage0_54[225], stage0_54[226], stage0_54[227], stage0_54[228]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[20],stage1_56[57],stage1_55[120],stage1_54[149]}
   );
   gpc606_5 gpc2103 (
      {stage0_54[229], stage0_54[230], stage0_54[231], stage0_54[232], stage0_54[233], stage0_54[234]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[21],stage1_56[58],stage1_55[121],stage1_54[150]}
   );
   gpc606_5 gpc2104 (
      {stage0_54[235], stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[22],stage1_56[59],stage1_55[122],stage1_54[151]}
   );
   gpc615_5 gpc2105 (
      {stage0_54[241], stage0_54[242], stage0_54[243], stage0_54[244], stage0_54[245]},
      {stage0_55[120]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[23],stage1_56[60],stage1_55[123],stage1_54[152]}
   );
   gpc615_5 gpc2106 (
      {stage0_54[246], stage0_54[247], stage0_54[248], stage0_54[249], stage0_54[250]},
      {stage0_55[121]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[24],stage1_56[61],stage1_55[124],stage1_54[153]}
   );
   gpc615_5 gpc2107 (
      {stage0_54[251], stage0_54[252], stage0_54[253], stage0_54[254], stage0_54[255]},
      {stage0_55[122]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[25],stage1_56[62],stage1_55[125],stage1_54[154]}
   );
   gpc615_5 gpc2108 (
      {stage0_54[256], stage0_54[257], stage0_54[258], stage0_54[259], stage0_54[260]},
      {stage0_55[123]},
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage1_58[6],stage1_57[26],stage1_56[63],stage1_55[126],stage1_54[155]}
   );
   gpc615_5 gpc2109 (
      {stage0_54[261], stage0_54[262], stage0_54[263], stage0_54[264], stage0_54[265]},
      {stage0_55[124]},
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage1_58[7],stage1_57[27],stage1_56[64],stage1_55[127],stage1_54[156]}
   );
   gpc615_5 gpc2110 (
      {stage0_54[266], stage0_54[267], stage0_54[268], stage0_54[269], stage0_54[270]},
      {stage0_55[125]},
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage1_58[8],stage1_57[28],stage1_56[65],stage1_55[128],stage1_54[157]}
   );
   gpc615_5 gpc2111 (
      {stage0_54[271], stage0_54[272], stage0_54[273], stage0_54[274], stage0_54[275]},
      {stage0_55[126]},
      {stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59]},
      {stage1_58[9],stage1_57[29],stage1_56[66],stage1_55[129],stage1_54[158]}
   );
   gpc615_5 gpc2112 (
      {stage0_54[276], stage0_54[277], stage0_54[278], stage0_54[279], stage0_54[280]},
      {stage0_55[127]},
      {stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65]},
      {stage1_58[10],stage1_57[30],stage1_56[67],stage1_55[130],stage1_54[159]}
   );
   gpc615_5 gpc2113 (
      {stage0_54[281], stage0_54[282], stage0_54[283], stage0_54[284], stage0_54[285]},
      {stage0_55[128]},
      {stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71]},
      {stage1_58[11],stage1_57[31],stage1_56[68],stage1_55[131],stage1_54[160]}
   );
   gpc615_5 gpc2114 (
      {stage0_54[286], stage0_54[287], stage0_54[288], stage0_54[289], stage0_54[290]},
      {stage0_55[129]},
      {stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77]},
      {stage1_58[12],stage1_57[32],stage1_56[69],stage1_55[132],stage1_54[161]}
   );
   gpc615_5 gpc2115 (
      {stage0_54[291], stage0_54[292], stage0_54[293], stage0_54[294], stage0_54[295]},
      {stage0_55[130]},
      {stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83]},
      {stage1_58[13],stage1_57[33],stage1_56[70],stage1_55[133],stage1_54[162]}
   );
   gpc615_5 gpc2116 (
      {stage0_54[296], stage0_54[297], stage0_54[298], stage0_54[299], stage0_54[300]},
      {stage0_55[131]},
      {stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89]},
      {stage1_58[14],stage1_57[34],stage1_56[71],stage1_55[134],stage1_54[163]}
   );
   gpc615_5 gpc2117 (
      {stage0_54[301], stage0_54[302], stage0_54[303], stage0_54[304], stage0_54[305]},
      {stage0_55[132]},
      {stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95]},
      {stage1_58[15],stage1_57[35],stage1_56[72],stage1_55[135],stage1_54[164]}
   );
   gpc615_5 gpc2118 (
      {stage0_54[306], stage0_54[307], stage0_54[308], stage0_54[309], stage0_54[310]},
      {stage0_55[133]},
      {stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101]},
      {stage1_58[16],stage1_57[36],stage1_56[73],stage1_55[136],stage1_54[165]}
   );
   gpc615_5 gpc2119 (
      {stage0_54[311], stage0_54[312], stage0_54[313], stage0_54[314], stage0_54[315]},
      {stage0_55[134]},
      {stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107]},
      {stage1_58[17],stage1_57[37],stage1_56[74],stage1_55[137],stage1_54[166]}
   );
   gpc615_5 gpc2120 (
      {stage0_54[316], stage0_54[317], stage0_54[318], stage0_54[319], stage0_54[320]},
      {stage0_55[135]},
      {stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113]},
      {stage1_58[18],stage1_57[38],stage1_56[75],stage1_55[138],stage1_54[167]}
   );
   gpc615_5 gpc2121 (
      {stage0_54[321], stage0_54[322], stage0_54[323], stage0_54[324], stage0_54[325]},
      {stage0_55[136]},
      {stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119]},
      {stage1_58[19],stage1_57[39],stage1_56[76],stage1_55[139],stage1_54[168]}
   );
   gpc615_5 gpc2122 (
      {stage0_54[326], stage0_54[327], stage0_54[328], stage0_54[329], stage0_54[330]},
      {stage0_55[137]},
      {stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125]},
      {stage1_58[20],stage1_57[40],stage1_56[77],stage1_55[140],stage1_54[169]}
   );
   gpc615_5 gpc2123 (
      {stage0_54[331], stage0_54[332], stage0_54[333], stage0_54[334], stage0_54[335]},
      {stage0_55[138]},
      {stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131]},
      {stage1_58[21],stage1_57[41],stage1_56[78],stage1_55[141],stage1_54[170]}
   );
   gpc615_5 gpc2124 (
      {stage0_54[336], stage0_54[337], stage0_54[338], stage0_54[339], stage0_54[340]},
      {stage0_55[139]},
      {stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137]},
      {stage1_58[22],stage1_57[42],stage1_56[79],stage1_55[142],stage1_54[171]}
   );
   gpc615_5 gpc2125 (
      {stage0_54[341], stage0_54[342], stage0_54[343], stage0_54[344], stage0_54[345]},
      {stage0_55[140]},
      {stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143]},
      {stage1_58[23],stage1_57[43],stage1_56[80],stage1_55[143],stage1_54[172]}
   );
   gpc615_5 gpc2126 (
      {stage0_54[346], stage0_54[347], stage0_54[348], stage0_54[349], stage0_54[350]},
      {stage0_55[141]},
      {stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149]},
      {stage1_58[24],stage1_57[44],stage1_56[81],stage1_55[144],stage1_54[173]}
   );
   gpc615_5 gpc2127 (
      {stage0_54[351], stage0_54[352], stage0_54[353], stage0_54[354], stage0_54[355]},
      {stage0_55[142]},
      {stage0_56[150], stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155]},
      {stage1_58[25],stage1_57[45],stage1_56[82],stage1_55[145],stage1_54[174]}
   );
   gpc615_5 gpc2128 (
      {stage0_54[356], stage0_54[357], stage0_54[358], stage0_54[359], stage0_54[360]},
      {stage0_55[143]},
      {stage0_56[156], stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161]},
      {stage1_58[26],stage1_57[46],stage1_56[83],stage1_55[146],stage1_54[175]}
   );
   gpc615_5 gpc2129 (
      {stage0_54[361], stage0_54[362], stage0_54[363], stage0_54[364], stage0_54[365]},
      {stage0_55[144]},
      {stage0_56[162], stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167]},
      {stage1_58[27],stage1_57[47],stage1_56[84],stage1_55[147],stage1_54[176]}
   );
   gpc615_5 gpc2130 (
      {stage0_54[366], stage0_54[367], stage0_54[368], stage0_54[369], stage0_54[370]},
      {stage0_55[145]},
      {stage0_56[168], stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173]},
      {stage1_58[28],stage1_57[48],stage1_56[85],stage1_55[148],stage1_54[177]}
   );
   gpc615_5 gpc2131 (
      {stage0_54[371], stage0_54[372], stage0_54[373], stage0_54[374], stage0_54[375]},
      {stage0_55[146]},
      {stage0_56[174], stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179]},
      {stage1_58[29],stage1_57[49],stage1_56[86],stage1_55[149],stage1_54[178]}
   );
   gpc615_5 gpc2132 (
      {stage0_54[376], stage0_54[377], stage0_54[378], stage0_54[379], stage0_54[380]},
      {stage0_55[147]},
      {stage0_56[180], stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185]},
      {stage1_58[30],stage1_57[50],stage1_56[87],stage1_55[150],stage1_54[179]}
   );
   gpc615_5 gpc2133 (
      {stage0_54[381], stage0_54[382], stage0_54[383], stage0_54[384], stage0_54[385]},
      {stage0_55[148]},
      {stage0_56[186], stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191]},
      {stage1_58[31],stage1_57[51],stage1_56[88],stage1_55[151],stage1_54[180]}
   );
   gpc615_5 gpc2134 (
      {stage0_54[386], stage0_54[387], stage0_54[388], stage0_54[389], stage0_54[390]},
      {stage0_55[149]},
      {stage0_56[192], stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197]},
      {stage1_58[32],stage1_57[52],stage1_56[89],stage1_55[152],stage1_54[181]}
   );
   gpc615_5 gpc2135 (
      {stage0_54[391], stage0_54[392], stage0_54[393], stage0_54[394], stage0_54[395]},
      {stage0_55[150]},
      {stage0_56[198], stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203]},
      {stage1_58[33],stage1_57[53],stage1_56[90],stage1_55[153],stage1_54[182]}
   );
   gpc615_5 gpc2136 (
      {stage0_54[396], stage0_54[397], stage0_54[398], stage0_54[399], stage0_54[400]},
      {stage0_55[151]},
      {stage0_56[204], stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209]},
      {stage1_58[34],stage1_57[54],stage1_56[91],stage1_55[154],stage1_54[183]}
   );
   gpc615_5 gpc2137 (
      {stage0_54[401], stage0_54[402], stage0_54[403], stage0_54[404], stage0_54[405]},
      {stage0_55[152]},
      {stage0_56[210], stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215]},
      {stage1_58[35],stage1_57[55],stage1_56[92],stage1_55[155],stage1_54[184]}
   );
   gpc615_5 gpc2138 (
      {stage0_54[406], stage0_54[407], stage0_54[408], stage0_54[409], stage0_54[410]},
      {stage0_55[153]},
      {stage0_56[216], stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221]},
      {stage1_58[36],stage1_57[56],stage1_56[93],stage1_55[156],stage1_54[185]}
   );
   gpc615_5 gpc2139 (
      {stage0_54[411], stage0_54[412], stage0_54[413], stage0_54[414], stage0_54[415]},
      {stage0_55[154]},
      {stage0_56[222], stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227]},
      {stage1_58[37],stage1_57[57],stage1_56[94],stage1_55[157],stage1_54[186]}
   );
   gpc615_5 gpc2140 (
      {stage0_54[416], stage0_54[417], stage0_54[418], stage0_54[419], stage0_54[420]},
      {stage0_55[155]},
      {stage0_56[228], stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233]},
      {stage1_58[38],stage1_57[58],stage1_56[95],stage1_55[158],stage1_54[187]}
   );
   gpc615_5 gpc2141 (
      {stage0_54[421], stage0_54[422], stage0_54[423], stage0_54[424], stage0_54[425]},
      {stage0_55[156]},
      {stage0_56[234], stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239]},
      {stage1_58[39],stage1_57[59],stage1_56[96],stage1_55[159],stage1_54[188]}
   );
   gpc615_5 gpc2142 (
      {stage0_54[426], stage0_54[427], stage0_54[428], stage0_54[429], stage0_54[430]},
      {stage0_55[157]},
      {stage0_56[240], stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245]},
      {stage1_58[40],stage1_57[60],stage1_56[97],stage1_55[160],stage1_54[189]}
   );
   gpc615_5 gpc2143 (
      {stage0_54[431], stage0_54[432], stage0_54[433], stage0_54[434], stage0_54[435]},
      {stage0_55[158]},
      {stage0_56[246], stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251]},
      {stage1_58[41],stage1_57[61],stage1_56[98],stage1_55[161],stage1_54[190]}
   );
   gpc615_5 gpc2144 (
      {stage0_54[436], stage0_54[437], stage0_54[438], stage0_54[439], stage0_54[440]},
      {stage0_55[159]},
      {stage0_56[252], stage0_56[253], stage0_56[254], stage0_56[255], stage0_56[256], stage0_56[257]},
      {stage1_58[42],stage1_57[62],stage1_56[99],stage1_55[162],stage1_54[191]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[160], stage0_55[161], stage0_55[162], stage0_55[163], stage0_55[164], stage0_55[165]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[43],stage1_57[63],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[166], stage0_55[167], stage0_55[168], stage0_55[169], stage0_55[170], stage0_55[171]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[44],stage1_57[64],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2147 (
      {stage0_55[172], stage0_55[173], stage0_55[174], stage0_55[175], stage0_55[176], stage0_55[177]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[45],stage1_57[65],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2148 (
      {stage0_55[178], stage0_55[179], stage0_55[180], stage0_55[181], stage0_55[182], stage0_55[183]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[46],stage1_57[66],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2149 (
      {stage0_55[184], stage0_55[185], stage0_55[186], stage0_55[187], stage0_55[188], stage0_55[189]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[47],stage1_57[67],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2150 (
      {stage0_55[190], stage0_55[191], stage0_55[192], stage0_55[193], stage0_55[194], stage0_55[195]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[48],stage1_57[68],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2151 (
      {stage0_55[196], stage0_55[197], stage0_55[198], stage0_55[199], stage0_55[200], stage0_55[201]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[49],stage1_57[69],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2152 (
      {stage0_55[202], stage0_55[203], stage0_55[204], stage0_55[205], stage0_55[206], stage0_55[207]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[50],stage1_57[70],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2153 (
      {stage0_55[208], stage0_55[209], stage0_55[210], stage0_55[211], stage0_55[212], stage0_55[213]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[51],stage1_57[71],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2154 (
      {stage0_55[214], stage0_55[215], stage0_55[216], stage0_55[217], stage0_55[218], stage0_55[219]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[52],stage1_57[72],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2155 (
      {stage0_55[220], stage0_55[221], stage0_55[222], stage0_55[223], stage0_55[224], stage0_55[225]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[53],stage1_57[73],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2156 (
      {stage0_55[226], stage0_55[227], stage0_55[228], stage0_55[229], stage0_55[230], stage0_55[231]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[54],stage1_57[74],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2157 (
      {stage0_55[232], stage0_55[233], stage0_55[234], stage0_55[235], stage0_55[236], stage0_55[237]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[55],stage1_57[75],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2158 (
      {stage0_55[238], stage0_55[239], stage0_55[240], stage0_55[241], stage0_55[242], stage0_55[243]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[56],stage1_57[76],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2159 (
      {stage0_55[244], stage0_55[245], stage0_55[246], stage0_55[247], stage0_55[248], stage0_55[249]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[57],stage1_57[77],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2160 (
      {stage0_55[250], stage0_55[251], stage0_55[252], stage0_55[253], stage0_55[254], stage0_55[255]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[58],stage1_57[78],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2161 (
      {stage0_55[256], stage0_55[257], stage0_55[258], stage0_55[259], stage0_55[260], stage0_55[261]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[59],stage1_57[79],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2162 (
      {stage0_55[262], stage0_55[263], stage0_55[264], stage0_55[265], stage0_55[266], stage0_55[267]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[60],stage1_57[80],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2163 (
      {stage0_55[268], stage0_55[269], stage0_55[270], stage0_55[271], stage0_55[272], stage0_55[273]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[61],stage1_57[81],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2164 (
      {stage0_55[274], stage0_55[275], stage0_55[276], stage0_55[277], stage0_55[278], stage0_55[279]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[62],stage1_57[82],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2165 (
      {stage0_55[280], stage0_55[281], stage0_55[282], stage0_55[283], stage0_55[284], stage0_55[285]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[63],stage1_57[83],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2166 (
      {stage0_55[286], stage0_55[287], stage0_55[288], stage0_55[289], stage0_55[290], stage0_55[291]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[64],stage1_57[84],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2167 (
      {stage0_55[292], stage0_55[293], stage0_55[294], stage0_55[295], stage0_55[296], stage0_55[297]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[65],stage1_57[85],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2168 (
      {stage0_55[298], stage0_55[299], stage0_55[300], stage0_55[301], stage0_55[302], stage0_55[303]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[66],stage1_57[86],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2169 (
      {stage0_55[304], stage0_55[305], stage0_55[306], stage0_55[307], stage0_55[308], stage0_55[309]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[67],stage1_57[87],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2170 (
      {stage0_55[310], stage0_55[311], stage0_55[312], stage0_55[313], stage0_55[314], stage0_55[315]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[68],stage1_57[88],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2171 (
      {stage0_55[316], stage0_55[317], stage0_55[318], stage0_55[319], stage0_55[320], stage0_55[321]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[69],stage1_57[89],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2172 (
      {stage0_55[322], stage0_55[323], stage0_55[324], stage0_55[325], stage0_55[326], stage0_55[327]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[70],stage1_57[90],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2173 (
      {stage0_55[328], stage0_55[329], stage0_55[330], stage0_55[331], stage0_55[332], stage0_55[333]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[71],stage1_57[91],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2174 (
      {stage0_55[334], stage0_55[335], stage0_55[336], stage0_55[337], stage0_55[338], stage0_55[339]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[72],stage1_57[92],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2175 (
      {stage0_55[340], stage0_55[341], stage0_55[342], stage0_55[343], stage0_55[344], stage0_55[345]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[73],stage1_57[93],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2176 (
      {stage0_55[346], stage0_55[347], stage0_55[348], stage0_55[349], stage0_55[350], stage0_55[351]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[74],stage1_57[94],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2177 (
      {stage0_55[352], stage0_55[353], stage0_55[354], stage0_55[355], stage0_55[356], stage0_55[357]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[75],stage1_57[95],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2178 (
      {stage0_55[358], stage0_55[359], stage0_55[360], stage0_55[361], stage0_55[362], stage0_55[363]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[76],stage1_57[96],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2179 (
      {stage0_55[364], stage0_55[365], stage0_55[366], stage0_55[367], stage0_55[368], stage0_55[369]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[77],stage1_57[97],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2180 (
      {stage0_55[370], stage0_55[371], stage0_55[372], stage0_55[373], stage0_55[374], stage0_55[375]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[78],stage1_57[98],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2181 (
      {stage0_55[376], stage0_55[377], stage0_55[378], stage0_55[379], stage0_55[380], stage0_55[381]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[79],stage1_57[99],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2182 (
      {stage0_55[382], stage0_55[383], stage0_55[384], stage0_55[385], stage0_55[386], stage0_55[387]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[80],stage1_57[100],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2183 (
      {stage0_55[388], stage0_55[389], stage0_55[390], stage0_55[391], stage0_55[392], stage0_55[393]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[81],stage1_57[101],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2184 (
      {stage0_55[394], stage0_55[395], stage0_55[396], stage0_55[397], stage0_55[398], stage0_55[399]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[82],stage1_57[102],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2185 (
      {stage0_55[400], stage0_55[401], stage0_55[402], stage0_55[403], stage0_55[404], stage0_55[405]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[83],stage1_57[103],stage1_56[140],stage1_55[203]}
   );
   gpc606_5 gpc2186 (
      {stage0_55[406], stage0_55[407], stage0_55[408], stage0_55[409], stage0_55[410], stage0_55[411]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[84],stage1_57[104],stage1_56[141],stage1_55[204]}
   );
   gpc606_5 gpc2187 (
      {stage0_55[412], stage0_55[413], stage0_55[414], stage0_55[415], stage0_55[416], stage0_55[417]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[85],stage1_57[105],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2188 (
      {stage0_55[418], stage0_55[419], stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[86],stage1_57[106],stage1_56[143],stage1_55[206]}
   );
   gpc606_5 gpc2189 (
      {stage0_55[424], stage0_55[425], stage0_55[426], stage0_55[427], stage0_55[428], stage0_55[429]},
      {stage0_57[264], stage0_57[265], stage0_57[266], stage0_57[267], stage0_57[268], stage0_57[269]},
      {stage1_59[44],stage1_58[87],stage1_57[107],stage1_56[144],stage1_55[207]}
   );
   gpc606_5 gpc2190 (
      {stage0_55[430], stage0_55[431], stage0_55[432], stage0_55[433], stage0_55[434], stage0_55[435]},
      {stage0_57[270], stage0_57[271], stage0_57[272], stage0_57[273], stage0_57[274], stage0_57[275]},
      {stage1_59[45],stage1_58[88],stage1_57[108],stage1_56[145],stage1_55[208]}
   );
   gpc606_5 gpc2191 (
      {stage0_55[436], stage0_55[437], stage0_55[438], stage0_55[439], stage0_55[440], stage0_55[441]},
      {stage0_57[276], stage0_57[277], stage0_57[278], stage0_57[279], stage0_57[280], stage0_57[281]},
      {stage1_59[46],stage1_58[89],stage1_57[109],stage1_56[146],stage1_55[209]}
   );
   gpc606_5 gpc2192 (
      {stage0_55[442], stage0_55[443], stage0_55[444], stage0_55[445], stage0_55[446], stage0_55[447]},
      {stage0_57[282], stage0_57[283], stage0_57[284], stage0_57[285], stage0_57[286], stage0_57[287]},
      {stage1_59[47],stage1_58[90],stage1_57[110],stage1_56[147],stage1_55[210]}
   );
   gpc606_5 gpc2193 (
      {stage0_55[448], stage0_55[449], stage0_55[450], stage0_55[451], stage0_55[452], stage0_55[453]},
      {stage0_57[288], stage0_57[289], stage0_57[290], stage0_57[291], stage0_57[292], stage0_57[293]},
      {stage1_59[48],stage1_58[91],stage1_57[111],stage1_56[148],stage1_55[211]}
   );
   gpc606_5 gpc2194 (
      {stage0_55[454], stage0_55[455], stage0_55[456], stage0_55[457], stage0_55[458], stage0_55[459]},
      {stage0_57[294], stage0_57[295], stage0_57[296], stage0_57[297], stage0_57[298], stage0_57[299]},
      {stage1_59[49],stage1_58[92],stage1_57[112],stage1_56[149],stage1_55[212]}
   );
   gpc606_5 gpc2195 (
      {stage0_55[460], stage0_55[461], stage0_55[462], stage0_55[463], stage0_55[464], stage0_55[465]},
      {stage0_57[300], stage0_57[301], stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305]},
      {stage1_59[50],stage1_58[93],stage1_57[113],stage1_56[150],stage1_55[213]}
   );
   gpc606_5 gpc2196 (
      {stage0_55[466], stage0_55[467], stage0_55[468], stage0_55[469], stage0_55[470], stage0_55[471]},
      {stage0_57[306], stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage1_59[51],stage1_58[94],stage1_57[114],stage1_56[151],stage1_55[214]}
   );
   gpc606_5 gpc2197 (
      {stage0_55[472], stage0_55[473], stage0_55[474], stage0_55[475], stage0_55[476], stage0_55[477]},
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316], stage0_57[317]},
      {stage1_59[52],stage1_58[95],stage1_57[115],stage1_56[152],stage1_55[215]}
   );
   gpc615_5 gpc2198 (
      {stage0_55[478], stage0_55[479], stage0_55[480], stage0_55[481], stage0_55[482]},
      {stage0_56[258]},
      {stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321], stage0_57[322], stage0_57[323]},
      {stage1_59[53],stage1_58[96],stage1_57[116],stage1_56[153],stage1_55[216]}
   );
   gpc615_5 gpc2199 (
      {stage0_55[483], stage0_55[484], stage0_55[485], stage0_55[486], stage0_55[487]},
      {stage0_56[259]},
      {stage0_57[324], stage0_57[325], stage0_57[326], stage0_57[327], stage0_57[328], stage0_57[329]},
      {stage1_59[54],stage1_58[97],stage1_57[117],stage1_56[154],stage1_55[217]}
   );
   gpc615_5 gpc2200 (
      {stage0_55[488], stage0_55[489], stage0_55[490], stage0_55[491], stage0_55[492]},
      {stage0_56[260]},
      {stage0_57[330], stage0_57[331], stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335]},
      {stage1_59[55],stage1_58[98],stage1_57[118],stage1_56[155],stage1_55[218]}
   );
   gpc615_5 gpc2201 (
      {stage0_55[493], stage0_55[494], stage0_55[495], stage0_55[496], stage0_55[497]},
      {stage0_56[261]},
      {stage0_57[336], stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage1_59[56],stage1_58[99],stage1_57[119],stage1_56[156],stage1_55[219]}
   );
   gpc615_5 gpc2202 (
      {stage0_55[498], stage0_55[499], stage0_55[500], stage0_55[501], stage0_55[502]},
      {stage0_56[262]},
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346], stage0_57[347]},
      {stage1_59[57],stage1_58[100],stage1_57[120],stage1_56[157],stage1_55[220]}
   );
   gpc615_5 gpc2203 (
      {stage0_55[503], stage0_55[504], stage0_55[505], stage0_55[506], stage0_55[507]},
      {stage0_56[263]},
      {stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351], stage0_57[352], stage0_57[353]},
      {stage1_59[58],stage1_58[101],stage1_57[121],stage1_56[158],stage1_55[221]}
   );
   gpc606_5 gpc2204 (
      {stage0_56[264], stage0_56[265], stage0_56[266], stage0_56[267], stage0_56[268], stage0_56[269]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[59],stage1_58[102],stage1_57[122],stage1_56[159]}
   );
   gpc606_5 gpc2205 (
      {stage0_56[270], stage0_56[271], stage0_56[272], stage0_56[273], stage0_56[274], stage0_56[275]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[60],stage1_58[103],stage1_57[123],stage1_56[160]}
   );
   gpc606_5 gpc2206 (
      {stage0_56[276], stage0_56[277], stage0_56[278], stage0_56[279], stage0_56[280], stage0_56[281]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[61],stage1_58[104],stage1_57[124],stage1_56[161]}
   );
   gpc606_5 gpc2207 (
      {stage0_56[282], stage0_56[283], stage0_56[284], stage0_56[285], stage0_56[286], stage0_56[287]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[62],stage1_58[105],stage1_57[125],stage1_56[162]}
   );
   gpc606_5 gpc2208 (
      {stage0_56[288], stage0_56[289], stage0_56[290], stage0_56[291], stage0_56[292], stage0_56[293]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[63],stage1_58[106],stage1_57[126],stage1_56[163]}
   );
   gpc606_5 gpc2209 (
      {stage0_56[294], stage0_56[295], stage0_56[296], stage0_56[297], stage0_56[298], stage0_56[299]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[64],stage1_58[107],stage1_57[127],stage1_56[164]}
   );
   gpc606_5 gpc2210 (
      {stage0_56[300], stage0_56[301], stage0_56[302], stage0_56[303], stage0_56[304], stage0_56[305]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[65],stage1_58[108],stage1_57[128],stage1_56[165]}
   );
   gpc606_5 gpc2211 (
      {stage0_56[306], stage0_56[307], stage0_56[308], stage0_56[309], stage0_56[310], stage0_56[311]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[66],stage1_58[109],stage1_57[129],stage1_56[166]}
   );
   gpc606_5 gpc2212 (
      {stage0_56[312], stage0_56[313], stage0_56[314], stage0_56[315], stage0_56[316], stage0_56[317]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[67],stage1_58[110],stage1_57[130],stage1_56[167]}
   );
   gpc606_5 gpc2213 (
      {stage0_56[318], stage0_56[319], stage0_56[320], stage0_56[321], stage0_56[322], stage0_56[323]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[68],stage1_58[111],stage1_57[131],stage1_56[168]}
   );
   gpc606_5 gpc2214 (
      {stage0_56[324], stage0_56[325], stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[69],stage1_58[112],stage1_57[132],stage1_56[169]}
   );
   gpc606_5 gpc2215 (
      {stage0_56[330], stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[70],stage1_58[113],stage1_57[133],stage1_56[170]}
   );
   gpc606_5 gpc2216 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340], stage0_56[341]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[71],stage1_58[114],stage1_57[134],stage1_56[171]}
   );
   gpc606_5 gpc2217 (
      {stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345], stage0_56[346], stage0_56[347]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[72],stage1_58[115],stage1_57[135],stage1_56[172]}
   );
   gpc606_5 gpc2218 (
      {stage0_56[348], stage0_56[349], stage0_56[350], stage0_56[351], stage0_56[352], stage0_56[353]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[73],stage1_58[116],stage1_57[136],stage1_56[173]}
   );
   gpc606_5 gpc2219 (
      {stage0_56[354], stage0_56[355], stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[74],stage1_58[117],stage1_57[137],stage1_56[174]}
   );
   gpc606_5 gpc2220 (
      {stage0_56[360], stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[75],stage1_58[118],stage1_57[138],stage1_56[175]}
   );
   gpc606_5 gpc2221 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370], stage0_56[371]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[76],stage1_58[119],stage1_57[139],stage1_56[176]}
   );
   gpc606_5 gpc2222 (
      {stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375], stage0_56[376], stage0_56[377]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[77],stage1_58[120],stage1_57[140],stage1_56[177]}
   );
   gpc606_5 gpc2223 (
      {stage0_56[378], stage0_56[379], stage0_56[380], stage0_56[381], stage0_56[382], stage0_56[383]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[78],stage1_58[121],stage1_57[141],stage1_56[178]}
   );
   gpc606_5 gpc2224 (
      {stage0_56[384], stage0_56[385], stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[79],stage1_58[122],stage1_57[142],stage1_56[179]}
   );
   gpc606_5 gpc2225 (
      {stage0_56[390], stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[80],stage1_58[123],stage1_57[143],stage1_56[180]}
   );
   gpc606_5 gpc2226 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400], stage0_56[401]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[81],stage1_58[124],stage1_57[144],stage1_56[181]}
   );
   gpc606_5 gpc2227 (
      {stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405], stage0_56[406], stage0_56[407]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[82],stage1_58[125],stage1_57[145],stage1_56[182]}
   );
   gpc606_5 gpc2228 (
      {stage0_56[408], stage0_56[409], stage0_56[410], stage0_56[411], stage0_56[412], stage0_56[413]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[83],stage1_58[126],stage1_57[146],stage1_56[183]}
   );
   gpc606_5 gpc2229 (
      {stage0_56[414], stage0_56[415], stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[84],stage1_58[127],stage1_57[147],stage1_56[184]}
   );
   gpc606_5 gpc2230 (
      {stage0_56[420], stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[85],stage1_58[128],stage1_57[148],stage1_56[185]}
   );
   gpc606_5 gpc2231 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430], stage0_56[431]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[86],stage1_58[129],stage1_57[149],stage1_56[186]}
   );
   gpc606_5 gpc2232 (
      {stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435], stage0_56[436], stage0_56[437]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[87],stage1_58[130],stage1_57[150],stage1_56[187]}
   );
   gpc606_5 gpc2233 (
      {stage0_56[438], stage0_56[439], stage0_56[440], stage0_56[441], stage0_56[442], stage0_56[443]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[88],stage1_58[131],stage1_57[151],stage1_56[188]}
   );
   gpc606_5 gpc2234 (
      {stage0_57[354], stage0_57[355], stage0_57[356], stage0_57[357], stage0_57[358], stage0_57[359]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[30],stage1_59[89],stage1_58[132],stage1_57[152]}
   );
   gpc606_5 gpc2235 (
      {stage0_57[360], stage0_57[361], stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[31],stage1_59[90],stage1_58[133],stage1_57[153]}
   );
   gpc606_5 gpc2236 (
      {stage0_57[366], stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[32],stage1_59[91],stage1_58[134],stage1_57[154]}
   );
   gpc606_5 gpc2237 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376], stage0_57[377]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[33],stage1_59[92],stage1_58[135],stage1_57[155]}
   );
   gpc606_5 gpc2238 (
      {stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381], stage0_57[382], stage0_57[383]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[34],stage1_59[93],stage1_58[136],stage1_57[156]}
   );
   gpc606_5 gpc2239 (
      {stage0_57[384], stage0_57[385], stage0_57[386], stage0_57[387], stage0_57[388], stage0_57[389]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[35],stage1_59[94],stage1_58[137],stage1_57[157]}
   );
   gpc606_5 gpc2240 (
      {stage0_57[390], stage0_57[391], stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[36],stage1_59[95],stage1_58[138],stage1_57[158]}
   );
   gpc606_5 gpc2241 (
      {stage0_57[396], stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[37],stage1_59[96],stage1_58[139],stage1_57[159]}
   );
   gpc606_5 gpc2242 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406], stage0_57[407]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[38],stage1_59[97],stage1_58[140],stage1_57[160]}
   );
   gpc606_5 gpc2243 (
      {stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411], stage0_57[412], stage0_57[413]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[39],stage1_59[98],stage1_58[141],stage1_57[161]}
   );
   gpc606_5 gpc2244 (
      {stage0_57[414], stage0_57[415], stage0_57[416], stage0_57[417], stage0_57[418], stage0_57[419]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[40],stage1_59[99],stage1_58[142],stage1_57[162]}
   );
   gpc606_5 gpc2245 (
      {stage0_57[420], stage0_57[421], stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[41],stage1_59[100],stage1_58[143],stage1_57[163]}
   );
   gpc606_5 gpc2246 (
      {stage0_57[426], stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[42],stage1_59[101],stage1_58[144],stage1_57[164]}
   );
   gpc606_5 gpc2247 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436], stage0_57[437]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[43],stage1_59[102],stage1_58[145],stage1_57[165]}
   );
   gpc606_5 gpc2248 (
      {stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441], stage0_57[442], stage0_57[443]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[44],stage1_59[103],stage1_58[146],stage1_57[166]}
   );
   gpc606_5 gpc2249 (
      {stage0_57[444], stage0_57[445], stage0_57[446], stage0_57[447], stage0_57[448], stage0_57[449]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[45],stage1_59[104],stage1_58[147],stage1_57[167]}
   );
   gpc606_5 gpc2250 (
      {stage0_57[450], stage0_57[451], stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[46],stage1_59[105],stage1_58[148],stage1_57[168]}
   );
   gpc606_5 gpc2251 (
      {stage0_57[456], stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[47],stage1_59[106],stage1_58[149],stage1_57[169]}
   );
   gpc606_5 gpc2252 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466], stage0_57[467]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[48],stage1_59[107],stage1_58[150],stage1_57[170]}
   );
   gpc606_5 gpc2253 (
      {stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471], stage0_57[472], stage0_57[473]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[49],stage1_59[108],stage1_58[151],stage1_57[171]}
   );
   gpc606_5 gpc2254 (
      {stage0_57[474], stage0_57[475], stage0_57[476], stage0_57[477], stage0_57[478], stage0_57[479]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[50],stage1_59[109],stage1_58[152],stage1_57[172]}
   );
   gpc606_5 gpc2255 (
      {stage0_57[480], stage0_57[481], stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[51],stage1_59[110],stage1_58[153],stage1_57[173]}
   );
   gpc606_5 gpc2256 (
      {stage0_57[486], stage0_57[487], stage0_57[488], stage0_57[489], stage0_57[490], stage0_57[491]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[52],stage1_59[111],stage1_58[154],stage1_57[174]}
   );
   gpc606_5 gpc2257 (
      {stage0_57[492], stage0_57[493], stage0_57[494], stage0_57[495], stage0_57[496], stage0_57[497]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[53],stage1_59[112],stage1_58[155],stage1_57[175]}
   );
   gpc606_5 gpc2258 (
      {stage0_57[498], stage0_57[499], stage0_57[500], stage0_57[501], stage0_57[502], stage0_57[503]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[54],stage1_59[113],stage1_58[156],stage1_57[176]}
   );
   gpc606_5 gpc2259 (
      {stage0_57[504], stage0_57[505], stage0_57[506], stage0_57[507], stage0_57[508], stage0_57[509]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[55],stage1_59[114],stage1_58[157],stage1_57[177]}
   );
   gpc2135_5 gpc2260 (
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184]},
      {stage0_59[156], stage0_59[157], stage0_59[158]},
      {stage0_60[0]},
      {stage0_61[0], stage0_61[1]},
      {stage1_62[0],stage1_61[26],stage1_60[56],stage1_59[115],stage1_58[158]}
   );
   gpc2135_5 gpc2261 (
      {stage0_58[185], stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189]},
      {stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage0_60[1]},
      {stage0_61[2], stage0_61[3]},
      {stage1_62[1],stage1_61[27],stage1_60[57],stage1_59[116],stage1_58[159]}
   );
   gpc2135_5 gpc2262 (
      {stage0_58[190], stage0_58[191], stage0_58[192], stage0_58[193], stage0_58[194]},
      {stage0_59[162], stage0_59[163], stage0_59[164]},
      {stage0_60[2]},
      {stage0_61[4], stage0_61[5]},
      {stage1_62[2],stage1_61[28],stage1_60[58],stage1_59[117],stage1_58[160]}
   );
   gpc2135_5 gpc2263 (
      {stage0_58[195], stage0_58[196], stage0_58[197], stage0_58[198], stage0_58[199]},
      {stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage0_60[3]},
      {stage0_61[6], stage0_61[7]},
      {stage1_62[3],stage1_61[29],stage1_60[59],stage1_59[118],stage1_58[161]}
   );
   gpc2135_5 gpc2264 (
      {stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203], stage0_58[204]},
      {stage0_59[168], stage0_59[169], stage0_59[170]},
      {stage0_60[4]},
      {stage0_61[8], stage0_61[9]},
      {stage1_62[4],stage1_61[30],stage1_60[60],stage1_59[119],stage1_58[162]}
   );
   gpc2135_5 gpc2265 (
      {stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage0_60[5]},
      {stage0_61[10], stage0_61[11]},
      {stage1_62[5],stage1_61[31],stage1_60[61],stage1_59[120],stage1_58[163]}
   );
   gpc2135_5 gpc2266 (
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214]},
      {stage0_59[174], stage0_59[175], stage0_59[176]},
      {stage0_60[6]},
      {stage0_61[12], stage0_61[13]},
      {stage1_62[6],stage1_61[32],stage1_60[62],stage1_59[121],stage1_58[164]}
   );
   gpc2135_5 gpc2267 (
      {stage0_58[215], stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219]},
      {stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage0_60[7]},
      {stage0_61[14], stage0_61[15]},
      {stage1_62[7],stage1_61[33],stage1_60[63],stage1_59[122],stage1_58[165]}
   );
   gpc2135_5 gpc2268 (
      {stage0_58[220], stage0_58[221], stage0_58[222], stage0_58[223], stage0_58[224]},
      {stage0_59[180], stage0_59[181], stage0_59[182]},
      {stage0_60[8]},
      {stage0_61[16], stage0_61[17]},
      {stage1_62[8],stage1_61[34],stage1_60[64],stage1_59[123],stage1_58[166]}
   );
   gpc2135_5 gpc2269 (
      {stage0_58[225], stage0_58[226], stage0_58[227], stage0_58[228], stage0_58[229]},
      {stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage0_60[9]},
      {stage0_61[18], stage0_61[19]},
      {stage1_62[9],stage1_61[35],stage1_60[65],stage1_59[124],stage1_58[167]}
   );
   gpc2135_5 gpc2270 (
      {stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233], stage0_58[234]},
      {stage0_59[186], stage0_59[187], stage0_59[188]},
      {stage0_60[10]},
      {stage0_61[20], stage0_61[21]},
      {stage1_62[10],stage1_61[36],stage1_60[66],stage1_59[125],stage1_58[168]}
   );
   gpc2135_5 gpc2271 (
      {stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage0_60[11]},
      {stage0_61[22], stage0_61[23]},
      {stage1_62[11],stage1_61[37],stage1_60[67],stage1_59[126],stage1_58[169]}
   );
   gpc2135_5 gpc2272 (
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244]},
      {stage0_59[192], stage0_59[193], stage0_59[194]},
      {stage0_60[12]},
      {stage0_61[24], stage0_61[25]},
      {stage1_62[12],stage1_61[38],stage1_60[68],stage1_59[127],stage1_58[170]}
   );
   gpc2135_5 gpc2273 (
      {stage0_58[245], stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249]},
      {stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage0_60[13]},
      {stage0_61[26], stage0_61[27]},
      {stage1_62[13],stage1_61[39],stage1_60[69],stage1_59[128],stage1_58[171]}
   );
   gpc2135_5 gpc2274 (
      {stage0_58[250], stage0_58[251], stage0_58[252], stage0_58[253], stage0_58[254]},
      {stage0_59[198], stage0_59[199], stage0_59[200]},
      {stage0_60[14]},
      {stage0_61[28], stage0_61[29]},
      {stage1_62[14],stage1_61[40],stage1_60[70],stage1_59[129],stage1_58[172]}
   );
   gpc2135_5 gpc2275 (
      {stage0_58[255], stage0_58[256], stage0_58[257], stage0_58[258], stage0_58[259]},
      {stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage0_60[15]},
      {stage0_61[30], stage0_61[31]},
      {stage1_62[15],stage1_61[41],stage1_60[71],stage1_59[130],stage1_58[173]}
   );
   gpc1163_5 gpc2276 (
      {stage0_58[260], stage0_58[261], stage0_58[262]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage0_60[16]},
      {stage0_61[32]},
      {stage1_62[16],stage1_61[42],stage1_60[72],stage1_59[131],stage1_58[174]}
   );
   gpc1163_5 gpc2277 (
      {stage0_58[263], stage0_58[264], stage0_58[265]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage0_60[17]},
      {stage0_61[33]},
      {stage1_62[17],stage1_61[43],stage1_60[73],stage1_59[132],stage1_58[175]}
   );
   gpc1163_5 gpc2278 (
      {stage0_58[266], stage0_58[267], stage0_58[268]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage0_60[18]},
      {stage0_61[34]},
      {stage1_62[18],stage1_61[44],stage1_60[74],stage1_59[133],stage1_58[176]}
   );
   gpc1163_5 gpc2279 (
      {stage0_58[269], stage0_58[270], stage0_58[271]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage0_60[19]},
      {stage0_61[35]},
      {stage1_62[19],stage1_61[45],stage1_60[75],stage1_59[134],stage1_58[177]}
   );
   gpc1163_5 gpc2280 (
      {stage0_58[272], stage0_58[273], stage0_58[274]},
      {stage0_59[228], stage0_59[229], stage0_59[230], stage0_59[231], stage0_59[232], stage0_59[233]},
      {stage0_60[20]},
      {stage0_61[36]},
      {stage1_62[20],stage1_61[46],stage1_60[76],stage1_59[135],stage1_58[178]}
   );
   gpc1163_5 gpc2281 (
      {stage0_58[275], stage0_58[276], stage0_58[277]},
      {stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238], stage0_59[239]},
      {stage0_60[21]},
      {stage0_61[37]},
      {stage1_62[21],stage1_61[47],stage1_60[77],stage1_59[136],stage1_58[179]}
   );
   gpc1163_5 gpc2282 (
      {stage0_58[278], stage0_58[279], stage0_58[280]},
      {stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[22]},
      {stage0_61[38]},
      {stage1_62[22],stage1_61[48],stage1_60[78],stage1_59[137],stage1_58[180]}
   );
   gpc1163_5 gpc2283 (
      {stage0_58[281], stage0_58[282], stage0_58[283]},
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251]},
      {stage0_60[23]},
      {stage0_61[39]},
      {stage1_62[23],stage1_61[49],stage1_60[79],stage1_59[138],stage1_58[181]}
   );
   gpc1163_5 gpc2284 (
      {stage0_58[284], stage0_58[285], stage0_58[286]},
      {stage0_59[252], stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257]},
      {stage0_60[24]},
      {stage0_61[40]},
      {stage1_62[24],stage1_61[50],stage1_60[80],stage1_59[139],stage1_58[182]}
   );
   gpc1163_5 gpc2285 (
      {stage0_58[287], stage0_58[288], stage0_58[289]},
      {stage0_59[258], stage0_59[259], stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263]},
      {stage0_60[25]},
      {stage0_61[41]},
      {stage1_62[25],stage1_61[51],stage1_60[81],stage1_59[140],stage1_58[183]}
   );
   gpc1163_5 gpc2286 (
      {stage0_58[290], stage0_58[291], stage0_58[292]},
      {stage0_59[264], stage0_59[265], stage0_59[266], stage0_59[267], stage0_59[268], stage0_59[269]},
      {stage0_60[26]},
      {stage0_61[42]},
      {stage1_62[26],stage1_61[52],stage1_60[82],stage1_59[141],stage1_58[184]}
   );
   gpc1163_5 gpc2287 (
      {stage0_58[293], stage0_58[294], stage0_58[295]},
      {stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273], stage0_59[274], stage0_59[275]},
      {stage0_60[27]},
      {stage0_61[43]},
      {stage1_62[27],stage1_61[53],stage1_60[83],stage1_59[142],stage1_58[185]}
   );
   gpc1163_5 gpc2288 (
      {stage0_58[296], stage0_58[297], stage0_58[298]},
      {stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280], stage0_59[281]},
      {stage0_60[28]},
      {stage0_61[44]},
      {stage1_62[28],stage1_61[54],stage1_60[84],stage1_59[143],stage1_58[186]}
   );
   gpc1163_5 gpc2289 (
      {stage0_58[299], stage0_58[300], stage0_58[301]},
      {stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[29]},
      {stage0_61[45]},
      {stage1_62[29],stage1_61[55],stage1_60[85],stage1_59[144],stage1_58[187]}
   );
   gpc1163_5 gpc2290 (
      {stage0_58[302], stage0_58[303], stage0_58[304]},
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293]},
      {stage0_60[30]},
      {stage0_61[46]},
      {stage1_62[30],stage1_61[56],stage1_60[86],stage1_59[145],stage1_58[188]}
   );
   gpc1163_5 gpc2291 (
      {stage0_58[305], stage0_58[306], stage0_58[307]},
      {stage0_59[294], stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299]},
      {stage0_60[31]},
      {stage0_61[47]},
      {stage1_62[31],stage1_61[57],stage1_60[87],stage1_59[146],stage1_58[189]}
   );
   gpc1163_5 gpc2292 (
      {stage0_58[308], stage0_58[309], stage0_58[310]},
      {stage0_59[300], stage0_59[301], stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305]},
      {stage0_60[32]},
      {stage0_61[48]},
      {stage1_62[32],stage1_61[58],stage1_60[88],stage1_59[147],stage1_58[190]}
   );
   gpc1163_5 gpc2293 (
      {stage0_58[311], stage0_58[312], stage0_58[313]},
      {stage0_59[306], stage0_59[307], stage0_59[308], stage0_59[309], stage0_59[310], stage0_59[311]},
      {stage0_60[33]},
      {stage0_61[49]},
      {stage1_62[33],stage1_61[59],stage1_60[89],stage1_59[148],stage1_58[191]}
   );
   gpc1163_5 gpc2294 (
      {stage0_58[314], stage0_58[315], stage0_58[316]},
      {stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315], stage0_59[316], stage0_59[317]},
      {stage0_60[34]},
      {stage0_61[50]},
      {stage1_62[34],stage1_61[60],stage1_60[90],stage1_59[149],stage1_58[192]}
   );
   gpc1163_5 gpc2295 (
      {stage0_58[317], stage0_58[318], stage0_58[319]},
      {stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322], stage0_59[323]},
      {stage0_60[35]},
      {stage0_61[51]},
      {stage1_62[35],stage1_61[61],stage1_60[91],stage1_59[150],stage1_58[193]}
   );
   gpc1163_5 gpc2296 (
      {stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[36]},
      {stage0_61[52]},
      {stage1_62[36],stage1_61[62],stage1_60[92],stage1_59[151],stage1_58[194]}
   );
   gpc606_5 gpc2297 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328]},
      {stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41], stage0_60[42]},
      {stage1_62[37],stage1_61[63],stage1_60[93],stage1_59[152],stage1_58[195]}
   );
   gpc606_5 gpc2298 (
      {stage0_58[329], stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334]},
      {stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47], stage0_60[48]},
      {stage1_62[38],stage1_61[64],stage1_60[94],stage1_59[153],stage1_58[196]}
   );
   gpc606_5 gpc2299 (
      {stage0_58[335], stage0_58[336], stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340]},
      {stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53], stage0_60[54]},
      {stage1_62[39],stage1_61[65],stage1_60[95],stage1_59[154],stage1_58[197]}
   );
   gpc606_5 gpc2300 (
      {stage0_58[341], stage0_58[342], stage0_58[343], stage0_58[344], stage0_58[345], stage0_58[346]},
      {stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59], stage0_60[60]},
      {stage1_62[40],stage1_61[66],stage1_60[96],stage1_59[155],stage1_58[198]}
   );
   gpc606_5 gpc2301 (
      {stage0_58[347], stage0_58[348], stage0_58[349], stage0_58[350], stage0_58[351], stage0_58[352]},
      {stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65], stage0_60[66]},
      {stage1_62[41],stage1_61[67],stage1_60[97],stage1_59[156],stage1_58[199]}
   );
   gpc606_5 gpc2302 (
      {stage0_58[353], stage0_58[354], stage0_58[355], stage0_58[356], stage0_58[357], stage0_58[358]},
      {stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71], stage0_60[72]},
      {stage1_62[42],stage1_61[68],stage1_60[98],stage1_59[157],stage1_58[200]}
   );
   gpc606_5 gpc2303 (
      {stage0_58[359], stage0_58[360], stage0_58[361], stage0_58[362], stage0_58[363], stage0_58[364]},
      {stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77], stage0_60[78]},
      {stage1_62[43],stage1_61[69],stage1_60[99],stage1_59[158],stage1_58[201]}
   );
   gpc606_5 gpc2304 (
      {stage0_58[365], stage0_58[366], stage0_58[367], stage0_58[368], stage0_58[369], stage0_58[370]},
      {stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83], stage0_60[84]},
      {stage1_62[44],stage1_61[70],stage1_60[100],stage1_59[159],stage1_58[202]}
   );
   gpc606_5 gpc2305 (
      {stage0_58[371], stage0_58[372], stage0_58[373], stage0_58[374], stage0_58[375], stage0_58[376]},
      {stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89], stage0_60[90]},
      {stage1_62[45],stage1_61[71],stage1_60[101],stage1_59[160],stage1_58[203]}
   );
   gpc606_5 gpc2306 (
      {stage0_58[377], stage0_58[378], stage0_58[379], stage0_58[380], stage0_58[381], stage0_58[382]},
      {stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95], stage0_60[96]},
      {stage1_62[46],stage1_61[72],stage1_60[102],stage1_59[161],stage1_58[204]}
   );
   gpc606_5 gpc2307 (
      {stage0_58[383], stage0_58[384], stage0_58[385], stage0_58[386], stage0_58[387], stage0_58[388]},
      {stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101], stage0_60[102]},
      {stage1_62[47],stage1_61[73],stage1_60[103],stage1_59[162],stage1_58[205]}
   );
   gpc606_5 gpc2308 (
      {stage0_58[389], stage0_58[390], stage0_58[391], stage0_58[392], stage0_58[393], stage0_58[394]},
      {stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107], stage0_60[108]},
      {stage1_62[48],stage1_61[74],stage1_60[104],stage1_59[163],stage1_58[206]}
   );
   gpc606_5 gpc2309 (
      {stage0_58[395], stage0_58[396], stage0_58[397], stage0_58[398], stage0_58[399], stage0_58[400]},
      {stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113], stage0_60[114]},
      {stage1_62[49],stage1_61[75],stage1_60[105],stage1_59[164],stage1_58[207]}
   );
   gpc606_5 gpc2310 (
      {stage0_58[401], stage0_58[402], stage0_58[403], stage0_58[404], stage0_58[405], stage0_58[406]},
      {stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119], stage0_60[120]},
      {stage1_62[50],stage1_61[76],stage1_60[106],stage1_59[165],stage1_58[208]}
   );
   gpc606_5 gpc2311 (
      {stage0_58[407], stage0_58[408], stage0_58[409], stage0_58[410], stage0_58[411], stage0_58[412]},
      {stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125], stage0_60[126]},
      {stage1_62[51],stage1_61[77],stage1_60[107],stage1_59[166],stage1_58[209]}
   );
   gpc606_5 gpc2312 (
      {stage0_58[413], stage0_58[414], stage0_58[415], stage0_58[416], stage0_58[417], stage0_58[418]},
      {stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131], stage0_60[132]},
      {stage1_62[52],stage1_61[78],stage1_60[108],stage1_59[167],stage1_58[210]}
   );
   gpc606_5 gpc2313 (
      {stage0_58[419], stage0_58[420], stage0_58[421], stage0_58[422], stage0_58[423], stage0_58[424]},
      {stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138]},
      {stage1_62[53],stage1_61[79],stage1_60[109],stage1_59[168],stage1_58[211]}
   );
   gpc606_5 gpc2314 (
      {stage0_58[425], stage0_58[426], stage0_58[427], stage0_58[428], stage0_58[429], stage0_58[430]},
      {stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144]},
      {stage1_62[54],stage1_61[80],stage1_60[110],stage1_59[169],stage1_58[212]}
   );
   gpc606_5 gpc2315 (
      {stage0_58[431], stage0_58[432], stage0_58[433], stage0_58[434], stage0_58[435], stage0_58[436]},
      {stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage1_62[55],stage1_61[81],stage1_60[111],stage1_59[170],stage1_58[213]}
   );
   gpc606_5 gpc2316 (
      {stage0_58[437], stage0_58[438], stage0_58[439], stage0_58[440], stage0_58[441], stage0_58[442]},
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155], stage0_60[156]},
      {stage1_62[56],stage1_61[82],stage1_60[112],stage1_59[171],stage1_58[214]}
   );
   gpc606_5 gpc2317 (
      {stage0_58[443], stage0_58[444], stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448]},
      {stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161], stage0_60[162]},
      {stage1_62[57],stage1_61[83],stage1_60[113],stage1_59[172],stage1_58[215]}
   );
   gpc606_5 gpc2318 (
      {stage0_58[449], stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_60[163], stage0_60[164], stage0_60[165], stage0_60[166], stage0_60[167], stage0_60[168]},
      {stage1_62[58],stage1_61[84],stage1_60[114],stage1_59[173],stage1_58[216]}
   );
   gpc606_5 gpc2319 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459], stage0_58[460]},
      {stage0_60[169], stage0_60[170], stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174]},
      {stage1_62[59],stage1_61[85],stage1_60[115],stage1_59[174],stage1_58[217]}
   );
   gpc606_5 gpc2320 (
      {stage0_58[461], stage0_58[462], stage0_58[463], stage0_58[464], stage0_58[465], stage0_58[466]},
      {stage0_60[175], stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage1_62[60],stage1_61[86],stage1_60[116],stage1_59[175],stage1_58[218]}
   );
   gpc606_5 gpc2321 (
      {stage0_58[467], stage0_58[468], stage0_58[469], stage0_58[470], stage0_58[471], stage0_58[472]},
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185], stage0_60[186]},
      {stage1_62[61],stage1_61[87],stage1_60[117],stage1_59[176],stage1_58[219]}
   );
   gpc615_5 gpc2322 (
      {stage0_58[473], stage0_58[474], stage0_58[475], stage0_58[476], stage0_58[477]},
      {stage0_59[330]},
      {stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190], stage0_60[191], stage0_60[192]},
      {stage1_62[62],stage1_61[88],stage1_60[118],stage1_59[177],stage1_58[220]}
   );
   gpc615_5 gpc2323 (
      {stage0_58[478], stage0_58[479], stage0_58[480], stage0_58[481], stage0_58[482]},
      {stage0_59[331]},
      {stage0_60[193], stage0_60[194], stage0_60[195], stage0_60[196], stage0_60[197], stage0_60[198]},
      {stage1_62[63],stage1_61[89],stage1_60[119],stage1_59[178],stage1_58[221]}
   );
   gpc615_5 gpc2324 (
      {stage0_58[483], stage0_58[484], stage0_58[485], stage0_58[486], stage0_58[487]},
      {stage0_59[332]},
      {stage0_60[199], stage0_60[200], stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204]},
      {stage1_62[64],stage1_61[90],stage1_60[120],stage1_59[179],stage1_58[222]}
   );
   gpc615_5 gpc2325 (
      {stage0_58[488], stage0_58[489], stage0_58[490], stage0_58[491], stage0_58[492]},
      {stage0_59[333]},
      {stage0_60[205], stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage1_62[65],stage1_61[91],stage1_60[121],stage1_59[180],stage1_58[223]}
   );
   gpc606_5 gpc2326 (
      {stage0_59[334], stage0_59[335], stage0_59[336], stage0_59[337], stage0_59[338], stage0_59[339]},
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58]},
      {stage1_63[0],stage1_62[66],stage1_61[92],stage1_60[122],stage1_59[181]}
   );
   gpc606_5 gpc2327 (
      {stage0_59[340], stage0_59[341], stage0_59[342], stage0_59[343], stage0_59[344], stage0_59[345]},
      {stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64]},
      {stage1_63[1],stage1_62[67],stage1_61[93],stage1_60[123],stage1_59[182]}
   );
   gpc606_5 gpc2328 (
      {stage0_59[346], stage0_59[347], stage0_59[348], stage0_59[349], stage0_59[350], stage0_59[351]},
      {stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70]},
      {stage1_63[2],stage1_62[68],stage1_61[94],stage1_60[124],stage1_59[183]}
   );
   gpc606_5 gpc2329 (
      {stage0_59[352], stage0_59[353], stage0_59[354], stage0_59[355], stage0_59[356], stage0_59[357]},
      {stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76]},
      {stage1_63[3],stage1_62[69],stage1_61[95],stage1_60[125],stage1_59[184]}
   );
   gpc606_5 gpc2330 (
      {stage0_59[358], stage0_59[359], stage0_59[360], stage0_59[361], stage0_59[362], stage0_59[363]},
      {stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82]},
      {stage1_63[4],stage1_62[70],stage1_61[96],stage1_60[126],stage1_59[185]}
   );
   gpc606_5 gpc2331 (
      {stage0_59[364], stage0_59[365], stage0_59[366], stage0_59[367], stage0_59[368], stage0_59[369]},
      {stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88]},
      {stage1_63[5],stage1_62[71],stage1_61[97],stage1_60[127],stage1_59[186]}
   );
   gpc606_5 gpc2332 (
      {stage0_59[370], stage0_59[371], stage0_59[372], stage0_59[373], stage0_59[374], stage0_59[375]},
      {stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94]},
      {stage1_63[6],stage1_62[72],stage1_61[98],stage1_60[128],stage1_59[187]}
   );
   gpc606_5 gpc2333 (
      {stage0_59[376], stage0_59[377], stage0_59[378], stage0_59[379], stage0_59[380], stage0_59[381]},
      {stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100]},
      {stage1_63[7],stage1_62[73],stage1_61[99],stage1_60[129],stage1_59[188]}
   );
   gpc606_5 gpc2334 (
      {stage0_59[382], stage0_59[383], stage0_59[384], stage0_59[385], stage0_59[386], stage0_59[387]},
      {stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106]},
      {stage1_63[8],stage1_62[74],stage1_61[100],stage1_60[130],stage1_59[189]}
   );
   gpc606_5 gpc2335 (
      {stage0_59[388], stage0_59[389], stage0_59[390], stage0_59[391], stage0_59[392], stage0_59[393]},
      {stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112]},
      {stage1_63[9],stage1_62[75],stage1_61[101],stage1_60[131],stage1_59[190]}
   );
   gpc606_5 gpc2336 (
      {stage0_59[394], stage0_59[395], stage0_59[396], stage0_59[397], stage0_59[398], stage0_59[399]},
      {stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118]},
      {stage1_63[10],stage1_62[76],stage1_61[102],stage1_60[132],stage1_59[191]}
   );
   gpc606_5 gpc2337 (
      {stage0_59[400], stage0_59[401], stage0_59[402], stage0_59[403], stage0_59[404], stage0_59[405]},
      {stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124]},
      {stage1_63[11],stage1_62[77],stage1_61[103],stage1_60[133],stage1_59[192]}
   );
   gpc606_5 gpc2338 (
      {stage0_59[406], stage0_59[407], stage0_59[408], stage0_59[409], stage0_59[410], stage0_59[411]},
      {stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130]},
      {stage1_63[12],stage1_62[78],stage1_61[104],stage1_60[134],stage1_59[193]}
   );
   gpc606_5 gpc2339 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215], stage0_60[216]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[13],stage1_62[79],stage1_61[105],stage1_60[135]}
   );
   gpc606_5 gpc2340 (
      {stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220], stage0_60[221], stage0_60[222]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[14],stage1_62[80],stage1_61[106],stage1_60[136]}
   );
   gpc606_5 gpc2341 (
      {stage0_60[223], stage0_60[224], stage0_60[225], stage0_60[226], stage0_60[227], stage0_60[228]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[15],stage1_62[81],stage1_61[107],stage1_60[137]}
   );
   gpc606_5 gpc2342 (
      {stage0_60[229], stage0_60[230], stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[16],stage1_62[82],stage1_61[108],stage1_60[138]}
   );
   gpc606_5 gpc2343 (
      {stage0_60[235], stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[17],stage1_62[83],stage1_61[109],stage1_60[139]}
   );
   gpc606_5 gpc2344 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245], stage0_60[246]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[18],stage1_62[84],stage1_61[110],stage1_60[140]}
   );
   gpc606_5 gpc2345 (
      {stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250], stage0_60[251], stage0_60[252]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[19],stage1_62[85],stage1_61[111],stage1_60[141]}
   );
   gpc606_5 gpc2346 (
      {stage0_60[253], stage0_60[254], stage0_60[255], stage0_60[256], stage0_60[257], stage0_60[258]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[20],stage1_62[86],stage1_61[112],stage1_60[142]}
   );
   gpc606_5 gpc2347 (
      {stage0_60[259], stage0_60[260], stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[21],stage1_62[87],stage1_61[113],stage1_60[143]}
   );
   gpc606_5 gpc2348 (
      {stage0_60[265], stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[22],stage1_62[88],stage1_61[114],stage1_60[144]}
   );
   gpc606_5 gpc2349 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275], stage0_60[276]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[23],stage1_62[89],stage1_61[115],stage1_60[145]}
   );
   gpc606_5 gpc2350 (
      {stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280], stage0_60[281], stage0_60[282]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[24],stage1_62[90],stage1_61[116],stage1_60[146]}
   );
   gpc606_5 gpc2351 (
      {stage0_60[283], stage0_60[284], stage0_60[285], stage0_60[286], stage0_60[287], stage0_60[288]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[25],stage1_62[91],stage1_61[117],stage1_60[147]}
   );
   gpc606_5 gpc2352 (
      {stage0_60[289], stage0_60[290], stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[26],stage1_62[92],stage1_61[118],stage1_60[148]}
   );
   gpc606_5 gpc2353 (
      {stage0_60[295], stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[27],stage1_62[93],stage1_61[119],stage1_60[149]}
   );
   gpc606_5 gpc2354 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305], stage0_60[306]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[28],stage1_62[94],stage1_61[120],stage1_60[150]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310], stage0_60[311]},
      {stage0_61[131]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[29],stage1_62[95],stage1_61[121],stage1_60[151]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315], stage0_60[316]},
      {stage0_61[132]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[30],stage1_62[96],stage1_61[122],stage1_60[152]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320], stage0_60[321]},
      {stage0_61[133]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[31],stage1_62[97],stage1_61[123],stage1_60[153]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325], stage0_60[326]},
      {stage0_61[134]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[32],stage1_62[98],stage1_61[124],stage1_60[154]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330], stage0_60[331]},
      {stage0_61[135]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[33],stage1_62[99],stage1_61[125],stage1_60[155]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335], stage0_60[336]},
      {stage0_61[136]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[34],stage1_62[100],stage1_61[126],stage1_60[156]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340], stage0_60[341]},
      {stage0_61[137]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[35],stage1_62[101],stage1_61[127],stage1_60[157]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345], stage0_60[346]},
      {stage0_61[138]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[36],stage1_62[102],stage1_61[128],stage1_60[158]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350], stage0_60[351]},
      {stage0_61[139]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[37],stage1_62[103],stage1_61[129],stage1_60[159]}
   );
   gpc615_5 gpc2364 (
      {stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355], stage0_60[356]},
      {stage0_61[140]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[38],stage1_62[104],stage1_61[130],stage1_60[160]}
   );
   gpc615_5 gpc2365 (
      {stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360], stage0_60[361]},
      {stage0_61[141]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[39],stage1_62[105],stage1_61[131],stage1_60[161]}
   );
   gpc615_5 gpc2366 (
      {stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365], stage0_60[366]},
      {stage0_61[142]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[40],stage1_62[106],stage1_61[132],stage1_60[162]}
   );
   gpc615_5 gpc2367 (
      {stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370], stage0_60[371]},
      {stage0_61[143]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[41],stage1_62[107],stage1_61[133],stage1_60[163]}
   );
   gpc615_5 gpc2368 (
      {stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375], stage0_60[376]},
      {stage0_61[144]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[42],stage1_62[108],stage1_61[134],stage1_60[164]}
   );
   gpc615_5 gpc2369 (
      {stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380], stage0_60[381]},
      {stage0_61[145]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[43],stage1_62[109],stage1_61[135],stage1_60[165]}
   );
   gpc615_5 gpc2370 (
      {stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385], stage0_60[386]},
      {stage0_61[146]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[44],stage1_62[110],stage1_61[136],stage1_60[166]}
   );
   gpc615_5 gpc2371 (
      {stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390], stage0_60[391]},
      {stage0_61[147]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[45],stage1_62[111],stage1_61[137],stage1_60[167]}
   );
   gpc615_5 gpc2372 (
      {stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395], stage0_60[396]},
      {stage0_61[148]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[46],stage1_62[112],stage1_61[138],stage1_60[168]}
   );
   gpc615_5 gpc2373 (
      {stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400], stage0_60[401]},
      {stage0_61[149]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[47],stage1_62[113],stage1_61[139],stage1_60[169]}
   );
   gpc615_5 gpc2374 (
      {stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405], stage0_60[406]},
      {stage0_61[150]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[48],stage1_62[114],stage1_61[140],stage1_60[170]}
   );
   gpc615_5 gpc2375 (
      {stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410], stage0_60[411]},
      {stage0_61[151]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[49],stage1_62[115],stage1_61[141],stage1_60[171]}
   );
   gpc615_5 gpc2376 (
      {stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415], stage0_60[416]},
      {stage0_61[152]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[50],stage1_62[116],stage1_61[142],stage1_60[172]}
   );
   gpc615_5 gpc2377 (
      {stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420], stage0_60[421]},
      {stage0_61[153]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[51],stage1_62[117],stage1_61[143],stage1_60[173]}
   );
   gpc615_5 gpc2378 (
      {stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425], stage0_60[426]},
      {stage0_61[154]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[52],stage1_62[118],stage1_61[144],stage1_60[174]}
   );
   gpc615_5 gpc2379 (
      {stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430], stage0_60[431]},
      {stage0_61[155]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[53],stage1_62[119],stage1_61[145],stage1_60[175]}
   );
   gpc615_5 gpc2380 (
      {stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435], stage0_60[436]},
      {stage0_61[156]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[54],stage1_62[120],stage1_61[146],stage1_60[176]}
   );
   gpc615_5 gpc2381 (
      {stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440], stage0_60[441]},
      {stage0_61[157]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[55],stage1_62[121],stage1_61[147],stage1_60[177]}
   );
   gpc615_5 gpc2382 (
      {stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445], stage0_60[446]},
      {stage0_61[158]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[56],stage1_62[122],stage1_61[148],stage1_60[178]}
   );
   gpc615_5 gpc2383 (
      {stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450], stage0_60[451]},
      {stage0_61[159]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[57],stage1_62[123],stage1_61[149],stage1_60[179]}
   );
   gpc615_5 gpc2384 (
      {stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455], stage0_60[456]},
      {stage0_61[160]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[58],stage1_62[124],stage1_61[150],stage1_60[180]}
   );
   gpc615_5 gpc2385 (
      {stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460], stage0_60[461]},
      {stage0_61[161]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[59],stage1_62[125],stage1_61[151],stage1_60[181]}
   );
   gpc615_5 gpc2386 (
      {stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465], stage0_60[466]},
      {stage0_61[162]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[60],stage1_62[126],stage1_61[152],stage1_60[182]}
   );
   gpc615_5 gpc2387 (
      {stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470], stage0_60[471]},
      {stage0_61[163]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[61],stage1_62[127],stage1_61[153],stage1_60[183]}
   );
   gpc615_5 gpc2388 (
      {stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475], stage0_60[476]},
      {stage0_61[164]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[62],stage1_62[128],stage1_61[154],stage1_60[184]}
   );
   gpc615_5 gpc2389 (
      {stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480], stage0_60[481]},
      {stage0_61[165]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[63],stage1_62[129],stage1_61[155],stage1_60[185]}
   );
   gpc615_5 gpc2390 (
      {stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485], stage0_60[486]},
      {stage0_61[166]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[64],stage1_62[130],stage1_61[156],stage1_60[186]}
   );
   gpc615_5 gpc2391 (
      {stage0_60[487], stage0_60[488], stage0_60[489], stage0_60[490], stage0_60[491]},
      {stage0_61[167]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[65],stage1_62[131],stage1_61[157],stage1_60[187]}
   );
   gpc615_5 gpc2392 (
      {stage0_60[492], stage0_60[493], stage0_60[494], stage0_60[495], stage0_60[496]},
      {stage0_61[168]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[66],stage1_62[132],stage1_61[158],stage1_60[188]}
   );
   gpc615_5 gpc2393 (
      {stage0_60[497], stage0_60[498], stage0_60[499], stage0_60[500], stage0_60[501]},
      {stage0_61[169]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[67],stage1_62[133],stage1_61[159],stage1_60[189]}
   );
   gpc606_5 gpc2394 (
      {stage0_61[170], stage0_61[171], stage0_61[172], stage0_61[173], stage0_61[174], stage0_61[175]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[55],stage1_63[68],stage1_62[134],stage1_61[160]}
   );
   gpc606_5 gpc2395 (
      {stage0_61[176], stage0_61[177], stage0_61[178], stage0_61[179], stage0_61[180], stage0_61[181]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[56],stage1_63[69],stage1_62[135],stage1_61[161]}
   );
   gpc606_5 gpc2396 (
      {stage0_61[182], stage0_61[183], stage0_61[184], stage0_61[185], stage0_61[186], stage0_61[187]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[57],stage1_63[70],stage1_62[136],stage1_61[162]}
   );
   gpc606_5 gpc2397 (
      {stage0_61[188], stage0_61[189], stage0_61[190], stage0_61[191], stage0_61[192], stage0_61[193]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[58],stage1_63[71],stage1_62[137],stage1_61[163]}
   );
   gpc606_5 gpc2398 (
      {stage0_61[194], stage0_61[195], stage0_61[196], stage0_61[197], stage0_61[198], stage0_61[199]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[59],stage1_63[72],stage1_62[138],stage1_61[164]}
   );
   gpc606_5 gpc2399 (
      {stage0_61[200], stage0_61[201], stage0_61[202], stage0_61[203], stage0_61[204], stage0_61[205]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[60],stage1_63[73],stage1_62[139],stage1_61[165]}
   );
   gpc606_5 gpc2400 (
      {stage0_61[206], stage0_61[207], stage0_61[208], stage0_61[209], stage0_61[210], stage0_61[211]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[61],stage1_63[74],stage1_62[140],stage1_61[166]}
   );
   gpc606_5 gpc2401 (
      {stage0_61[212], stage0_61[213], stage0_61[214], stage0_61[215], stage0_61[216], stage0_61[217]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[62],stage1_63[75],stage1_62[141],stage1_61[167]}
   );
   gpc606_5 gpc2402 (
      {stage0_61[218], stage0_61[219], stage0_61[220], stage0_61[221], stage0_61[222], stage0_61[223]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[63],stage1_63[76],stage1_62[142],stage1_61[168]}
   );
   gpc606_5 gpc2403 (
      {stage0_61[224], stage0_61[225], stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[64],stage1_63[77],stage1_62[143],stage1_61[169]}
   );
   gpc606_5 gpc2404 (
      {stage0_61[230], stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[65],stage1_63[78],stage1_62[144],stage1_61[170]}
   );
   gpc606_5 gpc2405 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240], stage0_61[241]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[66],stage1_63[79],stage1_62[145],stage1_61[171]}
   );
   gpc606_5 gpc2406 (
      {stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245], stage0_61[246], stage0_61[247]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[67],stage1_63[80],stage1_62[146],stage1_61[172]}
   );
   gpc606_5 gpc2407 (
      {stage0_61[248], stage0_61[249], stage0_61[250], stage0_61[251], stage0_61[252], stage0_61[253]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[68],stage1_63[81],stage1_62[147],stage1_61[173]}
   );
   gpc606_5 gpc2408 (
      {stage0_61[254], stage0_61[255], stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[69],stage1_63[82],stage1_62[148],stage1_61[174]}
   );
   gpc606_5 gpc2409 (
      {stage0_61[260], stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[70],stage1_63[83],stage1_62[149],stage1_61[175]}
   );
   gpc606_5 gpc2410 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270], stage0_61[271]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[71],stage1_63[84],stage1_62[150],stage1_61[176]}
   );
   gpc606_5 gpc2411 (
      {stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275], stage0_61[276], stage0_61[277]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[72],stage1_63[85],stage1_62[151],stage1_61[177]}
   );
   gpc606_5 gpc2412 (
      {stage0_61[278], stage0_61[279], stage0_61[280], stage0_61[281], stage0_61[282], stage0_61[283]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[73],stage1_63[86],stage1_62[152],stage1_61[178]}
   );
   gpc606_5 gpc2413 (
      {stage0_61[284], stage0_61[285], stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[74],stage1_63[87],stage1_62[153],stage1_61[179]}
   );
   gpc606_5 gpc2414 (
      {stage0_61[290], stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[75],stage1_63[88],stage1_62[154],stage1_61[180]}
   );
   gpc606_5 gpc2415 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300], stage0_61[301]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[76],stage1_63[89],stage1_62[155],stage1_61[181]}
   );
   gpc606_5 gpc2416 (
      {stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305], stage0_61[306], stage0_61[307]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[77],stage1_63[90],stage1_62[156],stage1_61[182]}
   );
   gpc606_5 gpc2417 (
      {stage0_61[308], stage0_61[309], stage0_61[310], stage0_61[311], stage0_61[312], stage0_61[313]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[78],stage1_63[91],stage1_62[157],stage1_61[183]}
   );
   gpc606_5 gpc2418 (
      {stage0_61[314], stage0_61[315], stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[79],stage1_63[92],stage1_62[158],stage1_61[184]}
   );
   gpc606_5 gpc2419 (
      {stage0_61[320], stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[80],stage1_63[93],stage1_62[159],stage1_61[185]}
   );
   gpc606_5 gpc2420 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330], stage0_61[331]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[81],stage1_63[94],stage1_62[160],stage1_61[186]}
   );
   gpc606_5 gpc2421 (
      {stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335], stage0_61[336], stage0_61[337]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[82],stage1_63[95],stage1_62[161],stage1_61[187]}
   );
   gpc606_5 gpc2422 (
      {stage0_61[338], stage0_61[339], stage0_61[340], stage0_61[341], stage0_61[342], stage0_61[343]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[83],stage1_63[96],stage1_62[162],stage1_61[188]}
   );
   gpc606_5 gpc2423 (
      {stage0_61[344], stage0_61[345], stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[84],stage1_63[97],stage1_62[163],stage1_61[189]}
   );
   gpc606_5 gpc2424 (
      {stage0_61[350], stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[85],stage1_63[98],stage1_62[164],stage1_61[190]}
   );
   gpc606_5 gpc2425 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360], stage0_61[361]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[86],stage1_63[99],stage1_62[165],stage1_61[191]}
   );
   gpc606_5 gpc2426 (
      {stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365], stage0_61[366], stage0_61[367]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[87],stage1_63[100],stage1_62[166],stage1_61[192]}
   );
   gpc606_5 gpc2427 (
      {stage0_61[368], stage0_61[369], stage0_61[370], stage0_61[371], stage0_61[372], stage0_61[373]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[88],stage1_63[101],stage1_62[167],stage1_61[193]}
   );
   gpc606_5 gpc2428 (
      {stage0_61[374], stage0_61[375], stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[89],stage1_63[102],stage1_62[168],stage1_61[194]}
   );
   gpc606_5 gpc2429 (
      {stage0_61[380], stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[90],stage1_63[103],stage1_62[169],stage1_61[195]}
   );
   gpc606_5 gpc2430 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390], stage0_61[391]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[91],stage1_63[104],stage1_62[170],stage1_61[196]}
   );
   gpc606_5 gpc2431 (
      {stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395], stage0_61[396], stage0_61[397]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[92],stage1_63[105],stage1_62[171],stage1_61[197]}
   );
   gpc606_5 gpc2432 (
      {stage0_61[398], stage0_61[399], stage0_61[400], stage0_61[401], stage0_61[402], stage0_61[403]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[93],stage1_63[106],stage1_62[172],stage1_61[198]}
   );
   gpc606_5 gpc2433 (
      {stage0_61[404], stage0_61[405], stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[94],stage1_63[107],stage1_62[173],stage1_61[199]}
   );
   gpc606_5 gpc2434 (
      {stage0_61[410], stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[95],stage1_63[108],stage1_62[174],stage1_61[200]}
   );
   gpc606_5 gpc2435 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420], stage0_61[421]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[96],stage1_63[109],stage1_62[175],stage1_61[201]}
   );
   gpc606_5 gpc2436 (
      {stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425], stage0_61[426], stage0_61[427]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[97],stage1_63[110],stage1_62[176],stage1_61[202]}
   );
   gpc606_5 gpc2437 (
      {stage0_61[428], stage0_61[429], stage0_61[430], stage0_61[431], stage0_61[432], stage0_61[433]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[98],stage1_63[111],stage1_62[177],stage1_61[203]}
   );
   gpc606_5 gpc2438 (
      {stage0_61[434], stage0_61[435], stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[99],stage1_63[112],stage1_62[178],stage1_61[204]}
   );
   gpc606_5 gpc2439 (
      {stage0_61[440], stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[100],stage1_63[113],stage1_62[179],stage1_61[205]}
   );
   gpc606_5 gpc2440 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450], stage0_61[451]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[101],stage1_63[114],stage1_62[180],stage1_61[206]}
   );
   gpc606_5 gpc2441 (
      {stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455], stage0_61[456], stage0_61[457]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[102],stage1_63[115],stage1_62[181],stage1_61[207]}
   );
   gpc606_5 gpc2442 (
      {stage0_61[458], stage0_61[459], stage0_61[460], stage0_61[461], stage0_61[462], stage0_61[463]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[103],stage1_63[116],stage1_62[182],stage1_61[208]}
   );
   gpc606_5 gpc2443 (
      {stage0_61[464], stage0_61[465], stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[104],stage1_63[117],stage1_62[183],stage1_61[209]}
   );
   gpc606_5 gpc2444 (
      {stage0_61[470], stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[105],stage1_63[118],stage1_62[184],stage1_61[210]}
   );
   gpc606_5 gpc2445 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480], stage0_61[481]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[106],stage1_63[119],stage1_62[185],stage1_61[211]}
   );
   gpc606_5 gpc2446 (
      {stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485], stage0_61[486], stage0_61[487]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[107],stage1_63[120],stage1_62[186],stage1_61[212]}
   );
   gpc606_5 gpc2447 (
      {stage0_61[488], stage0_61[489], stage0_61[490], stage0_61[491], stage0_61[492], stage0_61[493]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[108],stage1_63[121],stage1_62[187],stage1_61[213]}
   );
   gpc606_5 gpc2448 (
      {stage0_61[494], stage0_61[495], stage0_61[496], stage0_61[497], stage0_61[498], stage0_61[499]},
      {stage0_63[324], stage0_63[325], stage0_63[326], stage0_63[327], stage0_63[328], stage0_63[329]},
      {stage1_65[54],stage1_64[109],stage1_63[122],stage1_62[188],stage1_61[214]}
   );
   gpc606_5 gpc2449 (
      {stage0_61[500], stage0_61[501], stage0_61[502], stage0_61[503], stage0_61[504], stage0_61[505]},
      {stage0_63[330], stage0_63[331], stage0_63[332], stage0_63[333], stage0_63[334], stage0_63[335]},
      {stage1_65[55],stage1_64[110],stage1_63[123],stage1_62[189],stage1_61[215]}
   );
   gpc606_5 gpc2450 (
      {stage0_61[506], stage0_61[507], stage0_61[508], stage0_61[509], stage0_61[510], stage0_61[511]},
      {stage0_63[336], stage0_63[337], stage0_63[338], stage0_63[339], stage0_63[340], stage0_63[341]},
      {stage1_65[56],stage1_64[111],stage1_63[124],stage1_62[190],stage1_61[216]}
   );
   gpc1_1 gpc2451 (
      {stage0_1[481]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2452 (
      {stage0_1[482]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2453 (
      {stage0_1[483]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2454 (
      {stage0_1[484]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2455 (
      {stage0_1[485]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[486]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[487]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[488]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[489]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[490]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[491]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[492]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[493]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[494]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[495]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[496]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[497]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[498]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[499]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[500]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[501]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[502]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[503]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[504]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[505]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[506]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[507]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[508]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[509]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[510]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[511]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2482 (
      {stage0_2[429]},
      {stage1_2[138]}
   );
   gpc1_1 gpc2483 (
      {stage0_2[430]},
      {stage1_2[139]}
   );
   gpc1_1 gpc2484 (
      {stage0_2[431]},
      {stage1_2[140]}
   );
   gpc1_1 gpc2485 (
      {stage0_2[432]},
      {stage1_2[141]}
   );
   gpc1_1 gpc2486 (
      {stage0_2[433]},
      {stage1_2[142]}
   );
   gpc1_1 gpc2487 (
      {stage0_2[434]},
      {stage1_2[143]}
   );
   gpc1_1 gpc2488 (
      {stage0_2[435]},
      {stage1_2[144]}
   );
   gpc1_1 gpc2489 (
      {stage0_2[436]},
      {stage1_2[145]}
   );
   gpc1_1 gpc2490 (
      {stage0_2[437]},
      {stage1_2[146]}
   );
   gpc1_1 gpc2491 (
      {stage0_2[438]},
      {stage1_2[147]}
   );
   gpc1_1 gpc2492 (
      {stage0_2[439]},
      {stage1_2[148]}
   );
   gpc1_1 gpc2493 (
      {stage0_2[440]},
      {stage1_2[149]}
   );
   gpc1_1 gpc2494 (
      {stage0_2[441]},
      {stage1_2[150]}
   );
   gpc1_1 gpc2495 (
      {stage0_2[442]},
      {stage1_2[151]}
   );
   gpc1_1 gpc2496 (
      {stage0_2[443]},
      {stage1_2[152]}
   );
   gpc1_1 gpc2497 (
      {stage0_2[444]},
      {stage1_2[153]}
   );
   gpc1_1 gpc2498 (
      {stage0_2[445]},
      {stage1_2[154]}
   );
   gpc1_1 gpc2499 (
      {stage0_2[446]},
      {stage1_2[155]}
   );
   gpc1_1 gpc2500 (
      {stage0_2[447]},
      {stage1_2[156]}
   );
   gpc1_1 gpc2501 (
      {stage0_2[448]},
      {stage1_2[157]}
   );
   gpc1_1 gpc2502 (
      {stage0_2[449]},
      {stage1_2[158]}
   );
   gpc1_1 gpc2503 (
      {stage0_2[450]},
      {stage1_2[159]}
   );
   gpc1_1 gpc2504 (
      {stage0_2[451]},
      {stage1_2[160]}
   );
   gpc1_1 gpc2505 (
      {stage0_2[452]},
      {stage1_2[161]}
   );
   gpc1_1 gpc2506 (
      {stage0_2[453]},
      {stage1_2[162]}
   );
   gpc1_1 gpc2507 (
      {stage0_2[454]},
      {stage1_2[163]}
   );
   gpc1_1 gpc2508 (
      {stage0_2[455]},
      {stage1_2[164]}
   );
   gpc1_1 gpc2509 (
      {stage0_2[456]},
      {stage1_2[165]}
   );
   gpc1_1 gpc2510 (
      {stage0_2[457]},
      {stage1_2[166]}
   );
   gpc1_1 gpc2511 (
      {stage0_2[458]},
      {stage1_2[167]}
   );
   gpc1_1 gpc2512 (
      {stage0_2[459]},
      {stage1_2[168]}
   );
   gpc1_1 gpc2513 (
      {stage0_2[460]},
      {stage1_2[169]}
   );
   gpc1_1 gpc2514 (
      {stage0_2[461]},
      {stage1_2[170]}
   );
   gpc1_1 gpc2515 (
      {stage0_2[462]},
      {stage1_2[171]}
   );
   gpc1_1 gpc2516 (
      {stage0_2[463]},
      {stage1_2[172]}
   );
   gpc1_1 gpc2517 (
      {stage0_2[464]},
      {stage1_2[173]}
   );
   gpc1_1 gpc2518 (
      {stage0_2[465]},
      {stage1_2[174]}
   );
   gpc1_1 gpc2519 (
      {stage0_2[466]},
      {stage1_2[175]}
   );
   gpc1_1 gpc2520 (
      {stage0_2[467]},
      {stage1_2[176]}
   );
   gpc1_1 gpc2521 (
      {stage0_2[468]},
      {stage1_2[177]}
   );
   gpc1_1 gpc2522 (
      {stage0_2[469]},
      {stage1_2[178]}
   );
   gpc1_1 gpc2523 (
      {stage0_2[470]},
      {stage1_2[179]}
   );
   gpc1_1 gpc2524 (
      {stage0_2[471]},
      {stage1_2[180]}
   );
   gpc1_1 gpc2525 (
      {stage0_2[472]},
      {stage1_2[181]}
   );
   gpc1_1 gpc2526 (
      {stage0_2[473]},
      {stage1_2[182]}
   );
   gpc1_1 gpc2527 (
      {stage0_2[474]},
      {stage1_2[183]}
   );
   gpc1_1 gpc2528 (
      {stage0_2[475]},
      {stage1_2[184]}
   );
   gpc1_1 gpc2529 (
      {stage0_2[476]},
      {stage1_2[185]}
   );
   gpc1_1 gpc2530 (
      {stage0_2[477]},
      {stage1_2[186]}
   );
   gpc1_1 gpc2531 (
      {stage0_2[478]},
      {stage1_2[187]}
   );
   gpc1_1 gpc2532 (
      {stage0_2[479]},
      {stage1_2[188]}
   );
   gpc1_1 gpc2533 (
      {stage0_2[480]},
      {stage1_2[189]}
   );
   gpc1_1 gpc2534 (
      {stage0_2[481]},
      {stage1_2[190]}
   );
   gpc1_1 gpc2535 (
      {stage0_2[482]},
      {stage1_2[191]}
   );
   gpc1_1 gpc2536 (
      {stage0_2[483]},
      {stage1_2[192]}
   );
   gpc1_1 gpc2537 (
      {stage0_2[484]},
      {stage1_2[193]}
   );
   gpc1_1 gpc2538 (
      {stage0_2[485]},
      {stage1_2[194]}
   );
   gpc1_1 gpc2539 (
      {stage0_2[486]},
      {stage1_2[195]}
   );
   gpc1_1 gpc2540 (
      {stage0_2[487]},
      {stage1_2[196]}
   );
   gpc1_1 gpc2541 (
      {stage0_2[488]},
      {stage1_2[197]}
   );
   gpc1_1 gpc2542 (
      {stage0_2[489]},
      {stage1_2[198]}
   );
   gpc1_1 gpc2543 (
      {stage0_2[490]},
      {stage1_2[199]}
   );
   gpc1_1 gpc2544 (
      {stage0_2[491]},
      {stage1_2[200]}
   );
   gpc1_1 gpc2545 (
      {stage0_2[492]},
      {stage1_2[201]}
   );
   gpc1_1 gpc2546 (
      {stage0_2[493]},
      {stage1_2[202]}
   );
   gpc1_1 gpc2547 (
      {stage0_2[494]},
      {stage1_2[203]}
   );
   gpc1_1 gpc2548 (
      {stage0_2[495]},
      {stage1_2[204]}
   );
   gpc1_1 gpc2549 (
      {stage0_2[496]},
      {stage1_2[205]}
   );
   gpc1_1 gpc2550 (
      {stage0_2[497]},
      {stage1_2[206]}
   );
   gpc1_1 gpc2551 (
      {stage0_2[498]},
      {stage1_2[207]}
   );
   gpc1_1 gpc2552 (
      {stage0_2[499]},
      {stage1_2[208]}
   );
   gpc1_1 gpc2553 (
      {stage0_2[500]},
      {stage1_2[209]}
   );
   gpc1_1 gpc2554 (
      {stage0_2[501]},
      {stage1_2[210]}
   );
   gpc1_1 gpc2555 (
      {stage0_2[502]},
      {stage1_2[211]}
   );
   gpc1_1 gpc2556 (
      {stage0_2[503]},
      {stage1_2[212]}
   );
   gpc1_1 gpc2557 (
      {stage0_2[504]},
      {stage1_2[213]}
   );
   gpc1_1 gpc2558 (
      {stage0_2[505]},
      {stage1_2[214]}
   );
   gpc1_1 gpc2559 (
      {stage0_2[506]},
      {stage1_2[215]}
   );
   gpc1_1 gpc2560 (
      {stage0_2[507]},
      {stage1_2[216]}
   );
   gpc1_1 gpc2561 (
      {stage0_2[508]},
      {stage1_2[217]}
   );
   gpc1_1 gpc2562 (
      {stage0_2[509]},
      {stage1_2[218]}
   );
   gpc1_1 gpc2563 (
      {stage0_2[510]},
      {stage1_2[219]}
   );
   gpc1_1 gpc2564 (
      {stage0_2[511]},
      {stage1_2[220]}
   );
   gpc1_1 gpc2565 (
      {stage0_3[372]},
      {stage1_3[182]}
   );
   gpc1_1 gpc2566 (
      {stage0_3[373]},
      {stage1_3[183]}
   );
   gpc1_1 gpc2567 (
      {stage0_3[374]},
      {stage1_3[184]}
   );
   gpc1_1 gpc2568 (
      {stage0_3[375]},
      {stage1_3[185]}
   );
   gpc1_1 gpc2569 (
      {stage0_3[376]},
      {stage1_3[186]}
   );
   gpc1_1 gpc2570 (
      {stage0_3[377]},
      {stage1_3[187]}
   );
   gpc1_1 gpc2571 (
      {stage0_3[378]},
      {stage1_3[188]}
   );
   gpc1_1 gpc2572 (
      {stage0_3[379]},
      {stage1_3[189]}
   );
   gpc1_1 gpc2573 (
      {stage0_3[380]},
      {stage1_3[190]}
   );
   gpc1_1 gpc2574 (
      {stage0_3[381]},
      {stage1_3[191]}
   );
   gpc1_1 gpc2575 (
      {stage0_3[382]},
      {stage1_3[192]}
   );
   gpc1_1 gpc2576 (
      {stage0_3[383]},
      {stage1_3[193]}
   );
   gpc1_1 gpc2577 (
      {stage0_3[384]},
      {stage1_3[194]}
   );
   gpc1_1 gpc2578 (
      {stage0_3[385]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2579 (
      {stage0_3[386]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2580 (
      {stage0_3[387]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2581 (
      {stage0_3[388]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2582 (
      {stage0_3[389]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2583 (
      {stage0_3[390]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2584 (
      {stage0_3[391]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2585 (
      {stage0_3[392]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2586 (
      {stage0_3[393]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2587 (
      {stage0_3[394]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2588 (
      {stage0_3[395]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2589 (
      {stage0_3[396]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2590 (
      {stage0_3[397]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2591 (
      {stage0_3[398]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2592 (
      {stage0_3[399]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2593 (
      {stage0_3[400]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2594 (
      {stage0_3[401]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2595 (
      {stage0_3[402]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2596 (
      {stage0_3[403]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2597 (
      {stage0_3[404]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2598 (
      {stage0_3[405]},
      {stage1_3[215]}
   );
   gpc1_1 gpc2599 (
      {stage0_3[406]},
      {stage1_3[216]}
   );
   gpc1_1 gpc2600 (
      {stage0_3[407]},
      {stage1_3[217]}
   );
   gpc1_1 gpc2601 (
      {stage0_3[408]},
      {stage1_3[218]}
   );
   gpc1_1 gpc2602 (
      {stage0_3[409]},
      {stage1_3[219]}
   );
   gpc1_1 gpc2603 (
      {stage0_3[410]},
      {stage1_3[220]}
   );
   gpc1_1 gpc2604 (
      {stage0_3[411]},
      {stage1_3[221]}
   );
   gpc1_1 gpc2605 (
      {stage0_3[412]},
      {stage1_3[222]}
   );
   gpc1_1 gpc2606 (
      {stage0_3[413]},
      {stage1_3[223]}
   );
   gpc1_1 gpc2607 (
      {stage0_3[414]},
      {stage1_3[224]}
   );
   gpc1_1 gpc2608 (
      {stage0_3[415]},
      {stage1_3[225]}
   );
   gpc1_1 gpc2609 (
      {stage0_3[416]},
      {stage1_3[226]}
   );
   gpc1_1 gpc2610 (
      {stage0_3[417]},
      {stage1_3[227]}
   );
   gpc1_1 gpc2611 (
      {stage0_3[418]},
      {stage1_3[228]}
   );
   gpc1_1 gpc2612 (
      {stage0_3[419]},
      {stage1_3[229]}
   );
   gpc1_1 gpc2613 (
      {stage0_3[420]},
      {stage1_3[230]}
   );
   gpc1_1 gpc2614 (
      {stage0_3[421]},
      {stage1_3[231]}
   );
   gpc1_1 gpc2615 (
      {stage0_3[422]},
      {stage1_3[232]}
   );
   gpc1_1 gpc2616 (
      {stage0_3[423]},
      {stage1_3[233]}
   );
   gpc1_1 gpc2617 (
      {stage0_3[424]},
      {stage1_3[234]}
   );
   gpc1_1 gpc2618 (
      {stage0_3[425]},
      {stage1_3[235]}
   );
   gpc1_1 gpc2619 (
      {stage0_3[426]},
      {stage1_3[236]}
   );
   gpc1_1 gpc2620 (
      {stage0_3[427]},
      {stage1_3[237]}
   );
   gpc1_1 gpc2621 (
      {stage0_3[428]},
      {stage1_3[238]}
   );
   gpc1_1 gpc2622 (
      {stage0_3[429]},
      {stage1_3[239]}
   );
   gpc1_1 gpc2623 (
      {stage0_3[430]},
      {stage1_3[240]}
   );
   gpc1_1 gpc2624 (
      {stage0_3[431]},
      {stage1_3[241]}
   );
   gpc1_1 gpc2625 (
      {stage0_3[432]},
      {stage1_3[242]}
   );
   gpc1_1 gpc2626 (
      {stage0_3[433]},
      {stage1_3[243]}
   );
   gpc1_1 gpc2627 (
      {stage0_3[434]},
      {stage1_3[244]}
   );
   gpc1_1 gpc2628 (
      {stage0_3[435]},
      {stage1_3[245]}
   );
   gpc1_1 gpc2629 (
      {stage0_3[436]},
      {stage1_3[246]}
   );
   gpc1_1 gpc2630 (
      {stage0_3[437]},
      {stage1_3[247]}
   );
   gpc1_1 gpc2631 (
      {stage0_3[438]},
      {stage1_3[248]}
   );
   gpc1_1 gpc2632 (
      {stage0_3[439]},
      {stage1_3[249]}
   );
   gpc1_1 gpc2633 (
      {stage0_3[440]},
      {stage1_3[250]}
   );
   gpc1_1 gpc2634 (
      {stage0_3[441]},
      {stage1_3[251]}
   );
   gpc1_1 gpc2635 (
      {stage0_3[442]},
      {stage1_3[252]}
   );
   gpc1_1 gpc2636 (
      {stage0_3[443]},
      {stage1_3[253]}
   );
   gpc1_1 gpc2637 (
      {stage0_3[444]},
      {stage1_3[254]}
   );
   gpc1_1 gpc2638 (
      {stage0_3[445]},
      {stage1_3[255]}
   );
   gpc1_1 gpc2639 (
      {stage0_3[446]},
      {stage1_3[256]}
   );
   gpc1_1 gpc2640 (
      {stage0_3[447]},
      {stage1_3[257]}
   );
   gpc1_1 gpc2641 (
      {stage0_3[448]},
      {stage1_3[258]}
   );
   gpc1_1 gpc2642 (
      {stage0_3[449]},
      {stage1_3[259]}
   );
   gpc1_1 gpc2643 (
      {stage0_3[450]},
      {stage1_3[260]}
   );
   gpc1_1 gpc2644 (
      {stage0_3[451]},
      {stage1_3[261]}
   );
   gpc1_1 gpc2645 (
      {stage0_3[452]},
      {stage1_3[262]}
   );
   gpc1_1 gpc2646 (
      {stage0_3[453]},
      {stage1_3[263]}
   );
   gpc1_1 gpc2647 (
      {stage0_3[454]},
      {stage1_3[264]}
   );
   gpc1_1 gpc2648 (
      {stage0_3[455]},
      {stage1_3[265]}
   );
   gpc1_1 gpc2649 (
      {stage0_3[456]},
      {stage1_3[266]}
   );
   gpc1_1 gpc2650 (
      {stage0_3[457]},
      {stage1_3[267]}
   );
   gpc1_1 gpc2651 (
      {stage0_3[458]},
      {stage1_3[268]}
   );
   gpc1_1 gpc2652 (
      {stage0_3[459]},
      {stage1_3[269]}
   );
   gpc1_1 gpc2653 (
      {stage0_3[460]},
      {stage1_3[270]}
   );
   gpc1_1 gpc2654 (
      {stage0_3[461]},
      {stage1_3[271]}
   );
   gpc1_1 gpc2655 (
      {stage0_3[462]},
      {stage1_3[272]}
   );
   gpc1_1 gpc2656 (
      {stage0_3[463]},
      {stage1_3[273]}
   );
   gpc1_1 gpc2657 (
      {stage0_3[464]},
      {stage1_3[274]}
   );
   gpc1_1 gpc2658 (
      {stage0_3[465]},
      {stage1_3[275]}
   );
   gpc1_1 gpc2659 (
      {stage0_3[466]},
      {stage1_3[276]}
   );
   gpc1_1 gpc2660 (
      {stage0_3[467]},
      {stage1_3[277]}
   );
   gpc1_1 gpc2661 (
      {stage0_3[468]},
      {stage1_3[278]}
   );
   gpc1_1 gpc2662 (
      {stage0_3[469]},
      {stage1_3[279]}
   );
   gpc1_1 gpc2663 (
      {stage0_3[470]},
      {stage1_3[280]}
   );
   gpc1_1 gpc2664 (
      {stage0_3[471]},
      {stage1_3[281]}
   );
   gpc1_1 gpc2665 (
      {stage0_3[472]},
      {stage1_3[282]}
   );
   gpc1_1 gpc2666 (
      {stage0_3[473]},
      {stage1_3[283]}
   );
   gpc1_1 gpc2667 (
      {stage0_3[474]},
      {stage1_3[284]}
   );
   gpc1_1 gpc2668 (
      {stage0_3[475]},
      {stage1_3[285]}
   );
   gpc1_1 gpc2669 (
      {stage0_3[476]},
      {stage1_3[286]}
   );
   gpc1_1 gpc2670 (
      {stage0_3[477]},
      {stage1_3[287]}
   );
   gpc1_1 gpc2671 (
      {stage0_3[478]},
      {stage1_3[288]}
   );
   gpc1_1 gpc2672 (
      {stage0_3[479]},
      {stage1_3[289]}
   );
   gpc1_1 gpc2673 (
      {stage0_3[480]},
      {stage1_3[290]}
   );
   gpc1_1 gpc2674 (
      {stage0_3[481]},
      {stage1_3[291]}
   );
   gpc1_1 gpc2675 (
      {stage0_3[482]},
      {stage1_3[292]}
   );
   gpc1_1 gpc2676 (
      {stage0_3[483]},
      {stage1_3[293]}
   );
   gpc1_1 gpc2677 (
      {stage0_3[484]},
      {stage1_3[294]}
   );
   gpc1_1 gpc2678 (
      {stage0_3[485]},
      {stage1_3[295]}
   );
   gpc1_1 gpc2679 (
      {stage0_3[486]},
      {stage1_3[296]}
   );
   gpc1_1 gpc2680 (
      {stage0_3[487]},
      {stage1_3[297]}
   );
   gpc1_1 gpc2681 (
      {stage0_3[488]},
      {stage1_3[298]}
   );
   gpc1_1 gpc2682 (
      {stage0_3[489]},
      {stage1_3[299]}
   );
   gpc1_1 gpc2683 (
      {stage0_3[490]},
      {stage1_3[300]}
   );
   gpc1_1 gpc2684 (
      {stage0_3[491]},
      {stage1_3[301]}
   );
   gpc1_1 gpc2685 (
      {stage0_3[492]},
      {stage1_3[302]}
   );
   gpc1_1 gpc2686 (
      {stage0_3[493]},
      {stage1_3[303]}
   );
   gpc1_1 gpc2687 (
      {stage0_3[494]},
      {stage1_3[304]}
   );
   gpc1_1 gpc2688 (
      {stage0_3[495]},
      {stage1_3[305]}
   );
   gpc1_1 gpc2689 (
      {stage0_3[496]},
      {stage1_3[306]}
   );
   gpc1_1 gpc2690 (
      {stage0_3[497]},
      {stage1_3[307]}
   );
   gpc1_1 gpc2691 (
      {stage0_3[498]},
      {stage1_3[308]}
   );
   gpc1_1 gpc2692 (
      {stage0_3[499]},
      {stage1_3[309]}
   );
   gpc1_1 gpc2693 (
      {stage0_3[500]},
      {stage1_3[310]}
   );
   gpc1_1 gpc2694 (
      {stage0_3[501]},
      {stage1_3[311]}
   );
   gpc1_1 gpc2695 (
      {stage0_3[502]},
      {stage1_3[312]}
   );
   gpc1_1 gpc2696 (
      {stage0_3[503]},
      {stage1_3[313]}
   );
   gpc1_1 gpc2697 (
      {stage0_3[504]},
      {stage1_3[314]}
   );
   gpc1_1 gpc2698 (
      {stage0_3[505]},
      {stage1_3[315]}
   );
   gpc1_1 gpc2699 (
      {stage0_3[506]},
      {stage1_3[316]}
   );
   gpc1_1 gpc2700 (
      {stage0_3[507]},
      {stage1_3[317]}
   );
   gpc1_1 gpc2701 (
      {stage0_3[508]},
      {stage1_3[318]}
   );
   gpc1_1 gpc2702 (
      {stage0_3[509]},
      {stage1_3[319]}
   );
   gpc1_1 gpc2703 (
      {stage0_3[510]},
      {stage1_3[320]}
   );
   gpc1_1 gpc2704 (
      {stage0_3[511]},
      {stage1_3[321]}
   );
   gpc1_1 gpc2705 (
      {stage0_5[468]},
      {stage1_5[173]}
   );
   gpc1_1 gpc2706 (
      {stage0_5[469]},
      {stage1_5[174]}
   );
   gpc1_1 gpc2707 (
      {stage0_5[470]},
      {stage1_5[175]}
   );
   gpc1_1 gpc2708 (
      {stage0_5[471]},
      {stage1_5[176]}
   );
   gpc1_1 gpc2709 (
      {stage0_5[472]},
      {stage1_5[177]}
   );
   gpc1_1 gpc2710 (
      {stage0_5[473]},
      {stage1_5[178]}
   );
   gpc1_1 gpc2711 (
      {stage0_5[474]},
      {stage1_5[179]}
   );
   gpc1_1 gpc2712 (
      {stage0_5[475]},
      {stage1_5[180]}
   );
   gpc1_1 gpc2713 (
      {stage0_5[476]},
      {stage1_5[181]}
   );
   gpc1_1 gpc2714 (
      {stage0_5[477]},
      {stage1_5[182]}
   );
   gpc1_1 gpc2715 (
      {stage0_5[478]},
      {stage1_5[183]}
   );
   gpc1_1 gpc2716 (
      {stage0_5[479]},
      {stage1_5[184]}
   );
   gpc1_1 gpc2717 (
      {stage0_5[480]},
      {stage1_5[185]}
   );
   gpc1_1 gpc2718 (
      {stage0_5[481]},
      {stage1_5[186]}
   );
   gpc1_1 gpc2719 (
      {stage0_5[482]},
      {stage1_5[187]}
   );
   gpc1_1 gpc2720 (
      {stage0_5[483]},
      {stage1_5[188]}
   );
   gpc1_1 gpc2721 (
      {stage0_5[484]},
      {stage1_5[189]}
   );
   gpc1_1 gpc2722 (
      {stage0_5[485]},
      {stage1_5[190]}
   );
   gpc1_1 gpc2723 (
      {stage0_5[486]},
      {stage1_5[191]}
   );
   gpc1_1 gpc2724 (
      {stage0_5[487]},
      {stage1_5[192]}
   );
   gpc1_1 gpc2725 (
      {stage0_5[488]},
      {stage1_5[193]}
   );
   gpc1_1 gpc2726 (
      {stage0_5[489]},
      {stage1_5[194]}
   );
   gpc1_1 gpc2727 (
      {stage0_5[490]},
      {stage1_5[195]}
   );
   gpc1_1 gpc2728 (
      {stage0_5[491]},
      {stage1_5[196]}
   );
   gpc1_1 gpc2729 (
      {stage0_5[492]},
      {stage1_5[197]}
   );
   gpc1_1 gpc2730 (
      {stage0_5[493]},
      {stage1_5[198]}
   );
   gpc1_1 gpc2731 (
      {stage0_5[494]},
      {stage1_5[199]}
   );
   gpc1_1 gpc2732 (
      {stage0_5[495]},
      {stage1_5[200]}
   );
   gpc1_1 gpc2733 (
      {stage0_5[496]},
      {stage1_5[201]}
   );
   gpc1_1 gpc2734 (
      {stage0_5[497]},
      {stage1_5[202]}
   );
   gpc1_1 gpc2735 (
      {stage0_5[498]},
      {stage1_5[203]}
   );
   gpc1_1 gpc2736 (
      {stage0_5[499]},
      {stage1_5[204]}
   );
   gpc1_1 gpc2737 (
      {stage0_5[500]},
      {stage1_5[205]}
   );
   gpc1_1 gpc2738 (
      {stage0_5[501]},
      {stage1_5[206]}
   );
   gpc1_1 gpc2739 (
      {stage0_5[502]},
      {stage1_5[207]}
   );
   gpc1_1 gpc2740 (
      {stage0_5[503]},
      {stage1_5[208]}
   );
   gpc1_1 gpc2741 (
      {stage0_5[504]},
      {stage1_5[209]}
   );
   gpc1_1 gpc2742 (
      {stage0_5[505]},
      {stage1_5[210]}
   );
   gpc1_1 gpc2743 (
      {stage0_5[506]},
      {stage1_5[211]}
   );
   gpc1_1 gpc2744 (
      {stage0_5[507]},
      {stage1_5[212]}
   );
   gpc1_1 gpc2745 (
      {stage0_5[508]},
      {stage1_5[213]}
   );
   gpc1_1 gpc2746 (
      {stage0_5[509]},
      {stage1_5[214]}
   );
   gpc1_1 gpc2747 (
      {stage0_5[510]},
      {stage1_5[215]}
   );
   gpc1_1 gpc2748 (
      {stage0_5[511]},
      {stage1_5[216]}
   );
   gpc1_1 gpc2749 (
      {stage0_6[493]},
      {stage1_6[161]}
   );
   gpc1_1 gpc2750 (
      {stage0_6[494]},
      {stage1_6[162]}
   );
   gpc1_1 gpc2751 (
      {stage0_6[495]},
      {stage1_6[163]}
   );
   gpc1_1 gpc2752 (
      {stage0_6[496]},
      {stage1_6[164]}
   );
   gpc1_1 gpc2753 (
      {stage0_6[497]},
      {stage1_6[165]}
   );
   gpc1_1 gpc2754 (
      {stage0_6[498]},
      {stage1_6[166]}
   );
   gpc1_1 gpc2755 (
      {stage0_6[499]},
      {stage1_6[167]}
   );
   gpc1_1 gpc2756 (
      {stage0_6[500]},
      {stage1_6[168]}
   );
   gpc1_1 gpc2757 (
      {stage0_6[501]},
      {stage1_6[169]}
   );
   gpc1_1 gpc2758 (
      {stage0_6[502]},
      {stage1_6[170]}
   );
   gpc1_1 gpc2759 (
      {stage0_6[503]},
      {stage1_6[171]}
   );
   gpc1_1 gpc2760 (
      {stage0_6[504]},
      {stage1_6[172]}
   );
   gpc1_1 gpc2761 (
      {stage0_6[505]},
      {stage1_6[173]}
   );
   gpc1_1 gpc2762 (
      {stage0_6[506]},
      {stage1_6[174]}
   );
   gpc1_1 gpc2763 (
      {stage0_6[507]},
      {stage1_6[175]}
   );
   gpc1_1 gpc2764 (
      {stage0_6[508]},
      {stage1_6[176]}
   );
   gpc1_1 gpc2765 (
      {stage0_6[509]},
      {stage1_6[177]}
   );
   gpc1_1 gpc2766 (
      {stage0_6[510]},
      {stage1_6[178]}
   );
   gpc1_1 gpc2767 (
      {stage0_6[511]},
      {stage1_6[179]}
   );
   gpc1_1 gpc2768 (
      {stage0_7[364]},
      {stage1_7[192]}
   );
   gpc1_1 gpc2769 (
      {stage0_7[365]},
      {stage1_7[193]}
   );
   gpc1_1 gpc2770 (
      {stage0_7[366]},
      {stage1_7[194]}
   );
   gpc1_1 gpc2771 (
      {stage0_7[367]},
      {stage1_7[195]}
   );
   gpc1_1 gpc2772 (
      {stage0_7[368]},
      {stage1_7[196]}
   );
   gpc1_1 gpc2773 (
      {stage0_7[369]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2774 (
      {stage0_7[370]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2775 (
      {stage0_7[371]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2776 (
      {stage0_7[372]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2777 (
      {stage0_7[373]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2778 (
      {stage0_7[374]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2779 (
      {stage0_7[375]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2780 (
      {stage0_7[376]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2781 (
      {stage0_7[377]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2782 (
      {stage0_7[378]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2783 (
      {stage0_7[379]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2784 (
      {stage0_7[380]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2785 (
      {stage0_7[381]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2786 (
      {stage0_7[382]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2787 (
      {stage0_7[383]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2788 (
      {stage0_7[384]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2789 (
      {stage0_7[385]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2790 (
      {stage0_7[386]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2791 (
      {stage0_7[387]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2792 (
      {stage0_7[388]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2793 (
      {stage0_7[389]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2794 (
      {stage0_7[390]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2795 (
      {stage0_7[391]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2796 (
      {stage0_7[392]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2797 (
      {stage0_7[393]},
      {stage1_7[221]}
   );
   gpc1_1 gpc2798 (
      {stage0_7[394]},
      {stage1_7[222]}
   );
   gpc1_1 gpc2799 (
      {stage0_7[395]},
      {stage1_7[223]}
   );
   gpc1_1 gpc2800 (
      {stage0_7[396]},
      {stage1_7[224]}
   );
   gpc1_1 gpc2801 (
      {stage0_7[397]},
      {stage1_7[225]}
   );
   gpc1_1 gpc2802 (
      {stage0_7[398]},
      {stage1_7[226]}
   );
   gpc1_1 gpc2803 (
      {stage0_7[399]},
      {stage1_7[227]}
   );
   gpc1_1 gpc2804 (
      {stage0_7[400]},
      {stage1_7[228]}
   );
   gpc1_1 gpc2805 (
      {stage0_7[401]},
      {stage1_7[229]}
   );
   gpc1_1 gpc2806 (
      {stage0_7[402]},
      {stage1_7[230]}
   );
   gpc1_1 gpc2807 (
      {stage0_7[403]},
      {stage1_7[231]}
   );
   gpc1_1 gpc2808 (
      {stage0_7[404]},
      {stage1_7[232]}
   );
   gpc1_1 gpc2809 (
      {stage0_7[405]},
      {stage1_7[233]}
   );
   gpc1_1 gpc2810 (
      {stage0_7[406]},
      {stage1_7[234]}
   );
   gpc1_1 gpc2811 (
      {stage0_7[407]},
      {stage1_7[235]}
   );
   gpc1_1 gpc2812 (
      {stage0_7[408]},
      {stage1_7[236]}
   );
   gpc1_1 gpc2813 (
      {stage0_7[409]},
      {stage1_7[237]}
   );
   gpc1_1 gpc2814 (
      {stage0_7[410]},
      {stage1_7[238]}
   );
   gpc1_1 gpc2815 (
      {stage0_7[411]},
      {stage1_7[239]}
   );
   gpc1_1 gpc2816 (
      {stage0_7[412]},
      {stage1_7[240]}
   );
   gpc1_1 gpc2817 (
      {stage0_7[413]},
      {stage1_7[241]}
   );
   gpc1_1 gpc2818 (
      {stage0_7[414]},
      {stage1_7[242]}
   );
   gpc1_1 gpc2819 (
      {stage0_7[415]},
      {stage1_7[243]}
   );
   gpc1_1 gpc2820 (
      {stage0_7[416]},
      {stage1_7[244]}
   );
   gpc1_1 gpc2821 (
      {stage0_7[417]},
      {stage1_7[245]}
   );
   gpc1_1 gpc2822 (
      {stage0_7[418]},
      {stage1_7[246]}
   );
   gpc1_1 gpc2823 (
      {stage0_7[419]},
      {stage1_7[247]}
   );
   gpc1_1 gpc2824 (
      {stage0_7[420]},
      {stage1_7[248]}
   );
   gpc1_1 gpc2825 (
      {stage0_7[421]},
      {stage1_7[249]}
   );
   gpc1_1 gpc2826 (
      {stage0_7[422]},
      {stage1_7[250]}
   );
   gpc1_1 gpc2827 (
      {stage0_7[423]},
      {stage1_7[251]}
   );
   gpc1_1 gpc2828 (
      {stage0_7[424]},
      {stage1_7[252]}
   );
   gpc1_1 gpc2829 (
      {stage0_7[425]},
      {stage1_7[253]}
   );
   gpc1_1 gpc2830 (
      {stage0_7[426]},
      {stage1_7[254]}
   );
   gpc1_1 gpc2831 (
      {stage0_7[427]},
      {stage1_7[255]}
   );
   gpc1_1 gpc2832 (
      {stage0_7[428]},
      {stage1_7[256]}
   );
   gpc1_1 gpc2833 (
      {stage0_7[429]},
      {stage1_7[257]}
   );
   gpc1_1 gpc2834 (
      {stage0_7[430]},
      {stage1_7[258]}
   );
   gpc1_1 gpc2835 (
      {stage0_7[431]},
      {stage1_7[259]}
   );
   gpc1_1 gpc2836 (
      {stage0_7[432]},
      {stage1_7[260]}
   );
   gpc1_1 gpc2837 (
      {stage0_7[433]},
      {stage1_7[261]}
   );
   gpc1_1 gpc2838 (
      {stage0_7[434]},
      {stage1_7[262]}
   );
   gpc1_1 gpc2839 (
      {stage0_7[435]},
      {stage1_7[263]}
   );
   gpc1_1 gpc2840 (
      {stage0_7[436]},
      {stage1_7[264]}
   );
   gpc1_1 gpc2841 (
      {stage0_7[437]},
      {stage1_7[265]}
   );
   gpc1_1 gpc2842 (
      {stage0_7[438]},
      {stage1_7[266]}
   );
   gpc1_1 gpc2843 (
      {stage0_7[439]},
      {stage1_7[267]}
   );
   gpc1_1 gpc2844 (
      {stage0_7[440]},
      {stage1_7[268]}
   );
   gpc1_1 gpc2845 (
      {stage0_7[441]},
      {stage1_7[269]}
   );
   gpc1_1 gpc2846 (
      {stage0_7[442]},
      {stage1_7[270]}
   );
   gpc1_1 gpc2847 (
      {stage0_7[443]},
      {stage1_7[271]}
   );
   gpc1_1 gpc2848 (
      {stage0_7[444]},
      {stage1_7[272]}
   );
   gpc1_1 gpc2849 (
      {stage0_7[445]},
      {stage1_7[273]}
   );
   gpc1_1 gpc2850 (
      {stage0_7[446]},
      {stage1_7[274]}
   );
   gpc1_1 gpc2851 (
      {stage0_7[447]},
      {stage1_7[275]}
   );
   gpc1_1 gpc2852 (
      {stage0_7[448]},
      {stage1_7[276]}
   );
   gpc1_1 gpc2853 (
      {stage0_7[449]},
      {stage1_7[277]}
   );
   gpc1_1 gpc2854 (
      {stage0_7[450]},
      {stage1_7[278]}
   );
   gpc1_1 gpc2855 (
      {stage0_7[451]},
      {stage1_7[279]}
   );
   gpc1_1 gpc2856 (
      {stage0_7[452]},
      {stage1_7[280]}
   );
   gpc1_1 gpc2857 (
      {stage0_7[453]},
      {stage1_7[281]}
   );
   gpc1_1 gpc2858 (
      {stage0_7[454]},
      {stage1_7[282]}
   );
   gpc1_1 gpc2859 (
      {stage0_7[455]},
      {stage1_7[283]}
   );
   gpc1_1 gpc2860 (
      {stage0_7[456]},
      {stage1_7[284]}
   );
   gpc1_1 gpc2861 (
      {stage0_7[457]},
      {stage1_7[285]}
   );
   gpc1_1 gpc2862 (
      {stage0_7[458]},
      {stage1_7[286]}
   );
   gpc1_1 gpc2863 (
      {stage0_7[459]},
      {stage1_7[287]}
   );
   gpc1_1 gpc2864 (
      {stage0_7[460]},
      {stage1_7[288]}
   );
   gpc1_1 gpc2865 (
      {stage0_7[461]},
      {stage1_7[289]}
   );
   gpc1_1 gpc2866 (
      {stage0_7[462]},
      {stage1_7[290]}
   );
   gpc1_1 gpc2867 (
      {stage0_7[463]},
      {stage1_7[291]}
   );
   gpc1_1 gpc2868 (
      {stage0_7[464]},
      {stage1_7[292]}
   );
   gpc1_1 gpc2869 (
      {stage0_7[465]},
      {stage1_7[293]}
   );
   gpc1_1 gpc2870 (
      {stage0_7[466]},
      {stage1_7[294]}
   );
   gpc1_1 gpc2871 (
      {stage0_7[467]},
      {stage1_7[295]}
   );
   gpc1_1 gpc2872 (
      {stage0_7[468]},
      {stage1_7[296]}
   );
   gpc1_1 gpc2873 (
      {stage0_7[469]},
      {stage1_7[297]}
   );
   gpc1_1 gpc2874 (
      {stage0_7[470]},
      {stage1_7[298]}
   );
   gpc1_1 gpc2875 (
      {stage0_7[471]},
      {stage1_7[299]}
   );
   gpc1_1 gpc2876 (
      {stage0_7[472]},
      {stage1_7[300]}
   );
   gpc1_1 gpc2877 (
      {stage0_7[473]},
      {stage1_7[301]}
   );
   gpc1_1 gpc2878 (
      {stage0_7[474]},
      {stage1_7[302]}
   );
   gpc1_1 gpc2879 (
      {stage0_7[475]},
      {stage1_7[303]}
   );
   gpc1_1 gpc2880 (
      {stage0_7[476]},
      {stage1_7[304]}
   );
   gpc1_1 gpc2881 (
      {stage0_7[477]},
      {stage1_7[305]}
   );
   gpc1_1 gpc2882 (
      {stage0_7[478]},
      {stage1_7[306]}
   );
   gpc1_1 gpc2883 (
      {stage0_7[479]},
      {stage1_7[307]}
   );
   gpc1_1 gpc2884 (
      {stage0_7[480]},
      {stage1_7[308]}
   );
   gpc1_1 gpc2885 (
      {stage0_7[481]},
      {stage1_7[309]}
   );
   gpc1_1 gpc2886 (
      {stage0_7[482]},
      {stage1_7[310]}
   );
   gpc1_1 gpc2887 (
      {stage0_7[483]},
      {stage1_7[311]}
   );
   gpc1_1 gpc2888 (
      {stage0_7[484]},
      {stage1_7[312]}
   );
   gpc1_1 gpc2889 (
      {stage0_7[485]},
      {stage1_7[313]}
   );
   gpc1_1 gpc2890 (
      {stage0_7[486]},
      {stage1_7[314]}
   );
   gpc1_1 gpc2891 (
      {stage0_7[487]},
      {stage1_7[315]}
   );
   gpc1_1 gpc2892 (
      {stage0_7[488]},
      {stage1_7[316]}
   );
   gpc1_1 gpc2893 (
      {stage0_7[489]},
      {stage1_7[317]}
   );
   gpc1_1 gpc2894 (
      {stage0_7[490]},
      {stage1_7[318]}
   );
   gpc1_1 gpc2895 (
      {stage0_7[491]},
      {stage1_7[319]}
   );
   gpc1_1 gpc2896 (
      {stage0_7[492]},
      {stage1_7[320]}
   );
   gpc1_1 gpc2897 (
      {stage0_7[493]},
      {stage1_7[321]}
   );
   gpc1_1 gpc2898 (
      {stage0_7[494]},
      {stage1_7[322]}
   );
   gpc1_1 gpc2899 (
      {stage0_7[495]},
      {stage1_7[323]}
   );
   gpc1_1 gpc2900 (
      {stage0_7[496]},
      {stage1_7[324]}
   );
   gpc1_1 gpc2901 (
      {stage0_7[497]},
      {stage1_7[325]}
   );
   gpc1_1 gpc2902 (
      {stage0_7[498]},
      {stage1_7[326]}
   );
   gpc1_1 gpc2903 (
      {stage0_7[499]},
      {stage1_7[327]}
   );
   gpc1_1 gpc2904 (
      {stage0_7[500]},
      {stage1_7[328]}
   );
   gpc1_1 gpc2905 (
      {stage0_7[501]},
      {stage1_7[329]}
   );
   gpc1_1 gpc2906 (
      {stage0_7[502]},
      {stage1_7[330]}
   );
   gpc1_1 gpc2907 (
      {stage0_7[503]},
      {stage1_7[331]}
   );
   gpc1_1 gpc2908 (
      {stage0_7[504]},
      {stage1_7[332]}
   );
   gpc1_1 gpc2909 (
      {stage0_7[505]},
      {stage1_7[333]}
   );
   gpc1_1 gpc2910 (
      {stage0_7[506]},
      {stage1_7[334]}
   );
   gpc1_1 gpc2911 (
      {stage0_7[507]},
      {stage1_7[335]}
   );
   gpc1_1 gpc2912 (
      {stage0_7[508]},
      {stage1_7[336]}
   );
   gpc1_1 gpc2913 (
      {stage0_7[509]},
      {stage1_7[337]}
   );
   gpc1_1 gpc2914 (
      {stage0_7[510]},
      {stage1_7[338]}
   );
   gpc1_1 gpc2915 (
      {stage0_7[511]},
      {stage1_7[339]}
   );
   gpc1_1 gpc2916 (
      {stage0_8[493]},
      {stage1_8[220]}
   );
   gpc1_1 gpc2917 (
      {stage0_8[494]},
      {stage1_8[221]}
   );
   gpc1_1 gpc2918 (
      {stage0_8[495]},
      {stage1_8[222]}
   );
   gpc1_1 gpc2919 (
      {stage0_8[496]},
      {stage1_8[223]}
   );
   gpc1_1 gpc2920 (
      {stage0_8[497]},
      {stage1_8[224]}
   );
   gpc1_1 gpc2921 (
      {stage0_8[498]},
      {stage1_8[225]}
   );
   gpc1_1 gpc2922 (
      {stage0_8[499]},
      {stage1_8[226]}
   );
   gpc1_1 gpc2923 (
      {stage0_8[500]},
      {stage1_8[227]}
   );
   gpc1_1 gpc2924 (
      {stage0_8[501]},
      {stage1_8[228]}
   );
   gpc1_1 gpc2925 (
      {stage0_8[502]},
      {stage1_8[229]}
   );
   gpc1_1 gpc2926 (
      {stage0_8[503]},
      {stage1_8[230]}
   );
   gpc1_1 gpc2927 (
      {stage0_8[504]},
      {stage1_8[231]}
   );
   gpc1_1 gpc2928 (
      {stage0_8[505]},
      {stage1_8[232]}
   );
   gpc1_1 gpc2929 (
      {stage0_8[506]},
      {stage1_8[233]}
   );
   gpc1_1 gpc2930 (
      {stage0_8[507]},
      {stage1_8[234]}
   );
   gpc1_1 gpc2931 (
      {stage0_8[508]},
      {stage1_8[235]}
   );
   gpc1_1 gpc2932 (
      {stage0_8[509]},
      {stage1_8[236]}
   );
   gpc1_1 gpc2933 (
      {stage0_8[510]},
      {stage1_8[237]}
   );
   gpc1_1 gpc2934 (
      {stage0_8[511]},
      {stage1_8[238]}
   );
   gpc1_1 gpc2935 (
      {stage0_9[312]},
      {stage1_9[163]}
   );
   gpc1_1 gpc2936 (
      {stage0_9[313]},
      {stage1_9[164]}
   );
   gpc1_1 gpc2937 (
      {stage0_9[314]},
      {stage1_9[165]}
   );
   gpc1_1 gpc2938 (
      {stage0_9[315]},
      {stage1_9[166]}
   );
   gpc1_1 gpc2939 (
      {stage0_9[316]},
      {stage1_9[167]}
   );
   gpc1_1 gpc2940 (
      {stage0_9[317]},
      {stage1_9[168]}
   );
   gpc1_1 gpc2941 (
      {stage0_9[318]},
      {stage1_9[169]}
   );
   gpc1_1 gpc2942 (
      {stage0_9[319]},
      {stage1_9[170]}
   );
   gpc1_1 gpc2943 (
      {stage0_9[320]},
      {stage1_9[171]}
   );
   gpc1_1 gpc2944 (
      {stage0_9[321]},
      {stage1_9[172]}
   );
   gpc1_1 gpc2945 (
      {stage0_9[322]},
      {stage1_9[173]}
   );
   gpc1_1 gpc2946 (
      {stage0_9[323]},
      {stage1_9[174]}
   );
   gpc1_1 gpc2947 (
      {stage0_9[324]},
      {stage1_9[175]}
   );
   gpc1_1 gpc2948 (
      {stage0_9[325]},
      {stage1_9[176]}
   );
   gpc1_1 gpc2949 (
      {stage0_9[326]},
      {stage1_9[177]}
   );
   gpc1_1 gpc2950 (
      {stage0_9[327]},
      {stage1_9[178]}
   );
   gpc1_1 gpc2951 (
      {stage0_9[328]},
      {stage1_9[179]}
   );
   gpc1_1 gpc2952 (
      {stage0_9[329]},
      {stage1_9[180]}
   );
   gpc1_1 gpc2953 (
      {stage0_9[330]},
      {stage1_9[181]}
   );
   gpc1_1 gpc2954 (
      {stage0_9[331]},
      {stage1_9[182]}
   );
   gpc1_1 gpc2955 (
      {stage0_9[332]},
      {stage1_9[183]}
   );
   gpc1_1 gpc2956 (
      {stage0_9[333]},
      {stage1_9[184]}
   );
   gpc1_1 gpc2957 (
      {stage0_9[334]},
      {stage1_9[185]}
   );
   gpc1_1 gpc2958 (
      {stage0_9[335]},
      {stage1_9[186]}
   );
   gpc1_1 gpc2959 (
      {stage0_9[336]},
      {stage1_9[187]}
   );
   gpc1_1 gpc2960 (
      {stage0_9[337]},
      {stage1_9[188]}
   );
   gpc1_1 gpc2961 (
      {stage0_9[338]},
      {stage1_9[189]}
   );
   gpc1_1 gpc2962 (
      {stage0_9[339]},
      {stage1_9[190]}
   );
   gpc1_1 gpc2963 (
      {stage0_9[340]},
      {stage1_9[191]}
   );
   gpc1_1 gpc2964 (
      {stage0_9[341]},
      {stage1_9[192]}
   );
   gpc1_1 gpc2965 (
      {stage0_9[342]},
      {stage1_9[193]}
   );
   gpc1_1 gpc2966 (
      {stage0_9[343]},
      {stage1_9[194]}
   );
   gpc1_1 gpc2967 (
      {stage0_9[344]},
      {stage1_9[195]}
   );
   gpc1_1 gpc2968 (
      {stage0_9[345]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2969 (
      {stage0_9[346]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2970 (
      {stage0_9[347]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2971 (
      {stage0_9[348]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2972 (
      {stage0_9[349]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2973 (
      {stage0_9[350]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2974 (
      {stage0_9[351]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2975 (
      {stage0_9[352]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2976 (
      {stage0_9[353]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2977 (
      {stage0_9[354]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2978 (
      {stage0_9[355]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2979 (
      {stage0_9[356]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2980 (
      {stage0_9[357]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2981 (
      {stage0_9[358]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2982 (
      {stage0_9[359]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2983 (
      {stage0_9[360]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2984 (
      {stage0_9[361]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2985 (
      {stage0_9[362]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2986 (
      {stage0_9[363]},
      {stage1_9[214]}
   );
   gpc1_1 gpc2987 (
      {stage0_9[364]},
      {stage1_9[215]}
   );
   gpc1_1 gpc2988 (
      {stage0_9[365]},
      {stage1_9[216]}
   );
   gpc1_1 gpc2989 (
      {stage0_9[366]},
      {stage1_9[217]}
   );
   gpc1_1 gpc2990 (
      {stage0_9[367]},
      {stage1_9[218]}
   );
   gpc1_1 gpc2991 (
      {stage0_9[368]},
      {stage1_9[219]}
   );
   gpc1_1 gpc2992 (
      {stage0_9[369]},
      {stage1_9[220]}
   );
   gpc1_1 gpc2993 (
      {stage0_9[370]},
      {stage1_9[221]}
   );
   gpc1_1 gpc2994 (
      {stage0_9[371]},
      {stage1_9[222]}
   );
   gpc1_1 gpc2995 (
      {stage0_9[372]},
      {stage1_9[223]}
   );
   gpc1_1 gpc2996 (
      {stage0_9[373]},
      {stage1_9[224]}
   );
   gpc1_1 gpc2997 (
      {stage0_9[374]},
      {stage1_9[225]}
   );
   gpc1_1 gpc2998 (
      {stage0_9[375]},
      {stage1_9[226]}
   );
   gpc1_1 gpc2999 (
      {stage0_9[376]},
      {stage1_9[227]}
   );
   gpc1_1 gpc3000 (
      {stage0_9[377]},
      {stage1_9[228]}
   );
   gpc1_1 gpc3001 (
      {stage0_9[378]},
      {stage1_9[229]}
   );
   gpc1_1 gpc3002 (
      {stage0_9[379]},
      {stage1_9[230]}
   );
   gpc1_1 gpc3003 (
      {stage0_9[380]},
      {stage1_9[231]}
   );
   gpc1_1 gpc3004 (
      {stage0_9[381]},
      {stage1_9[232]}
   );
   gpc1_1 gpc3005 (
      {stage0_9[382]},
      {stage1_9[233]}
   );
   gpc1_1 gpc3006 (
      {stage0_9[383]},
      {stage1_9[234]}
   );
   gpc1_1 gpc3007 (
      {stage0_9[384]},
      {stage1_9[235]}
   );
   gpc1_1 gpc3008 (
      {stage0_9[385]},
      {stage1_9[236]}
   );
   gpc1_1 gpc3009 (
      {stage0_9[386]},
      {stage1_9[237]}
   );
   gpc1_1 gpc3010 (
      {stage0_9[387]},
      {stage1_9[238]}
   );
   gpc1_1 gpc3011 (
      {stage0_9[388]},
      {stage1_9[239]}
   );
   gpc1_1 gpc3012 (
      {stage0_9[389]},
      {stage1_9[240]}
   );
   gpc1_1 gpc3013 (
      {stage0_9[390]},
      {stage1_9[241]}
   );
   gpc1_1 gpc3014 (
      {stage0_9[391]},
      {stage1_9[242]}
   );
   gpc1_1 gpc3015 (
      {stage0_9[392]},
      {stage1_9[243]}
   );
   gpc1_1 gpc3016 (
      {stage0_9[393]},
      {stage1_9[244]}
   );
   gpc1_1 gpc3017 (
      {stage0_9[394]},
      {stage1_9[245]}
   );
   gpc1_1 gpc3018 (
      {stage0_9[395]},
      {stage1_9[246]}
   );
   gpc1_1 gpc3019 (
      {stage0_9[396]},
      {stage1_9[247]}
   );
   gpc1_1 gpc3020 (
      {stage0_9[397]},
      {stage1_9[248]}
   );
   gpc1_1 gpc3021 (
      {stage0_9[398]},
      {stage1_9[249]}
   );
   gpc1_1 gpc3022 (
      {stage0_9[399]},
      {stage1_9[250]}
   );
   gpc1_1 gpc3023 (
      {stage0_9[400]},
      {stage1_9[251]}
   );
   gpc1_1 gpc3024 (
      {stage0_9[401]},
      {stage1_9[252]}
   );
   gpc1_1 gpc3025 (
      {stage0_9[402]},
      {stage1_9[253]}
   );
   gpc1_1 gpc3026 (
      {stage0_9[403]},
      {stage1_9[254]}
   );
   gpc1_1 gpc3027 (
      {stage0_9[404]},
      {stage1_9[255]}
   );
   gpc1_1 gpc3028 (
      {stage0_9[405]},
      {stage1_9[256]}
   );
   gpc1_1 gpc3029 (
      {stage0_9[406]},
      {stage1_9[257]}
   );
   gpc1_1 gpc3030 (
      {stage0_9[407]},
      {stage1_9[258]}
   );
   gpc1_1 gpc3031 (
      {stage0_9[408]},
      {stage1_9[259]}
   );
   gpc1_1 gpc3032 (
      {stage0_9[409]},
      {stage1_9[260]}
   );
   gpc1_1 gpc3033 (
      {stage0_9[410]},
      {stage1_9[261]}
   );
   gpc1_1 gpc3034 (
      {stage0_9[411]},
      {stage1_9[262]}
   );
   gpc1_1 gpc3035 (
      {stage0_9[412]},
      {stage1_9[263]}
   );
   gpc1_1 gpc3036 (
      {stage0_9[413]},
      {stage1_9[264]}
   );
   gpc1_1 gpc3037 (
      {stage0_9[414]},
      {stage1_9[265]}
   );
   gpc1_1 gpc3038 (
      {stage0_9[415]},
      {stage1_9[266]}
   );
   gpc1_1 gpc3039 (
      {stage0_9[416]},
      {stage1_9[267]}
   );
   gpc1_1 gpc3040 (
      {stage0_9[417]},
      {stage1_9[268]}
   );
   gpc1_1 gpc3041 (
      {stage0_9[418]},
      {stage1_9[269]}
   );
   gpc1_1 gpc3042 (
      {stage0_9[419]},
      {stage1_9[270]}
   );
   gpc1_1 gpc3043 (
      {stage0_9[420]},
      {stage1_9[271]}
   );
   gpc1_1 gpc3044 (
      {stage0_9[421]},
      {stage1_9[272]}
   );
   gpc1_1 gpc3045 (
      {stage0_9[422]},
      {stage1_9[273]}
   );
   gpc1_1 gpc3046 (
      {stage0_9[423]},
      {stage1_9[274]}
   );
   gpc1_1 gpc3047 (
      {stage0_9[424]},
      {stage1_9[275]}
   );
   gpc1_1 gpc3048 (
      {stage0_9[425]},
      {stage1_9[276]}
   );
   gpc1_1 gpc3049 (
      {stage0_9[426]},
      {stage1_9[277]}
   );
   gpc1_1 gpc3050 (
      {stage0_9[427]},
      {stage1_9[278]}
   );
   gpc1_1 gpc3051 (
      {stage0_9[428]},
      {stage1_9[279]}
   );
   gpc1_1 gpc3052 (
      {stage0_9[429]},
      {stage1_9[280]}
   );
   gpc1_1 gpc3053 (
      {stage0_9[430]},
      {stage1_9[281]}
   );
   gpc1_1 gpc3054 (
      {stage0_9[431]},
      {stage1_9[282]}
   );
   gpc1_1 gpc3055 (
      {stage0_9[432]},
      {stage1_9[283]}
   );
   gpc1_1 gpc3056 (
      {stage0_9[433]},
      {stage1_9[284]}
   );
   gpc1_1 gpc3057 (
      {stage0_9[434]},
      {stage1_9[285]}
   );
   gpc1_1 gpc3058 (
      {stage0_9[435]},
      {stage1_9[286]}
   );
   gpc1_1 gpc3059 (
      {stage0_9[436]},
      {stage1_9[287]}
   );
   gpc1_1 gpc3060 (
      {stage0_9[437]},
      {stage1_9[288]}
   );
   gpc1_1 gpc3061 (
      {stage0_9[438]},
      {stage1_9[289]}
   );
   gpc1_1 gpc3062 (
      {stage0_9[439]},
      {stage1_9[290]}
   );
   gpc1_1 gpc3063 (
      {stage0_9[440]},
      {stage1_9[291]}
   );
   gpc1_1 gpc3064 (
      {stage0_9[441]},
      {stage1_9[292]}
   );
   gpc1_1 gpc3065 (
      {stage0_9[442]},
      {stage1_9[293]}
   );
   gpc1_1 gpc3066 (
      {stage0_9[443]},
      {stage1_9[294]}
   );
   gpc1_1 gpc3067 (
      {stage0_9[444]},
      {stage1_9[295]}
   );
   gpc1_1 gpc3068 (
      {stage0_9[445]},
      {stage1_9[296]}
   );
   gpc1_1 gpc3069 (
      {stage0_9[446]},
      {stage1_9[297]}
   );
   gpc1_1 gpc3070 (
      {stage0_9[447]},
      {stage1_9[298]}
   );
   gpc1_1 gpc3071 (
      {stage0_9[448]},
      {stage1_9[299]}
   );
   gpc1_1 gpc3072 (
      {stage0_9[449]},
      {stage1_9[300]}
   );
   gpc1_1 gpc3073 (
      {stage0_9[450]},
      {stage1_9[301]}
   );
   gpc1_1 gpc3074 (
      {stage0_9[451]},
      {stage1_9[302]}
   );
   gpc1_1 gpc3075 (
      {stage0_9[452]},
      {stage1_9[303]}
   );
   gpc1_1 gpc3076 (
      {stage0_9[453]},
      {stage1_9[304]}
   );
   gpc1_1 gpc3077 (
      {stage0_9[454]},
      {stage1_9[305]}
   );
   gpc1_1 gpc3078 (
      {stage0_9[455]},
      {stage1_9[306]}
   );
   gpc1_1 gpc3079 (
      {stage0_9[456]},
      {stage1_9[307]}
   );
   gpc1_1 gpc3080 (
      {stage0_9[457]},
      {stage1_9[308]}
   );
   gpc1_1 gpc3081 (
      {stage0_9[458]},
      {stage1_9[309]}
   );
   gpc1_1 gpc3082 (
      {stage0_9[459]},
      {stage1_9[310]}
   );
   gpc1_1 gpc3083 (
      {stage0_9[460]},
      {stage1_9[311]}
   );
   gpc1_1 gpc3084 (
      {stage0_9[461]},
      {stage1_9[312]}
   );
   gpc1_1 gpc3085 (
      {stage0_9[462]},
      {stage1_9[313]}
   );
   gpc1_1 gpc3086 (
      {stage0_9[463]},
      {stage1_9[314]}
   );
   gpc1_1 gpc3087 (
      {stage0_9[464]},
      {stage1_9[315]}
   );
   gpc1_1 gpc3088 (
      {stage0_9[465]},
      {stage1_9[316]}
   );
   gpc1_1 gpc3089 (
      {stage0_9[466]},
      {stage1_9[317]}
   );
   gpc1_1 gpc3090 (
      {stage0_9[467]},
      {stage1_9[318]}
   );
   gpc1_1 gpc3091 (
      {stage0_9[468]},
      {stage1_9[319]}
   );
   gpc1_1 gpc3092 (
      {stage0_9[469]},
      {stage1_9[320]}
   );
   gpc1_1 gpc3093 (
      {stage0_9[470]},
      {stage1_9[321]}
   );
   gpc1_1 gpc3094 (
      {stage0_9[471]},
      {stage1_9[322]}
   );
   gpc1_1 gpc3095 (
      {stage0_9[472]},
      {stage1_9[323]}
   );
   gpc1_1 gpc3096 (
      {stage0_9[473]},
      {stage1_9[324]}
   );
   gpc1_1 gpc3097 (
      {stage0_9[474]},
      {stage1_9[325]}
   );
   gpc1_1 gpc3098 (
      {stage0_9[475]},
      {stage1_9[326]}
   );
   gpc1_1 gpc3099 (
      {stage0_9[476]},
      {stage1_9[327]}
   );
   gpc1_1 gpc3100 (
      {stage0_9[477]},
      {stage1_9[328]}
   );
   gpc1_1 gpc3101 (
      {stage0_9[478]},
      {stage1_9[329]}
   );
   gpc1_1 gpc3102 (
      {stage0_9[479]},
      {stage1_9[330]}
   );
   gpc1_1 gpc3103 (
      {stage0_9[480]},
      {stage1_9[331]}
   );
   gpc1_1 gpc3104 (
      {stage0_9[481]},
      {stage1_9[332]}
   );
   gpc1_1 gpc3105 (
      {stage0_9[482]},
      {stage1_9[333]}
   );
   gpc1_1 gpc3106 (
      {stage0_9[483]},
      {stage1_9[334]}
   );
   gpc1_1 gpc3107 (
      {stage0_9[484]},
      {stage1_9[335]}
   );
   gpc1_1 gpc3108 (
      {stage0_9[485]},
      {stage1_9[336]}
   );
   gpc1_1 gpc3109 (
      {stage0_9[486]},
      {stage1_9[337]}
   );
   gpc1_1 gpc3110 (
      {stage0_9[487]},
      {stage1_9[338]}
   );
   gpc1_1 gpc3111 (
      {stage0_9[488]},
      {stage1_9[339]}
   );
   gpc1_1 gpc3112 (
      {stage0_9[489]},
      {stage1_9[340]}
   );
   gpc1_1 gpc3113 (
      {stage0_9[490]},
      {stage1_9[341]}
   );
   gpc1_1 gpc3114 (
      {stage0_9[491]},
      {stage1_9[342]}
   );
   gpc1_1 gpc3115 (
      {stage0_9[492]},
      {stage1_9[343]}
   );
   gpc1_1 gpc3116 (
      {stage0_9[493]},
      {stage1_9[344]}
   );
   gpc1_1 gpc3117 (
      {stage0_9[494]},
      {stage1_9[345]}
   );
   gpc1_1 gpc3118 (
      {stage0_9[495]},
      {stage1_9[346]}
   );
   gpc1_1 gpc3119 (
      {stage0_9[496]},
      {stage1_9[347]}
   );
   gpc1_1 gpc3120 (
      {stage0_9[497]},
      {stage1_9[348]}
   );
   gpc1_1 gpc3121 (
      {stage0_9[498]},
      {stage1_9[349]}
   );
   gpc1_1 gpc3122 (
      {stage0_9[499]},
      {stage1_9[350]}
   );
   gpc1_1 gpc3123 (
      {stage0_9[500]},
      {stage1_9[351]}
   );
   gpc1_1 gpc3124 (
      {stage0_9[501]},
      {stage1_9[352]}
   );
   gpc1_1 gpc3125 (
      {stage0_9[502]},
      {stage1_9[353]}
   );
   gpc1_1 gpc3126 (
      {stage0_9[503]},
      {stage1_9[354]}
   );
   gpc1_1 gpc3127 (
      {stage0_9[504]},
      {stage1_9[355]}
   );
   gpc1_1 gpc3128 (
      {stage0_9[505]},
      {stage1_9[356]}
   );
   gpc1_1 gpc3129 (
      {stage0_9[506]},
      {stage1_9[357]}
   );
   gpc1_1 gpc3130 (
      {stage0_9[507]},
      {stage1_9[358]}
   );
   gpc1_1 gpc3131 (
      {stage0_9[508]},
      {stage1_9[359]}
   );
   gpc1_1 gpc3132 (
      {stage0_9[509]},
      {stage1_9[360]}
   );
   gpc1_1 gpc3133 (
      {stage0_9[510]},
      {stage1_9[361]}
   );
   gpc1_1 gpc3134 (
      {stage0_9[511]},
      {stage1_9[362]}
   );
   gpc1_1 gpc3135 (
      {stage0_10[502]},
      {stage1_10[143]}
   );
   gpc1_1 gpc3136 (
      {stage0_10[503]},
      {stage1_10[144]}
   );
   gpc1_1 gpc3137 (
      {stage0_10[504]},
      {stage1_10[145]}
   );
   gpc1_1 gpc3138 (
      {stage0_10[505]},
      {stage1_10[146]}
   );
   gpc1_1 gpc3139 (
      {stage0_10[506]},
      {stage1_10[147]}
   );
   gpc1_1 gpc3140 (
      {stage0_10[507]},
      {stage1_10[148]}
   );
   gpc1_1 gpc3141 (
      {stage0_10[508]},
      {stage1_10[149]}
   );
   gpc1_1 gpc3142 (
      {stage0_10[509]},
      {stage1_10[150]}
   );
   gpc1_1 gpc3143 (
      {stage0_10[510]},
      {stage1_10[151]}
   );
   gpc1_1 gpc3144 (
      {stage0_10[511]},
      {stage1_10[152]}
   );
   gpc1_1 gpc3145 (
      {stage0_11[380]},
      {stage1_11[186]}
   );
   gpc1_1 gpc3146 (
      {stage0_11[381]},
      {stage1_11[187]}
   );
   gpc1_1 gpc3147 (
      {stage0_11[382]},
      {stage1_11[188]}
   );
   gpc1_1 gpc3148 (
      {stage0_11[383]},
      {stage1_11[189]}
   );
   gpc1_1 gpc3149 (
      {stage0_11[384]},
      {stage1_11[190]}
   );
   gpc1_1 gpc3150 (
      {stage0_11[385]},
      {stage1_11[191]}
   );
   gpc1_1 gpc3151 (
      {stage0_11[386]},
      {stage1_11[192]}
   );
   gpc1_1 gpc3152 (
      {stage0_11[387]},
      {stage1_11[193]}
   );
   gpc1_1 gpc3153 (
      {stage0_11[388]},
      {stage1_11[194]}
   );
   gpc1_1 gpc3154 (
      {stage0_11[389]},
      {stage1_11[195]}
   );
   gpc1_1 gpc3155 (
      {stage0_11[390]},
      {stage1_11[196]}
   );
   gpc1_1 gpc3156 (
      {stage0_11[391]},
      {stage1_11[197]}
   );
   gpc1_1 gpc3157 (
      {stage0_11[392]},
      {stage1_11[198]}
   );
   gpc1_1 gpc3158 (
      {stage0_11[393]},
      {stage1_11[199]}
   );
   gpc1_1 gpc3159 (
      {stage0_11[394]},
      {stage1_11[200]}
   );
   gpc1_1 gpc3160 (
      {stage0_11[395]},
      {stage1_11[201]}
   );
   gpc1_1 gpc3161 (
      {stage0_11[396]},
      {stage1_11[202]}
   );
   gpc1_1 gpc3162 (
      {stage0_11[397]},
      {stage1_11[203]}
   );
   gpc1_1 gpc3163 (
      {stage0_11[398]},
      {stage1_11[204]}
   );
   gpc1_1 gpc3164 (
      {stage0_11[399]},
      {stage1_11[205]}
   );
   gpc1_1 gpc3165 (
      {stage0_11[400]},
      {stage1_11[206]}
   );
   gpc1_1 gpc3166 (
      {stage0_11[401]},
      {stage1_11[207]}
   );
   gpc1_1 gpc3167 (
      {stage0_11[402]},
      {stage1_11[208]}
   );
   gpc1_1 gpc3168 (
      {stage0_11[403]},
      {stage1_11[209]}
   );
   gpc1_1 gpc3169 (
      {stage0_11[404]},
      {stage1_11[210]}
   );
   gpc1_1 gpc3170 (
      {stage0_11[405]},
      {stage1_11[211]}
   );
   gpc1_1 gpc3171 (
      {stage0_11[406]},
      {stage1_11[212]}
   );
   gpc1_1 gpc3172 (
      {stage0_11[407]},
      {stage1_11[213]}
   );
   gpc1_1 gpc3173 (
      {stage0_11[408]},
      {stage1_11[214]}
   );
   gpc1_1 gpc3174 (
      {stage0_11[409]},
      {stage1_11[215]}
   );
   gpc1_1 gpc3175 (
      {stage0_11[410]},
      {stage1_11[216]}
   );
   gpc1_1 gpc3176 (
      {stage0_11[411]},
      {stage1_11[217]}
   );
   gpc1_1 gpc3177 (
      {stage0_11[412]},
      {stage1_11[218]}
   );
   gpc1_1 gpc3178 (
      {stage0_11[413]},
      {stage1_11[219]}
   );
   gpc1_1 gpc3179 (
      {stage0_11[414]},
      {stage1_11[220]}
   );
   gpc1_1 gpc3180 (
      {stage0_11[415]},
      {stage1_11[221]}
   );
   gpc1_1 gpc3181 (
      {stage0_11[416]},
      {stage1_11[222]}
   );
   gpc1_1 gpc3182 (
      {stage0_11[417]},
      {stage1_11[223]}
   );
   gpc1_1 gpc3183 (
      {stage0_11[418]},
      {stage1_11[224]}
   );
   gpc1_1 gpc3184 (
      {stage0_11[419]},
      {stage1_11[225]}
   );
   gpc1_1 gpc3185 (
      {stage0_11[420]},
      {stage1_11[226]}
   );
   gpc1_1 gpc3186 (
      {stage0_11[421]},
      {stage1_11[227]}
   );
   gpc1_1 gpc3187 (
      {stage0_11[422]},
      {stage1_11[228]}
   );
   gpc1_1 gpc3188 (
      {stage0_11[423]},
      {stage1_11[229]}
   );
   gpc1_1 gpc3189 (
      {stage0_11[424]},
      {stage1_11[230]}
   );
   gpc1_1 gpc3190 (
      {stage0_11[425]},
      {stage1_11[231]}
   );
   gpc1_1 gpc3191 (
      {stage0_11[426]},
      {stage1_11[232]}
   );
   gpc1_1 gpc3192 (
      {stage0_11[427]},
      {stage1_11[233]}
   );
   gpc1_1 gpc3193 (
      {stage0_11[428]},
      {stage1_11[234]}
   );
   gpc1_1 gpc3194 (
      {stage0_11[429]},
      {stage1_11[235]}
   );
   gpc1_1 gpc3195 (
      {stage0_11[430]},
      {stage1_11[236]}
   );
   gpc1_1 gpc3196 (
      {stage0_11[431]},
      {stage1_11[237]}
   );
   gpc1_1 gpc3197 (
      {stage0_11[432]},
      {stage1_11[238]}
   );
   gpc1_1 gpc3198 (
      {stage0_11[433]},
      {stage1_11[239]}
   );
   gpc1_1 gpc3199 (
      {stage0_11[434]},
      {stage1_11[240]}
   );
   gpc1_1 gpc3200 (
      {stage0_11[435]},
      {stage1_11[241]}
   );
   gpc1_1 gpc3201 (
      {stage0_11[436]},
      {stage1_11[242]}
   );
   gpc1_1 gpc3202 (
      {stage0_11[437]},
      {stage1_11[243]}
   );
   gpc1_1 gpc3203 (
      {stage0_11[438]},
      {stage1_11[244]}
   );
   gpc1_1 gpc3204 (
      {stage0_11[439]},
      {stage1_11[245]}
   );
   gpc1_1 gpc3205 (
      {stage0_11[440]},
      {stage1_11[246]}
   );
   gpc1_1 gpc3206 (
      {stage0_11[441]},
      {stage1_11[247]}
   );
   gpc1_1 gpc3207 (
      {stage0_11[442]},
      {stage1_11[248]}
   );
   gpc1_1 gpc3208 (
      {stage0_11[443]},
      {stage1_11[249]}
   );
   gpc1_1 gpc3209 (
      {stage0_11[444]},
      {stage1_11[250]}
   );
   gpc1_1 gpc3210 (
      {stage0_11[445]},
      {stage1_11[251]}
   );
   gpc1_1 gpc3211 (
      {stage0_11[446]},
      {stage1_11[252]}
   );
   gpc1_1 gpc3212 (
      {stage0_11[447]},
      {stage1_11[253]}
   );
   gpc1_1 gpc3213 (
      {stage0_11[448]},
      {stage1_11[254]}
   );
   gpc1_1 gpc3214 (
      {stage0_11[449]},
      {stage1_11[255]}
   );
   gpc1_1 gpc3215 (
      {stage0_11[450]},
      {stage1_11[256]}
   );
   gpc1_1 gpc3216 (
      {stage0_11[451]},
      {stage1_11[257]}
   );
   gpc1_1 gpc3217 (
      {stage0_11[452]},
      {stage1_11[258]}
   );
   gpc1_1 gpc3218 (
      {stage0_11[453]},
      {stage1_11[259]}
   );
   gpc1_1 gpc3219 (
      {stage0_11[454]},
      {stage1_11[260]}
   );
   gpc1_1 gpc3220 (
      {stage0_11[455]},
      {stage1_11[261]}
   );
   gpc1_1 gpc3221 (
      {stage0_11[456]},
      {stage1_11[262]}
   );
   gpc1_1 gpc3222 (
      {stage0_11[457]},
      {stage1_11[263]}
   );
   gpc1_1 gpc3223 (
      {stage0_11[458]},
      {stage1_11[264]}
   );
   gpc1_1 gpc3224 (
      {stage0_11[459]},
      {stage1_11[265]}
   );
   gpc1_1 gpc3225 (
      {stage0_11[460]},
      {stage1_11[266]}
   );
   gpc1_1 gpc3226 (
      {stage0_11[461]},
      {stage1_11[267]}
   );
   gpc1_1 gpc3227 (
      {stage0_11[462]},
      {stage1_11[268]}
   );
   gpc1_1 gpc3228 (
      {stage0_11[463]},
      {stage1_11[269]}
   );
   gpc1_1 gpc3229 (
      {stage0_11[464]},
      {stage1_11[270]}
   );
   gpc1_1 gpc3230 (
      {stage0_11[465]},
      {stage1_11[271]}
   );
   gpc1_1 gpc3231 (
      {stage0_11[466]},
      {stage1_11[272]}
   );
   gpc1_1 gpc3232 (
      {stage0_11[467]},
      {stage1_11[273]}
   );
   gpc1_1 gpc3233 (
      {stage0_11[468]},
      {stage1_11[274]}
   );
   gpc1_1 gpc3234 (
      {stage0_11[469]},
      {stage1_11[275]}
   );
   gpc1_1 gpc3235 (
      {stage0_11[470]},
      {stage1_11[276]}
   );
   gpc1_1 gpc3236 (
      {stage0_11[471]},
      {stage1_11[277]}
   );
   gpc1_1 gpc3237 (
      {stage0_11[472]},
      {stage1_11[278]}
   );
   gpc1_1 gpc3238 (
      {stage0_11[473]},
      {stage1_11[279]}
   );
   gpc1_1 gpc3239 (
      {stage0_11[474]},
      {stage1_11[280]}
   );
   gpc1_1 gpc3240 (
      {stage0_11[475]},
      {stage1_11[281]}
   );
   gpc1_1 gpc3241 (
      {stage0_11[476]},
      {stage1_11[282]}
   );
   gpc1_1 gpc3242 (
      {stage0_11[477]},
      {stage1_11[283]}
   );
   gpc1_1 gpc3243 (
      {stage0_11[478]},
      {stage1_11[284]}
   );
   gpc1_1 gpc3244 (
      {stage0_11[479]},
      {stage1_11[285]}
   );
   gpc1_1 gpc3245 (
      {stage0_11[480]},
      {stage1_11[286]}
   );
   gpc1_1 gpc3246 (
      {stage0_11[481]},
      {stage1_11[287]}
   );
   gpc1_1 gpc3247 (
      {stage0_11[482]},
      {stage1_11[288]}
   );
   gpc1_1 gpc3248 (
      {stage0_11[483]},
      {stage1_11[289]}
   );
   gpc1_1 gpc3249 (
      {stage0_11[484]},
      {stage1_11[290]}
   );
   gpc1_1 gpc3250 (
      {stage0_11[485]},
      {stage1_11[291]}
   );
   gpc1_1 gpc3251 (
      {stage0_11[486]},
      {stage1_11[292]}
   );
   gpc1_1 gpc3252 (
      {stage0_11[487]},
      {stage1_11[293]}
   );
   gpc1_1 gpc3253 (
      {stage0_11[488]},
      {stage1_11[294]}
   );
   gpc1_1 gpc3254 (
      {stage0_11[489]},
      {stage1_11[295]}
   );
   gpc1_1 gpc3255 (
      {stage0_11[490]},
      {stage1_11[296]}
   );
   gpc1_1 gpc3256 (
      {stage0_11[491]},
      {stage1_11[297]}
   );
   gpc1_1 gpc3257 (
      {stage0_11[492]},
      {stage1_11[298]}
   );
   gpc1_1 gpc3258 (
      {stage0_11[493]},
      {stage1_11[299]}
   );
   gpc1_1 gpc3259 (
      {stage0_11[494]},
      {stage1_11[300]}
   );
   gpc1_1 gpc3260 (
      {stage0_11[495]},
      {stage1_11[301]}
   );
   gpc1_1 gpc3261 (
      {stage0_11[496]},
      {stage1_11[302]}
   );
   gpc1_1 gpc3262 (
      {stage0_11[497]},
      {stage1_11[303]}
   );
   gpc1_1 gpc3263 (
      {stage0_11[498]},
      {stage1_11[304]}
   );
   gpc1_1 gpc3264 (
      {stage0_11[499]},
      {stage1_11[305]}
   );
   gpc1_1 gpc3265 (
      {stage0_11[500]},
      {stage1_11[306]}
   );
   gpc1_1 gpc3266 (
      {stage0_11[501]},
      {stage1_11[307]}
   );
   gpc1_1 gpc3267 (
      {stage0_11[502]},
      {stage1_11[308]}
   );
   gpc1_1 gpc3268 (
      {stage0_11[503]},
      {stage1_11[309]}
   );
   gpc1_1 gpc3269 (
      {stage0_11[504]},
      {stage1_11[310]}
   );
   gpc1_1 gpc3270 (
      {stage0_11[505]},
      {stage1_11[311]}
   );
   gpc1_1 gpc3271 (
      {stage0_11[506]},
      {stage1_11[312]}
   );
   gpc1_1 gpc3272 (
      {stage0_11[507]},
      {stage1_11[313]}
   );
   gpc1_1 gpc3273 (
      {stage0_11[508]},
      {stage1_11[314]}
   );
   gpc1_1 gpc3274 (
      {stage0_11[509]},
      {stage1_11[315]}
   );
   gpc1_1 gpc3275 (
      {stage0_11[510]},
      {stage1_11[316]}
   );
   gpc1_1 gpc3276 (
      {stage0_11[511]},
      {stage1_11[317]}
   );
   gpc1_1 gpc3277 (
      {stage0_14[429]},
      {stage1_14[173]}
   );
   gpc1_1 gpc3278 (
      {stage0_14[430]},
      {stage1_14[174]}
   );
   gpc1_1 gpc3279 (
      {stage0_14[431]},
      {stage1_14[175]}
   );
   gpc1_1 gpc3280 (
      {stage0_14[432]},
      {stage1_14[176]}
   );
   gpc1_1 gpc3281 (
      {stage0_14[433]},
      {stage1_14[177]}
   );
   gpc1_1 gpc3282 (
      {stage0_14[434]},
      {stage1_14[178]}
   );
   gpc1_1 gpc3283 (
      {stage0_14[435]},
      {stage1_14[179]}
   );
   gpc1_1 gpc3284 (
      {stage0_14[436]},
      {stage1_14[180]}
   );
   gpc1_1 gpc3285 (
      {stage0_14[437]},
      {stage1_14[181]}
   );
   gpc1_1 gpc3286 (
      {stage0_14[438]},
      {stage1_14[182]}
   );
   gpc1_1 gpc3287 (
      {stage0_14[439]},
      {stage1_14[183]}
   );
   gpc1_1 gpc3288 (
      {stage0_14[440]},
      {stage1_14[184]}
   );
   gpc1_1 gpc3289 (
      {stage0_14[441]},
      {stage1_14[185]}
   );
   gpc1_1 gpc3290 (
      {stage0_14[442]},
      {stage1_14[186]}
   );
   gpc1_1 gpc3291 (
      {stage0_14[443]},
      {stage1_14[187]}
   );
   gpc1_1 gpc3292 (
      {stage0_14[444]},
      {stage1_14[188]}
   );
   gpc1_1 gpc3293 (
      {stage0_14[445]},
      {stage1_14[189]}
   );
   gpc1_1 gpc3294 (
      {stage0_14[446]},
      {stage1_14[190]}
   );
   gpc1_1 gpc3295 (
      {stage0_14[447]},
      {stage1_14[191]}
   );
   gpc1_1 gpc3296 (
      {stage0_14[448]},
      {stage1_14[192]}
   );
   gpc1_1 gpc3297 (
      {stage0_14[449]},
      {stage1_14[193]}
   );
   gpc1_1 gpc3298 (
      {stage0_14[450]},
      {stage1_14[194]}
   );
   gpc1_1 gpc3299 (
      {stage0_14[451]},
      {stage1_14[195]}
   );
   gpc1_1 gpc3300 (
      {stage0_14[452]},
      {stage1_14[196]}
   );
   gpc1_1 gpc3301 (
      {stage0_14[453]},
      {stage1_14[197]}
   );
   gpc1_1 gpc3302 (
      {stage0_14[454]},
      {stage1_14[198]}
   );
   gpc1_1 gpc3303 (
      {stage0_14[455]},
      {stage1_14[199]}
   );
   gpc1_1 gpc3304 (
      {stage0_14[456]},
      {stage1_14[200]}
   );
   gpc1_1 gpc3305 (
      {stage0_14[457]},
      {stage1_14[201]}
   );
   gpc1_1 gpc3306 (
      {stage0_14[458]},
      {stage1_14[202]}
   );
   gpc1_1 gpc3307 (
      {stage0_14[459]},
      {stage1_14[203]}
   );
   gpc1_1 gpc3308 (
      {stage0_14[460]},
      {stage1_14[204]}
   );
   gpc1_1 gpc3309 (
      {stage0_14[461]},
      {stage1_14[205]}
   );
   gpc1_1 gpc3310 (
      {stage0_14[462]},
      {stage1_14[206]}
   );
   gpc1_1 gpc3311 (
      {stage0_14[463]},
      {stage1_14[207]}
   );
   gpc1_1 gpc3312 (
      {stage0_14[464]},
      {stage1_14[208]}
   );
   gpc1_1 gpc3313 (
      {stage0_14[465]},
      {stage1_14[209]}
   );
   gpc1_1 gpc3314 (
      {stage0_14[466]},
      {stage1_14[210]}
   );
   gpc1_1 gpc3315 (
      {stage0_14[467]},
      {stage1_14[211]}
   );
   gpc1_1 gpc3316 (
      {stage0_14[468]},
      {stage1_14[212]}
   );
   gpc1_1 gpc3317 (
      {stage0_14[469]},
      {stage1_14[213]}
   );
   gpc1_1 gpc3318 (
      {stage0_14[470]},
      {stage1_14[214]}
   );
   gpc1_1 gpc3319 (
      {stage0_14[471]},
      {stage1_14[215]}
   );
   gpc1_1 gpc3320 (
      {stage0_14[472]},
      {stage1_14[216]}
   );
   gpc1_1 gpc3321 (
      {stage0_14[473]},
      {stage1_14[217]}
   );
   gpc1_1 gpc3322 (
      {stage0_14[474]},
      {stage1_14[218]}
   );
   gpc1_1 gpc3323 (
      {stage0_14[475]},
      {stage1_14[219]}
   );
   gpc1_1 gpc3324 (
      {stage0_14[476]},
      {stage1_14[220]}
   );
   gpc1_1 gpc3325 (
      {stage0_14[477]},
      {stage1_14[221]}
   );
   gpc1_1 gpc3326 (
      {stage0_14[478]},
      {stage1_14[222]}
   );
   gpc1_1 gpc3327 (
      {stage0_14[479]},
      {stage1_14[223]}
   );
   gpc1_1 gpc3328 (
      {stage0_14[480]},
      {stage1_14[224]}
   );
   gpc1_1 gpc3329 (
      {stage0_14[481]},
      {stage1_14[225]}
   );
   gpc1_1 gpc3330 (
      {stage0_14[482]},
      {stage1_14[226]}
   );
   gpc1_1 gpc3331 (
      {stage0_14[483]},
      {stage1_14[227]}
   );
   gpc1_1 gpc3332 (
      {stage0_14[484]},
      {stage1_14[228]}
   );
   gpc1_1 gpc3333 (
      {stage0_14[485]},
      {stage1_14[229]}
   );
   gpc1_1 gpc3334 (
      {stage0_14[486]},
      {stage1_14[230]}
   );
   gpc1_1 gpc3335 (
      {stage0_14[487]},
      {stage1_14[231]}
   );
   gpc1_1 gpc3336 (
      {stage0_14[488]},
      {stage1_14[232]}
   );
   gpc1_1 gpc3337 (
      {stage0_14[489]},
      {stage1_14[233]}
   );
   gpc1_1 gpc3338 (
      {stage0_14[490]},
      {stage1_14[234]}
   );
   gpc1_1 gpc3339 (
      {stage0_14[491]},
      {stage1_14[235]}
   );
   gpc1_1 gpc3340 (
      {stage0_14[492]},
      {stage1_14[236]}
   );
   gpc1_1 gpc3341 (
      {stage0_14[493]},
      {stage1_14[237]}
   );
   gpc1_1 gpc3342 (
      {stage0_14[494]},
      {stage1_14[238]}
   );
   gpc1_1 gpc3343 (
      {stage0_14[495]},
      {stage1_14[239]}
   );
   gpc1_1 gpc3344 (
      {stage0_14[496]},
      {stage1_14[240]}
   );
   gpc1_1 gpc3345 (
      {stage0_14[497]},
      {stage1_14[241]}
   );
   gpc1_1 gpc3346 (
      {stage0_14[498]},
      {stage1_14[242]}
   );
   gpc1_1 gpc3347 (
      {stage0_14[499]},
      {stage1_14[243]}
   );
   gpc1_1 gpc3348 (
      {stage0_14[500]},
      {stage1_14[244]}
   );
   gpc1_1 gpc3349 (
      {stage0_14[501]},
      {stage1_14[245]}
   );
   gpc1_1 gpc3350 (
      {stage0_14[502]},
      {stage1_14[246]}
   );
   gpc1_1 gpc3351 (
      {stage0_14[503]},
      {stage1_14[247]}
   );
   gpc1_1 gpc3352 (
      {stage0_14[504]},
      {stage1_14[248]}
   );
   gpc1_1 gpc3353 (
      {stage0_14[505]},
      {stage1_14[249]}
   );
   gpc1_1 gpc3354 (
      {stage0_14[506]},
      {stage1_14[250]}
   );
   gpc1_1 gpc3355 (
      {stage0_14[507]},
      {stage1_14[251]}
   );
   gpc1_1 gpc3356 (
      {stage0_14[508]},
      {stage1_14[252]}
   );
   gpc1_1 gpc3357 (
      {stage0_14[509]},
      {stage1_14[253]}
   );
   gpc1_1 gpc3358 (
      {stage0_14[510]},
      {stage1_14[254]}
   );
   gpc1_1 gpc3359 (
      {stage0_14[511]},
      {stage1_14[255]}
   );
   gpc1_1 gpc3360 (
      {stage0_15[457]},
      {stage1_15[203]}
   );
   gpc1_1 gpc3361 (
      {stage0_15[458]},
      {stage1_15[204]}
   );
   gpc1_1 gpc3362 (
      {stage0_15[459]},
      {stage1_15[205]}
   );
   gpc1_1 gpc3363 (
      {stage0_15[460]},
      {stage1_15[206]}
   );
   gpc1_1 gpc3364 (
      {stage0_15[461]},
      {stage1_15[207]}
   );
   gpc1_1 gpc3365 (
      {stage0_15[462]},
      {stage1_15[208]}
   );
   gpc1_1 gpc3366 (
      {stage0_15[463]},
      {stage1_15[209]}
   );
   gpc1_1 gpc3367 (
      {stage0_15[464]},
      {stage1_15[210]}
   );
   gpc1_1 gpc3368 (
      {stage0_15[465]},
      {stage1_15[211]}
   );
   gpc1_1 gpc3369 (
      {stage0_15[466]},
      {stage1_15[212]}
   );
   gpc1_1 gpc3370 (
      {stage0_15[467]},
      {stage1_15[213]}
   );
   gpc1_1 gpc3371 (
      {stage0_15[468]},
      {stage1_15[214]}
   );
   gpc1_1 gpc3372 (
      {stage0_15[469]},
      {stage1_15[215]}
   );
   gpc1_1 gpc3373 (
      {stage0_15[470]},
      {stage1_15[216]}
   );
   gpc1_1 gpc3374 (
      {stage0_15[471]},
      {stage1_15[217]}
   );
   gpc1_1 gpc3375 (
      {stage0_15[472]},
      {stage1_15[218]}
   );
   gpc1_1 gpc3376 (
      {stage0_15[473]},
      {stage1_15[219]}
   );
   gpc1_1 gpc3377 (
      {stage0_15[474]},
      {stage1_15[220]}
   );
   gpc1_1 gpc3378 (
      {stage0_15[475]},
      {stage1_15[221]}
   );
   gpc1_1 gpc3379 (
      {stage0_15[476]},
      {stage1_15[222]}
   );
   gpc1_1 gpc3380 (
      {stage0_15[477]},
      {stage1_15[223]}
   );
   gpc1_1 gpc3381 (
      {stage0_15[478]},
      {stage1_15[224]}
   );
   gpc1_1 gpc3382 (
      {stage0_15[479]},
      {stage1_15[225]}
   );
   gpc1_1 gpc3383 (
      {stage0_15[480]},
      {stage1_15[226]}
   );
   gpc1_1 gpc3384 (
      {stage0_15[481]},
      {stage1_15[227]}
   );
   gpc1_1 gpc3385 (
      {stage0_15[482]},
      {stage1_15[228]}
   );
   gpc1_1 gpc3386 (
      {stage0_15[483]},
      {stage1_15[229]}
   );
   gpc1_1 gpc3387 (
      {stage0_15[484]},
      {stage1_15[230]}
   );
   gpc1_1 gpc3388 (
      {stage0_15[485]},
      {stage1_15[231]}
   );
   gpc1_1 gpc3389 (
      {stage0_15[486]},
      {stage1_15[232]}
   );
   gpc1_1 gpc3390 (
      {stage0_15[487]},
      {stage1_15[233]}
   );
   gpc1_1 gpc3391 (
      {stage0_15[488]},
      {stage1_15[234]}
   );
   gpc1_1 gpc3392 (
      {stage0_15[489]},
      {stage1_15[235]}
   );
   gpc1_1 gpc3393 (
      {stage0_15[490]},
      {stage1_15[236]}
   );
   gpc1_1 gpc3394 (
      {stage0_15[491]},
      {stage1_15[237]}
   );
   gpc1_1 gpc3395 (
      {stage0_15[492]},
      {stage1_15[238]}
   );
   gpc1_1 gpc3396 (
      {stage0_15[493]},
      {stage1_15[239]}
   );
   gpc1_1 gpc3397 (
      {stage0_15[494]},
      {stage1_15[240]}
   );
   gpc1_1 gpc3398 (
      {stage0_15[495]},
      {stage1_15[241]}
   );
   gpc1_1 gpc3399 (
      {stage0_15[496]},
      {stage1_15[242]}
   );
   gpc1_1 gpc3400 (
      {stage0_15[497]},
      {stage1_15[243]}
   );
   gpc1_1 gpc3401 (
      {stage0_15[498]},
      {stage1_15[244]}
   );
   gpc1_1 gpc3402 (
      {stage0_15[499]},
      {stage1_15[245]}
   );
   gpc1_1 gpc3403 (
      {stage0_15[500]},
      {stage1_15[246]}
   );
   gpc1_1 gpc3404 (
      {stage0_15[501]},
      {stage1_15[247]}
   );
   gpc1_1 gpc3405 (
      {stage0_15[502]},
      {stage1_15[248]}
   );
   gpc1_1 gpc3406 (
      {stage0_15[503]},
      {stage1_15[249]}
   );
   gpc1_1 gpc3407 (
      {stage0_15[504]},
      {stage1_15[250]}
   );
   gpc1_1 gpc3408 (
      {stage0_15[505]},
      {stage1_15[251]}
   );
   gpc1_1 gpc3409 (
      {stage0_15[506]},
      {stage1_15[252]}
   );
   gpc1_1 gpc3410 (
      {stage0_15[507]},
      {stage1_15[253]}
   );
   gpc1_1 gpc3411 (
      {stage0_15[508]},
      {stage1_15[254]}
   );
   gpc1_1 gpc3412 (
      {stage0_15[509]},
      {stage1_15[255]}
   );
   gpc1_1 gpc3413 (
      {stage0_15[510]},
      {stage1_15[256]}
   );
   gpc1_1 gpc3414 (
      {stage0_15[511]},
      {stage1_15[257]}
   );
   gpc1_1 gpc3415 (
      {stage0_17[492]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3416 (
      {stage0_17[493]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3417 (
      {stage0_17[494]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3418 (
      {stage0_17[495]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3419 (
      {stage0_17[496]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3420 (
      {stage0_17[497]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3421 (
      {stage0_17[498]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3422 (
      {stage0_17[499]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3423 (
      {stage0_17[500]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3424 (
      {stage0_17[501]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3425 (
      {stage0_17[502]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3426 (
      {stage0_17[503]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3427 (
      {stage0_17[504]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3428 (
      {stage0_17[505]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3429 (
      {stage0_17[506]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3430 (
      {stage0_17[507]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3431 (
      {stage0_17[508]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3432 (
      {stage0_17[509]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3433 (
      {stage0_17[510]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3434 (
      {stage0_17[511]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3435 (
      {stage0_18[434]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3436 (
      {stage0_18[435]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3437 (
      {stage0_18[436]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3438 (
      {stage0_18[437]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3439 (
      {stage0_18[438]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3440 (
      {stage0_18[439]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3441 (
      {stage0_18[440]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3442 (
      {stage0_18[441]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3443 (
      {stage0_18[442]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3444 (
      {stage0_18[443]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3445 (
      {stage0_18[444]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3446 (
      {stage0_18[445]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3447 (
      {stage0_18[446]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3448 (
      {stage0_18[447]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3449 (
      {stage0_18[448]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3450 (
      {stage0_18[449]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3451 (
      {stage0_18[450]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3452 (
      {stage0_18[451]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3453 (
      {stage0_18[452]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3454 (
      {stage0_18[453]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3455 (
      {stage0_18[454]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3456 (
      {stage0_18[455]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3457 (
      {stage0_18[456]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3458 (
      {stage0_18[457]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3459 (
      {stage0_18[458]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3460 (
      {stage0_18[459]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3461 (
      {stage0_18[460]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3462 (
      {stage0_18[461]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3463 (
      {stage0_18[462]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3464 (
      {stage0_18[463]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3465 (
      {stage0_18[464]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3466 (
      {stage0_18[465]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3467 (
      {stage0_18[466]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3468 (
      {stage0_18[467]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3469 (
      {stage0_18[468]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3470 (
      {stage0_18[469]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3471 (
      {stage0_18[470]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3472 (
      {stage0_18[471]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3473 (
      {stage0_18[472]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3474 (
      {stage0_18[473]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3475 (
      {stage0_18[474]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3476 (
      {stage0_18[475]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3477 (
      {stage0_18[476]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3478 (
      {stage0_18[477]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3479 (
      {stage0_18[478]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3480 (
      {stage0_18[479]},
      {stage1_18[209]}
   );
   gpc1_1 gpc3481 (
      {stage0_18[480]},
      {stage1_18[210]}
   );
   gpc1_1 gpc3482 (
      {stage0_18[481]},
      {stage1_18[211]}
   );
   gpc1_1 gpc3483 (
      {stage0_18[482]},
      {stage1_18[212]}
   );
   gpc1_1 gpc3484 (
      {stage0_18[483]},
      {stage1_18[213]}
   );
   gpc1_1 gpc3485 (
      {stage0_18[484]},
      {stage1_18[214]}
   );
   gpc1_1 gpc3486 (
      {stage0_18[485]},
      {stage1_18[215]}
   );
   gpc1_1 gpc3487 (
      {stage0_18[486]},
      {stage1_18[216]}
   );
   gpc1_1 gpc3488 (
      {stage0_18[487]},
      {stage1_18[217]}
   );
   gpc1_1 gpc3489 (
      {stage0_18[488]},
      {stage1_18[218]}
   );
   gpc1_1 gpc3490 (
      {stage0_18[489]},
      {stage1_18[219]}
   );
   gpc1_1 gpc3491 (
      {stage0_18[490]},
      {stage1_18[220]}
   );
   gpc1_1 gpc3492 (
      {stage0_18[491]},
      {stage1_18[221]}
   );
   gpc1_1 gpc3493 (
      {stage0_18[492]},
      {stage1_18[222]}
   );
   gpc1_1 gpc3494 (
      {stage0_18[493]},
      {stage1_18[223]}
   );
   gpc1_1 gpc3495 (
      {stage0_18[494]},
      {stage1_18[224]}
   );
   gpc1_1 gpc3496 (
      {stage0_18[495]},
      {stage1_18[225]}
   );
   gpc1_1 gpc3497 (
      {stage0_18[496]},
      {stage1_18[226]}
   );
   gpc1_1 gpc3498 (
      {stage0_18[497]},
      {stage1_18[227]}
   );
   gpc1_1 gpc3499 (
      {stage0_18[498]},
      {stage1_18[228]}
   );
   gpc1_1 gpc3500 (
      {stage0_18[499]},
      {stage1_18[229]}
   );
   gpc1_1 gpc3501 (
      {stage0_18[500]},
      {stage1_18[230]}
   );
   gpc1_1 gpc3502 (
      {stage0_18[501]},
      {stage1_18[231]}
   );
   gpc1_1 gpc3503 (
      {stage0_18[502]},
      {stage1_18[232]}
   );
   gpc1_1 gpc3504 (
      {stage0_18[503]},
      {stage1_18[233]}
   );
   gpc1_1 gpc3505 (
      {stage0_18[504]},
      {stage1_18[234]}
   );
   gpc1_1 gpc3506 (
      {stage0_18[505]},
      {stage1_18[235]}
   );
   gpc1_1 gpc3507 (
      {stage0_18[506]},
      {stage1_18[236]}
   );
   gpc1_1 gpc3508 (
      {stage0_18[507]},
      {stage1_18[237]}
   );
   gpc1_1 gpc3509 (
      {stage0_18[508]},
      {stage1_18[238]}
   );
   gpc1_1 gpc3510 (
      {stage0_18[509]},
      {stage1_18[239]}
   );
   gpc1_1 gpc3511 (
      {stage0_18[510]},
      {stage1_18[240]}
   );
   gpc1_1 gpc3512 (
      {stage0_18[511]},
      {stage1_18[241]}
   );
   gpc1_1 gpc3513 (
      {stage0_19[502]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3514 (
      {stage0_19[503]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3515 (
      {stage0_19[504]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3516 (
      {stage0_19[505]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3517 (
      {stage0_19[506]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3518 (
      {stage0_19[507]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3519 (
      {stage0_19[508]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3520 (
      {stage0_19[509]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3521 (
      {stage0_19[510]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3522 (
      {stage0_19[511]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3523 (
      {stage0_20[504]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3524 (
      {stage0_20[505]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3525 (
      {stage0_20[506]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3526 (
      {stage0_20[507]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3527 (
      {stage0_20[508]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3528 (
      {stage0_20[509]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3529 (
      {stage0_20[510]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3530 (
      {stage0_20[511]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3531 (
      {stage0_21[504]},
      {stage1_21[197]}
   );
   gpc1_1 gpc3532 (
      {stage0_21[505]},
      {stage1_21[198]}
   );
   gpc1_1 gpc3533 (
      {stage0_21[506]},
      {stage1_21[199]}
   );
   gpc1_1 gpc3534 (
      {stage0_21[507]},
      {stage1_21[200]}
   );
   gpc1_1 gpc3535 (
      {stage0_21[508]},
      {stage1_21[201]}
   );
   gpc1_1 gpc3536 (
      {stage0_21[509]},
      {stage1_21[202]}
   );
   gpc1_1 gpc3537 (
      {stage0_21[510]},
      {stage1_21[203]}
   );
   gpc1_1 gpc3538 (
      {stage0_21[511]},
      {stage1_21[204]}
   );
   gpc1_1 gpc3539 (
      {stage0_22[481]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3540 (
      {stage0_22[482]},
      {stage1_22[171]}
   );
   gpc1_1 gpc3541 (
      {stage0_22[483]},
      {stage1_22[172]}
   );
   gpc1_1 gpc3542 (
      {stage0_22[484]},
      {stage1_22[173]}
   );
   gpc1_1 gpc3543 (
      {stage0_22[485]},
      {stage1_22[174]}
   );
   gpc1_1 gpc3544 (
      {stage0_22[486]},
      {stage1_22[175]}
   );
   gpc1_1 gpc3545 (
      {stage0_22[487]},
      {stage1_22[176]}
   );
   gpc1_1 gpc3546 (
      {stage0_22[488]},
      {stage1_22[177]}
   );
   gpc1_1 gpc3547 (
      {stage0_22[489]},
      {stage1_22[178]}
   );
   gpc1_1 gpc3548 (
      {stage0_22[490]},
      {stage1_22[179]}
   );
   gpc1_1 gpc3549 (
      {stage0_22[491]},
      {stage1_22[180]}
   );
   gpc1_1 gpc3550 (
      {stage0_22[492]},
      {stage1_22[181]}
   );
   gpc1_1 gpc3551 (
      {stage0_22[493]},
      {stage1_22[182]}
   );
   gpc1_1 gpc3552 (
      {stage0_22[494]},
      {stage1_22[183]}
   );
   gpc1_1 gpc3553 (
      {stage0_22[495]},
      {stage1_22[184]}
   );
   gpc1_1 gpc3554 (
      {stage0_22[496]},
      {stage1_22[185]}
   );
   gpc1_1 gpc3555 (
      {stage0_22[497]},
      {stage1_22[186]}
   );
   gpc1_1 gpc3556 (
      {stage0_22[498]},
      {stage1_22[187]}
   );
   gpc1_1 gpc3557 (
      {stage0_22[499]},
      {stage1_22[188]}
   );
   gpc1_1 gpc3558 (
      {stage0_22[500]},
      {stage1_22[189]}
   );
   gpc1_1 gpc3559 (
      {stage0_22[501]},
      {stage1_22[190]}
   );
   gpc1_1 gpc3560 (
      {stage0_22[502]},
      {stage1_22[191]}
   );
   gpc1_1 gpc3561 (
      {stage0_22[503]},
      {stage1_22[192]}
   );
   gpc1_1 gpc3562 (
      {stage0_22[504]},
      {stage1_22[193]}
   );
   gpc1_1 gpc3563 (
      {stage0_22[505]},
      {stage1_22[194]}
   );
   gpc1_1 gpc3564 (
      {stage0_22[506]},
      {stage1_22[195]}
   );
   gpc1_1 gpc3565 (
      {stage0_22[507]},
      {stage1_22[196]}
   );
   gpc1_1 gpc3566 (
      {stage0_22[508]},
      {stage1_22[197]}
   );
   gpc1_1 gpc3567 (
      {stage0_22[509]},
      {stage1_22[198]}
   );
   gpc1_1 gpc3568 (
      {stage0_22[510]},
      {stage1_22[199]}
   );
   gpc1_1 gpc3569 (
      {stage0_22[511]},
      {stage1_22[200]}
   );
   gpc1_1 gpc3570 (
      {stage0_23[418]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3571 (
      {stage0_23[419]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3572 (
      {stage0_23[420]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3573 (
      {stage0_23[421]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3574 (
      {stage0_23[422]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3575 (
      {stage0_23[423]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3576 (
      {stage0_23[424]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3577 (
      {stage0_23[425]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3578 (
      {stage0_23[426]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3579 (
      {stage0_23[427]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3580 (
      {stage0_23[428]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3581 (
      {stage0_23[429]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3582 (
      {stage0_23[430]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3583 (
      {stage0_23[431]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3584 (
      {stage0_23[432]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3585 (
      {stage0_23[433]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3586 (
      {stage0_23[434]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3587 (
      {stage0_23[435]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3588 (
      {stage0_23[436]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3589 (
      {stage0_23[437]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3590 (
      {stage0_23[438]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3591 (
      {stage0_23[439]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3592 (
      {stage0_23[440]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3593 (
      {stage0_23[441]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3594 (
      {stage0_23[442]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3595 (
      {stage0_23[443]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3596 (
      {stage0_23[444]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3597 (
      {stage0_23[445]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3598 (
      {stage0_23[446]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3599 (
      {stage0_23[447]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3600 (
      {stage0_23[448]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3601 (
      {stage0_23[449]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3602 (
      {stage0_23[450]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3603 (
      {stage0_23[451]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3604 (
      {stage0_23[452]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3605 (
      {stage0_23[453]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3606 (
      {stage0_23[454]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3607 (
      {stage0_23[455]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3608 (
      {stage0_23[456]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3609 (
      {stage0_23[457]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3610 (
      {stage0_23[458]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3611 (
      {stage0_23[459]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3612 (
      {stage0_23[460]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3613 (
      {stage0_23[461]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3614 (
      {stage0_23[462]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3615 (
      {stage0_23[463]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3616 (
      {stage0_23[464]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3617 (
      {stage0_23[465]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3618 (
      {stage0_23[466]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3619 (
      {stage0_23[467]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3620 (
      {stage0_23[468]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3621 (
      {stage0_23[469]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3622 (
      {stage0_23[470]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3623 (
      {stage0_23[471]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3624 (
      {stage0_23[472]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3625 (
      {stage0_23[473]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3626 (
      {stage0_23[474]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3627 (
      {stage0_23[475]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3628 (
      {stage0_23[476]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3629 (
      {stage0_23[477]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3630 (
      {stage0_23[478]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3631 (
      {stage0_23[479]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3632 (
      {stage0_23[480]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3633 (
      {stage0_23[481]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3634 (
      {stage0_23[482]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3635 (
      {stage0_23[483]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3636 (
      {stage0_23[484]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3637 (
      {stage0_23[485]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3638 (
      {stage0_23[486]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3639 (
      {stage0_23[487]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3640 (
      {stage0_23[488]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3641 (
      {stage0_23[489]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3642 (
      {stage0_23[490]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3643 (
      {stage0_23[491]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3644 (
      {stage0_23[492]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3645 (
      {stage0_23[493]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3646 (
      {stage0_23[494]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3647 (
      {stage0_23[495]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3648 (
      {stage0_23[496]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3649 (
      {stage0_23[497]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3650 (
      {stage0_23[498]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3651 (
      {stage0_23[499]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3652 (
      {stage0_23[500]},
      {stage1_23[287]}
   );
   gpc1_1 gpc3653 (
      {stage0_23[501]},
      {stage1_23[288]}
   );
   gpc1_1 gpc3654 (
      {stage0_23[502]},
      {stage1_23[289]}
   );
   gpc1_1 gpc3655 (
      {stage0_23[503]},
      {stage1_23[290]}
   );
   gpc1_1 gpc3656 (
      {stage0_23[504]},
      {stage1_23[291]}
   );
   gpc1_1 gpc3657 (
      {stage0_23[505]},
      {stage1_23[292]}
   );
   gpc1_1 gpc3658 (
      {stage0_23[506]},
      {stage1_23[293]}
   );
   gpc1_1 gpc3659 (
      {stage0_23[507]},
      {stage1_23[294]}
   );
   gpc1_1 gpc3660 (
      {stage0_23[508]},
      {stage1_23[295]}
   );
   gpc1_1 gpc3661 (
      {stage0_23[509]},
      {stage1_23[296]}
   );
   gpc1_1 gpc3662 (
      {stage0_23[510]},
      {stage1_23[297]}
   );
   gpc1_1 gpc3663 (
      {stage0_23[511]},
      {stage1_23[298]}
   );
   gpc1_1 gpc3664 (
      {stage0_24[499]},
      {stage1_24[222]}
   );
   gpc1_1 gpc3665 (
      {stage0_24[500]},
      {stage1_24[223]}
   );
   gpc1_1 gpc3666 (
      {stage0_24[501]},
      {stage1_24[224]}
   );
   gpc1_1 gpc3667 (
      {stage0_24[502]},
      {stage1_24[225]}
   );
   gpc1_1 gpc3668 (
      {stage0_24[503]},
      {stage1_24[226]}
   );
   gpc1_1 gpc3669 (
      {stage0_24[504]},
      {stage1_24[227]}
   );
   gpc1_1 gpc3670 (
      {stage0_24[505]},
      {stage1_24[228]}
   );
   gpc1_1 gpc3671 (
      {stage0_24[506]},
      {stage1_24[229]}
   );
   gpc1_1 gpc3672 (
      {stage0_24[507]},
      {stage1_24[230]}
   );
   gpc1_1 gpc3673 (
      {stage0_24[508]},
      {stage1_24[231]}
   );
   gpc1_1 gpc3674 (
      {stage0_24[509]},
      {stage1_24[232]}
   );
   gpc1_1 gpc3675 (
      {stage0_24[510]},
      {stage1_24[233]}
   );
   gpc1_1 gpc3676 (
      {stage0_24[511]},
      {stage1_24[234]}
   );
   gpc1_1 gpc3677 (
      {stage0_25[506]},
      {stage1_25[205]}
   );
   gpc1_1 gpc3678 (
      {stage0_25[507]},
      {stage1_25[206]}
   );
   gpc1_1 gpc3679 (
      {stage0_25[508]},
      {stage1_25[207]}
   );
   gpc1_1 gpc3680 (
      {stage0_25[509]},
      {stage1_25[208]}
   );
   gpc1_1 gpc3681 (
      {stage0_25[510]},
      {stage1_25[209]}
   );
   gpc1_1 gpc3682 (
      {stage0_25[511]},
      {stage1_25[210]}
   );
   gpc1_1 gpc3683 (
      {stage0_26[503]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3684 (
      {stage0_26[504]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3685 (
      {stage0_26[505]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3686 (
      {stage0_26[506]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3687 (
      {stage0_26[507]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3688 (
      {stage0_26[508]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3689 (
      {stage0_26[509]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3690 (
      {stage0_26[510]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3691 (
      {stage0_26[511]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3692 (
      {stage0_27[503]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3693 (
      {stage0_27[504]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3694 (
      {stage0_27[505]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3695 (
      {stage0_27[506]},
      {stage1_27[206]}
   );
   gpc1_1 gpc3696 (
      {stage0_27[507]},
      {stage1_27[207]}
   );
   gpc1_1 gpc3697 (
      {stage0_27[508]},
      {stage1_27[208]}
   );
   gpc1_1 gpc3698 (
      {stage0_27[509]},
      {stage1_27[209]}
   );
   gpc1_1 gpc3699 (
      {stage0_27[510]},
      {stage1_27[210]}
   );
   gpc1_1 gpc3700 (
      {stage0_27[511]},
      {stage1_27[211]}
   );
   gpc1_1 gpc3701 (
      {stage0_28[500]},
      {stage1_28[237]}
   );
   gpc1_1 gpc3702 (
      {stage0_28[501]},
      {stage1_28[238]}
   );
   gpc1_1 gpc3703 (
      {stage0_28[502]},
      {stage1_28[239]}
   );
   gpc1_1 gpc3704 (
      {stage0_28[503]},
      {stage1_28[240]}
   );
   gpc1_1 gpc3705 (
      {stage0_28[504]},
      {stage1_28[241]}
   );
   gpc1_1 gpc3706 (
      {stage0_28[505]},
      {stage1_28[242]}
   );
   gpc1_1 gpc3707 (
      {stage0_28[506]},
      {stage1_28[243]}
   );
   gpc1_1 gpc3708 (
      {stage0_28[507]},
      {stage1_28[244]}
   );
   gpc1_1 gpc3709 (
      {stage0_28[508]},
      {stage1_28[245]}
   );
   gpc1_1 gpc3710 (
      {stage0_28[509]},
      {stage1_28[246]}
   );
   gpc1_1 gpc3711 (
      {stage0_28[510]},
      {stage1_28[247]}
   );
   gpc1_1 gpc3712 (
      {stage0_28[511]},
      {stage1_28[248]}
   );
   gpc1_1 gpc3713 (
      {stage0_29[510]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3714 (
      {stage0_29[511]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3715 (
      {stage0_30[443]},
      {stage1_30[164]}
   );
   gpc1_1 gpc3716 (
      {stage0_30[444]},
      {stage1_30[165]}
   );
   gpc1_1 gpc3717 (
      {stage0_30[445]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3718 (
      {stage0_30[446]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3719 (
      {stage0_30[447]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3720 (
      {stage0_30[448]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3721 (
      {stage0_30[449]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3722 (
      {stage0_30[450]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3723 (
      {stage0_30[451]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3724 (
      {stage0_30[452]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3725 (
      {stage0_30[453]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3726 (
      {stage0_30[454]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3727 (
      {stage0_30[455]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3728 (
      {stage0_30[456]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3729 (
      {stage0_30[457]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3730 (
      {stage0_30[458]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3731 (
      {stage0_30[459]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3732 (
      {stage0_30[460]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3733 (
      {stage0_30[461]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3734 (
      {stage0_30[462]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3735 (
      {stage0_30[463]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3736 (
      {stage0_30[464]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3737 (
      {stage0_30[465]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3738 (
      {stage0_30[466]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3739 (
      {stage0_30[467]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3740 (
      {stage0_30[468]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3741 (
      {stage0_30[469]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3742 (
      {stage0_30[470]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3743 (
      {stage0_30[471]},
      {stage1_30[192]}
   );
   gpc1_1 gpc3744 (
      {stage0_30[472]},
      {stage1_30[193]}
   );
   gpc1_1 gpc3745 (
      {stage0_30[473]},
      {stage1_30[194]}
   );
   gpc1_1 gpc3746 (
      {stage0_30[474]},
      {stage1_30[195]}
   );
   gpc1_1 gpc3747 (
      {stage0_30[475]},
      {stage1_30[196]}
   );
   gpc1_1 gpc3748 (
      {stage0_30[476]},
      {stage1_30[197]}
   );
   gpc1_1 gpc3749 (
      {stage0_30[477]},
      {stage1_30[198]}
   );
   gpc1_1 gpc3750 (
      {stage0_30[478]},
      {stage1_30[199]}
   );
   gpc1_1 gpc3751 (
      {stage0_30[479]},
      {stage1_30[200]}
   );
   gpc1_1 gpc3752 (
      {stage0_30[480]},
      {stage1_30[201]}
   );
   gpc1_1 gpc3753 (
      {stage0_30[481]},
      {stage1_30[202]}
   );
   gpc1_1 gpc3754 (
      {stage0_30[482]},
      {stage1_30[203]}
   );
   gpc1_1 gpc3755 (
      {stage0_30[483]},
      {stage1_30[204]}
   );
   gpc1_1 gpc3756 (
      {stage0_30[484]},
      {stage1_30[205]}
   );
   gpc1_1 gpc3757 (
      {stage0_30[485]},
      {stage1_30[206]}
   );
   gpc1_1 gpc3758 (
      {stage0_30[486]},
      {stage1_30[207]}
   );
   gpc1_1 gpc3759 (
      {stage0_30[487]},
      {stage1_30[208]}
   );
   gpc1_1 gpc3760 (
      {stage0_30[488]},
      {stage1_30[209]}
   );
   gpc1_1 gpc3761 (
      {stage0_30[489]},
      {stage1_30[210]}
   );
   gpc1_1 gpc3762 (
      {stage0_30[490]},
      {stage1_30[211]}
   );
   gpc1_1 gpc3763 (
      {stage0_30[491]},
      {stage1_30[212]}
   );
   gpc1_1 gpc3764 (
      {stage0_30[492]},
      {stage1_30[213]}
   );
   gpc1_1 gpc3765 (
      {stage0_30[493]},
      {stage1_30[214]}
   );
   gpc1_1 gpc3766 (
      {stage0_30[494]},
      {stage1_30[215]}
   );
   gpc1_1 gpc3767 (
      {stage0_30[495]},
      {stage1_30[216]}
   );
   gpc1_1 gpc3768 (
      {stage0_30[496]},
      {stage1_30[217]}
   );
   gpc1_1 gpc3769 (
      {stage0_30[497]},
      {stage1_30[218]}
   );
   gpc1_1 gpc3770 (
      {stage0_30[498]},
      {stage1_30[219]}
   );
   gpc1_1 gpc3771 (
      {stage0_30[499]},
      {stage1_30[220]}
   );
   gpc1_1 gpc3772 (
      {stage0_30[500]},
      {stage1_30[221]}
   );
   gpc1_1 gpc3773 (
      {stage0_30[501]},
      {stage1_30[222]}
   );
   gpc1_1 gpc3774 (
      {stage0_30[502]},
      {stage1_30[223]}
   );
   gpc1_1 gpc3775 (
      {stage0_30[503]},
      {stage1_30[224]}
   );
   gpc1_1 gpc3776 (
      {stage0_30[504]},
      {stage1_30[225]}
   );
   gpc1_1 gpc3777 (
      {stage0_30[505]},
      {stage1_30[226]}
   );
   gpc1_1 gpc3778 (
      {stage0_30[506]},
      {stage1_30[227]}
   );
   gpc1_1 gpc3779 (
      {stage0_30[507]},
      {stage1_30[228]}
   );
   gpc1_1 gpc3780 (
      {stage0_30[508]},
      {stage1_30[229]}
   );
   gpc1_1 gpc3781 (
      {stage0_30[509]},
      {stage1_30[230]}
   );
   gpc1_1 gpc3782 (
      {stage0_30[510]},
      {stage1_30[231]}
   );
   gpc1_1 gpc3783 (
      {stage0_30[511]},
      {stage1_30[232]}
   );
   gpc1_1 gpc3784 (
      {stage0_31[494]},
      {stage1_31[194]}
   );
   gpc1_1 gpc3785 (
      {stage0_31[495]},
      {stage1_31[195]}
   );
   gpc1_1 gpc3786 (
      {stage0_31[496]},
      {stage1_31[196]}
   );
   gpc1_1 gpc3787 (
      {stage0_31[497]},
      {stage1_31[197]}
   );
   gpc1_1 gpc3788 (
      {stage0_31[498]},
      {stage1_31[198]}
   );
   gpc1_1 gpc3789 (
      {stage0_31[499]},
      {stage1_31[199]}
   );
   gpc1_1 gpc3790 (
      {stage0_31[500]},
      {stage1_31[200]}
   );
   gpc1_1 gpc3791 (
      {stage0_31[501]},
      {stage1_31[201]}
   );
   gpc1_1 gpc3792 (
      {stage0_31[502]},
      {stage1_31[202]}
   );
   gpc1_1 gpc3793 (
      {stage0_31[503]},
      {stage1_31[203]}
   );
   gpc1_1 gpc3794 (
      {stage0_31[504]},
      {stage1_31[204]}
   );
   gpc1_1 gpc3795 (
      {stage0_31[505]},
      {stage1_31[205]}
   );
   gpc1_1 gpc3796 (
      {stage0_31[506]},
      {stage1_31[206]}
   );
   gpc1_1 gpc3797 (
      {stage0_31[507]},
      {stage1_31[207]}
   );
   gpc1_1 gpc3798 (
      {stage0_31[508]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3799 (
      {stage0_31[509]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3800 (
      {stage0_31[510]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3801 (
      {stage0_31[511]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3802 (
      {stage0_32[303]},
      {stage1_32[206]}
   );
   gpc1_1 gpc3803 (
      {stage0_32[304]},
      {stage1_32[207]}
   );
   gpc1_1 gpc3804 (
      {stage0_32[305]},
      {stage1_32[208]}
   );
   gpc1_1 gpc3805 (
      {stage0_32[306]},
      {stage1_32[209]}
   );
   gpc1_1 gpc3806 (
      {stage0_32[307]},
      {stage1_32[210]}
   );
   gpc1_1 gpc3807 (
      {stage0_32[308]},
      {stage1_32[211]}
   );
   gpc1_1 gpc3808 (
      {stage0_32[309]},
      {stage1_32[212]}
   );
   gpc1_1 gpc3809 (
      {stage0_32[310]},
      {stage1_32[213]}
   );
   gpc1_1 gpc3810 (
      {stage0_32[311]},
      {stage1_32[214]}
   );
   gpc1_1 gpc3811 (
      {stage0_32[312]},
      {stage1_32[215]}
   );
   gpc1_1 gpc3812 (
      {stage0_32[313]},
      {stage1_32[216]}
   );
   gpc1_1 gpc3813 (
      {stage0_32[314]},
      {stage1_32[217]}
   );
   gpc1_1 gpc3814 (
      {stage0_32[315]},
      {stage1_32[218]}
   );
   gpc1_1 gpc3815 (
      {stage0_32[316]},
      {stage1_32[219]}
   );
   gpc1_1 gpc3816 (
      {stage0_32[317]},
      {stage1_32[220]}
   );
   gpc1_1 gpc3817 (
      {stage0_32[318]},
      {stage1_32[221]}
   );
   gpc1_1 gpc3818 (
      {stage0_32[319]},
      {stage1_32[222]}
   );
   gpc1_1 gpc3819 (
      {stage0_32[320]},
      {stage1_32[223]}
   );
   gpc1_1 gpc3820 (
      {stage0_32[321]},
      {stage1_32[224]}
   );
   gpc1_1 gpc3821 (
      {stage0_32[322]},
      {stage1_32[225]}
   );
   gpc1_1 gpc3822 (
      {stage0_32[323]},
      {stage1_32[226]}
   );
   gpc1_1 gpc3823 (
      {stage0_32[324]},
      {stage1_32[227]}
   );
   gpc1_1 gpc3824 (
      {stage0_32[325]},
      {stage1_32[228]}
   );
   gpc1_1 gpc3825 (
      {stage0_32[326]},
      {stage1_32[229]}
   );
   gpc1_1 gpc3826 (
      {stage0_32[327]},
      {stage1_32[230]}
   );
   gpc1_1 gpc3827 (
      {stage0_32[328]},
      {stage1_32[231]}
   );
   gpc1_1 gpc3828 (
      {stage0_32[329]},
      {stage1_32[232]}
   );
   gpc1_1 gpc3829 (
      {stage0_32[330]},
      {stage1_32[233]}
   );
   gpc1_1 gpc3830 (
      {stage0_32[331]},
      {stage1_32[234]}
   );
   gpc1_1 gpc3831 (
      {stage0_32[332]},
      {stage1_32[235]}
   );
   gpc1_1 gpc3832 (
      {stage0_32[333]},
      {stage1_32[236]}
   );
   gpc1_1 gpc3833 (
      {stage0_32[334]},
      {stage1_32[237]}
   );
   gpc1_1 gpc3834 (
      {stage0_32[335]},
      {stage1_32[238]}
   );
   gpc1_1 gpc3835 (
      {stage0_32[336]},
      {stage1_32[239]}
   );
   gpc1_1 gpc3836 (
      {stage0_32[337]},
      {stage1_32[240]}
   );
   gpc1_1 gpc3837 (
      {stage0_32[338]},
      {stage1_32[241]}
   );
   gpc1_1 gpc3838 (
      {stage0_32[339]},
      {stage1_32[242]}
   );
   gpc1_1 gpc3839 (
      {stage0_32[340]},
      {stage1_32[243]}
   );
   gpc1_1 gpc3840 (
      {stage0_32[341]},
      {stage1_32[244]}
   );
   gpc1_1 gpc3841 (
      {stage0_32[342]},
      {stage1_32[245]}
   );
   gpc1_1 gpc3842 (
      {stage0_32[343]},
      {stage1_32[246]}
   );
   gpc1_1 gpc3843 (
      {stage0_32[344]},
      {stage1_32[247]}
   );
   gpc1_1 gpc3844 (
      {stage0_32[345]},
      {stage1_32[248]}
   );
   gpc1_1 gpc3845 (
      {stage0_32[346]},
      {stage1_32[249]}
   );
   gpc1_1 gpc3846 (
      {stage0_32[347]},
      {stage1_32[250]}
   );
   gpc1_1 gpc3847 (
      {stage0_32[348]},
      {stage1_32[251]}
   );
   gpc1_1 gpc3848 (
      {stage0_32[349]},
      {stage1_32[252]}
   );
   gpc1_1 gpc3849 (
      {stage0_32[350]},
      {stage1_32[253]}
   );
   gpc1_1 gpc3850 (
      {stage0_32[351]},
      {stage1_32[254]}
   );
   gpc1_1 gpc3851 (
      {stage0_32[352]},
      {stage1_32[255]}
   );
   gpc1_1 gpc3852 (
      {stage0_32[353]},
      {stage1_32[256]}
   );
   gpc1_1 gpc3853 (
      {stage0_32[354]},
      {stage1_32[257]}
   );
   gpc1_1 gpc3854 (
      {stage0_32[355]},
      {stage1_32[258]}
   );
   gpc1_1 gpc3855 (
      {stage0_32[356]},
      {stage1_32[259]}
   );
   gpc1_1 gpc3856 (
      {stage0_32[357]},
      {stage1_32[260]}
   );
   gpc1_1 gpc3857 (
      {stage0_32[358]},
      {stage1_32[261]}
   );
   gpc1_1 gpc3858 (
      {stage0_32[359]},
      {stage1_32[262]}
   );
   gpc1_1 gpc3859 (
      {stage0_32[360]},
      {stage1_32[263]}
   );
   gpc1_1 gpc3860 (
      {stage0_32[361]},
      {stage1_32[264]}
   );
   gpc1_1 gpc3861 (
      {stage0_32[362]},
      {stage1_32[265]}
   );
   gpc1_1 gpc3862 (
      {stage0_32[363]},
      {stage1_32[266]}
   );
   gpc1_1 gpc3863 (
      {stage0_32[364]},
      {stage1_32[267]}
   );
   gpc1_1 gpc3864 (
      {stage0_32[365]},
      {stage1_32[268]}
   );
   gpc1_1 gpc3865 (
      {stage0_32[366]},
      {stage1_32[269]}
   );
   gpc1_1 gpc3866 (
      {stage0_32[367]},
      {stage1_32[270]}
   );
   gpc1_1 gpc3867 (
      {stage0_32[368]},
      {stage1_32[271]}
   );
   gpc1_1 gpc3868 (
      {stage0_32[369]},
      {stage1_32[272]}
   );
   gpc1_1 gpc3869 (
      {stage0_32[370]},
      {stage1_32[273]}
   );
   gpc1_1 gpc3870 (
      {stage0_32[371]},
      {stage1_32[274]}
   );
   gpc1_1 gpc3871 (
      {stage0_32[372]},
      {stage1_32[275]}
   );
   gpc1_1 gpc3872 (
      {stage0_32[373]},
      {stage1_32[276]}
   );
   gpc1_1 gpc3873 (
      {stage0_32[374]},
      {stage1_32[277]}
   );
   gpc1_1 gpc3874 (
      {stage0_32[375]},
      {stage1_32[278]}
   );
   gpc1_1 gpc3875 (
      {stage0_32[376]},
      {stage1_32[279]}
   );
   gpc1_1 gpc3876 (
      {stage0_32[377]},
      {stage1_32[280]}
   );
   gpc1_1 gpc3877 (
      {stage0_32[378]},
      {stage1_32[281]}
   );
   gpc1_1 gpc3878 (
      {stage0_32[379]},
      {stage1_32[282]}
   );
   gpc1_1 gpc3879 (
      {stage0_32[380]},
      {stage1_32[283]}
   );
   gpc1_1 gpc3880 (
      {stage0_32[381]},
      {stage1_32[284]}
   );
   gpc1_1 gpc3881 (
      {stage0_32[382]},
      {stage1_32[285]}
   );
   gpc1_1 gpc3882 (
      {stage0_32[383]},
      {stage1_32[286]}
   );
   gpc1_1 gpc3883 (
      {stage0_32[384]},
      {stage1_32[287]}
   );
   gpc1_1 gpc3884 (
      {stage0_32[385]},
      {stage1_32[288]}
   );
   gpc1_1 gpc3885 (
      {stage0_32[386]},
      {stage1_32[289]}
   );
   gpc1_1 gpc3886 (
      {stage0_32[387]},
      {stage1_32[290]}
   );
   gpc1_1 gpc3887 (
      {stage0_32[388]},
      {stage1_32[291]}
   );
   gpc1_1 gpc3888 (
      {stage0_32[389]},
      {stage1_32[292]}
   );
   gpc1_1 gpc3889 (
      {stage0_32[390]},
      {stage1_32[293]}
   );
   gpc1_1 gpc3890 (
      {stage0_32[391]},
      {stage1_32[294]}
   );
   gpc1_1 gpc3891 (
      {stage0_32[392]},
      {stage1_32[295]}
   );
   gpc1_1 gpc3892 (
      {stage0_32[393]},
      {stage1_32[296]}
   );
   gpc1_1 gpc3893 (
      {stage0_32[394]},
      {stage1_32[297]}
   );
   gpc1_1 gpc3894 (
      {stage0_32[395]},
      {stage1_32[298]}
   );
   gpc1_1 gpc3895 (
      {stage0_32[396]},
      {stage1_32[299]}
   );
   gpc1_1 gpc3896 (
      {stage0_32[397]},
      {stage1_32[300]}
   );
   gpc1_1 gpc3897 (
      {stage0_32[398]},
      {stage1_32[301]}
   );
   gpc1_1 gpc3898 (
      {stage0_32[399]},
      {stage1_32[302]}
   );
   gpc1_1 gpc3899 (
      {stage0_32[400]},
      {stage1_32[303]}
   );
   gpc1_1 gpc3900 (
      {stage0_32[401]},
      {stage1_32[304]}
   );
   gpc1_1 gpc3901 (
      {stage0_32[402]},
      {stage1_32[305]}
   );
   gpc1_1 gpc3902 (
      {stage0_32[403]},
      {stage1_32[306]}
   );
   gpc1_1 gpc3903 (
      {stage0_32[404]},
      {stage1_32[307]}
   );
   gpc1_1 gpc3904 (
      {stage0_32[405]},
      {stage1_32[308]}
   );
   gpc1_1 gpc3905 (
      {stage0_32[406]},
      {stage1_32[309]}
   );
   gpc1_1 gpc3906 (
      {stage0_32[407]},
      {stage1_32[310]}
   );
   gpc1_1 gpc3907 (
      {stage0_32[408]},
      {stage1_32[311]}
   );
   gpc1_1 gpc3908 (
      {stage0_32[409]},
      {stage1_32[312]}
   );
   gpc1_1 gpc3909 (
      {stage0_32[410]},
      {stage1_32[313]}
   );
   gpc1_1 gpc3910 (
      {stage0_32[411]},
      {stage1_32[314]}
   );
   gpc1_1 gpc3911 (
      {stage0_32[412]},
      {stage1_32[315]}
   );
   gpc1_1 gpc3912 (
      {stage0_32[413]},
      {stage1_32[316]}
   );
   gpc1_1 gpc3913 (
      {stage0_32[414]},
      {stage1_32[317]}
   );
   gpc1_1 gpc3914 (
      {stage0_32[415]},
      {stage1_32[318]}
   );
   gpc1_1 gpc3915 (
      {stage0_32[416]},
      {stage1_32[319]}
   );
   gpc1_1 gpc3916 (
      {stage0_32[417]},
      {stage1_32[320]}
   );
   gpc1_1 gpc3917 (
      {stage0_32[418]},
      {stage1_32[321]}
   );
   gpc1_1 gpc3918 (
      {stage0_32[419]},
      {stage1_32[322]}
   );
   gpc1_1 gpc3919 (
      {stage0_32[420]},
      {stage1_32[323]}
   );
   gpc1_1 gpc3920 (
      {stage0_32[421]},
      {stage1_32[324]}
   );
   gpc1_1 gpc3921 (
      {stage0_32[422]},
      {stage1_32[325]}
   );
   gpc1_1 gpc3922 (
      {stage0_32[423]},
      {stage1_32[326]}
   );
   gpc1_1 gpc3923 (
      {stage0_32[424]},
      {stage1_32[327]}
   );
   gpc1_1 gpc3924 (
      {stage0_32[425]},
      {stage1_32[328]}
   );
   gpc1_1 gpc3925 (
      {stage0_32[426]},
      {stage1_32[329]}
   );
   gpc1_1 gpc3926 (
      {stage0_32[427]},
      {stage1_32[330]}
   );
   gpc1_1 gpc3927 (
      {stage0_32[428]},
      {stage1_32[331]}
   );
   gpc1_1 gpc3928 (
      {stage0_32[429]},
      {stage1_32[332]}
   );
   gpc1_1 gpc3929 (
      {stage0_32[430]},
      {stage1_32[333]}
   );
   gpc1_1 gpc3930 (
      {stage0_32[431]},
      {stage1_32[334]}
   );
   gpc1_1 gpc3931 (
      {stage0_32[432]},
      {stage1_32[335]}
   );
   gpc1_1 gpc3932 (
      {stage0_32[433]},
      {stage1_32[336]}
   );
   gpc1_1 gpc3933 (
      {stage0_32[434]},
      {stage1_32[337]}
   );
   gpc1_1 gpc3934 (
      {stage0_32[435]},
      {stage1_32[338]}
   );
   gpc1_1 gpc3935 (
      {stage0_32[436]},
      {stage1_32[339]}
   );
   gpc1_1 gpc3936 (
      {stage0_32[437]},
      {stage1_32[340]}
   );
   gpc1_1 gpc3937 (
      {stage0_32[438]},
      {stage1_32[341]}
   );
   gpc1_1 gpc3938 (
      {stage0_32[439]},
      {stage1_32[342]}
   );
   gpc1_1 gpc3939 (
      {stage0_32[440]},
      {stage1_32[343]}
   );
   gpc1_1 gpc3940 (
      {stage0_32[441]},
      {stage1_32[344]}
   );
   gpc1_1 gpc3941 (
      {stage0_32[442]},
      {stage1_32[345]}
   );
   gpc1_1 gpc3942 (
      {stage0_32[443]},
      {stage1_32[346]}
   );
   gpc1_1 gpc3943 (
      {stage0_32[444]},
      {stage1_32[347]}
   );
   gpc1_1 gpc3944 (
      {stage0_32[445]},
      {stage1_32[348]}
   );
   gpc1_1 gpc3945 (
      {stage0_32[446]},
      {stage1_32[349]}
   );
   gpc1_1 gpc3946 (
      {stage0_32[447]},
      {stage1_32[350]}
   );
   gpc1_1 gpc3947 (
      {stage0_32[448]},
      {stage1_32[351]}
   );
   gpc1_1 gpc3948 (
      {stage0_32[449]},
      {stage1_32[352]}
   );
   gpc1_1 gpc3949 (
      {stage0_32[450]},
      {stage1_32[353]}
   );
   gpc1_1 gpc3950 (
      {stage0_32[451]},
      {stage1_32[354]}
   );
   gpc1_1 gpc3951 (
      {stage0_32[452]},
      {stage1_32[355]}
   );
   gpc1_1 gpc3952 (
      {stage0_32[453]},
      {stage1_32[356]}
   );
   gpc1_1 gpc3953 (
      {stage0_32[454]},
      {stage1_32[357]}
   );
   gpc1_1 gpc3954 (
      {stage0_32[455]},
      {stage1_32[358]}
   );
   gpc1_1 gpc3955 (
      {stage0_32[456]},
      {stage1_32[359]}
   );
   gpc1_1 gpc3956 (
      {stage0_32[457]},
      {stage1_32[360]}
   );
   gpc1_1 gpc3957 (
      {stage0_32[458]},
      {stage1_32[361]}
   );
   gpc1_1 gpc3958 (
      {stage0_32[459]},
      {stage1_32[362]}
   );
   gpc1_1 gpc3959 (
      {stage0_32[460]},
      {stage1_32[363]}
   );
   gpc1_1 gpc3960 (
      {stage0_32[461]},
      {stage1_32[364]}
   );
   gpc1_1 gpc3961 (
      {stage0_32[462]},
      {stage1_32[365]}
   );
   gpc1_1 gpc3962 (
      {stage0_32[463]},
      {stage1_32[366]}
   );
   gpc1_1 gpc3963 (
      {stage0_32[464]},
      {stage1_32[367]}
   );
   gpc1_1 gpc3964 (
      {stage0_32[465]},
      {stage1_32[368]}
   );
   gpc1_1 gpc3965 (
      {stage0_32[466]},
      {stage1_32[369]}
   );
   gpc1_1 gpc3966 (
      {stage0_32[467]},
      {stage1_32[370]}
   );
   gpc1_1 gpc3967 (
      {stage0_32[468]},
      {stage1_32[371]}
   );
   gpc1_1 gpc3968 (
      {stage0_32[469]},
      {stage1_32[372]}
   );
   gpc1_1 gpc3969 (
      {stage0_32[470]},
      {stage1_32[373]}
   );
   gpc1_1 gpc3970 (
      {stage0_32[471]},
      {stage1_32[374]}
   );
   gpc1_1 gpc3971 (
      {stage0_32[472]},
      {stage1_32[375]}
   );
   gpc1_1 gpc3972 (
      {stage0_32[473]},
      {stage1_32[376]}
   );
   gpc1_1 gpc3973 (
      {stage0_32[474]},
      {stage1_32[377]}
   );
   gpc1_1 gpc3974 (
      {stage0_32[475]},
      {stage1_32[378]}
   );
   gpc1_1 gpc3975 (
      {stage0_32[476]},
      {stage1_32[379]}
   );
   gpc1_1 gpc3976 (
      {stage0_32[477]},
      {stage1_32[380]}
   );
   gpc1_1 gpc3977 (
      {stage0_32[478]},
      {stage1_32[381]}
   );
   gpc1_1 gpc3978 (
      {stage0_32[479]},
      {stage1_32[382]}
   );
   gpc1_1 gpc3979 (
      {stage0_32[480]},
      {stage1_32[383]}
   );
   gpc1_1 gpc3980 (
      {stage0_32[481]},
      {stage1_32[384]}
   );
   gpc1_1 gpc3981 (
      {stage0_32[482]},
      {stage1_32[385]}
   );
   gpc1_1 gpc3982 (
      {stage0_32[483]},
      {stage1_32[386]}
   );
   gpc1_1 gpc3983 (
      {stage0_32[484]},
      {stage1_32[387]}
   );
   gpc1_1 gpc3984 (
      {stage0_32[485]},
      {stage1_32[388]}
   );
   gpc1_1 gpc3985 (
      {stage0_32[486]},
      {stage1_32[389]}
   );
   gpc1_1 gpc3986 (
      {stage0_32[487]},
      {stage1_32[390]}
   );
   gpc1_1 gpc3987 (
      {stage0_32[488]},
      {stage1_32[391]}
   );
   gpc1_1 gpc3988 (
      {stage0_32[489]},
      {stage1_32[392]}
   );
   gpc1_1 gpc3989 (
      {stage0_32[490]},
      {stage1_32[393]}
   );
   gpc1_1 gpc3990 (
      {stage0_32[491]},
      {stage1_32[394]}
   );
   gpc1_1 gpc3991 (
      {stage0_32[492]},
      {stage1_32[395]}
   );
   gpc1_1 gpc3992 (
      {stage0_32[493]},
      {stage1_32[396]}
   );
   gpc1_1 gpc3993 (
      {stage0_32[494]},
      {stage1_32[397]}
   );
   gpc1_1 gpc3994 (
      {stage0_32[495]},
      {stage1_32[398]}
   );
   gpc1_1 gpc3995 (
      {stage0_32[496]},
      {stage1_32[399]}
   );
   gpc1_1 gpc3996 (
      {stage0_32[497]},
      {stage1_32[400]}
   );
   gpc1_1 gpc3997 (
      {stage0_32[498]},
      {stage1_32[401]}
   );
   gpc1_1 gpc3998 (
      {stage0_32[499]},
      {stage1_32[402]}
   );
   gpc1_1 gpc3999 (
      {stage0_32[500]},
      {stage1_32[403]}
   );
   gpc1_1 gpc4000 (
      {stage0_32[501]},
      {stage1_32[404]}
   );
   gpc1_1 gpc4001 (
      {stage0_32[502]},
      {stage1_32[405]}
   );
   gpc1_1 gpc4002 (
      {stage0_32[503]},
      {stage1_32[406]}
   );
   gpc1_1 gpc4003 (
      {stage0_32[504]},
      {stage1_32[407]}
   );
   gpc1_1 gpc4004 (
      {stage0_32[505]},
      {stage1_32[408]}
   );
   gpc1_1 gpc4005 (
      {stage0_32[506]},
      {stage1_32[409]}
   );
   gpc1_1 gpc4006 (
      {stage0_32[507]},
      {stage1_32[410]}
   );
   gpc1_1 gpc4007 (
      {stage0_32[508]},
      {stage1_32[411]}
   );
   gpc1_1 gpc4008 (
      {stage0_32[509]},
      {stage1_32[412]}
   );
   gpc1_1 gpc4009 (
      {stage0_32[510]},
      {stage1_32[413]}
   );
   gpc1_1 gpc4010 (
      {stage0_32[511]},
      {stage1_32[414]}
   );
   gpc1_1 gpc4011 (
      {stage0_33[491]},
      {stage1_33[189]}
   );
   gpc1_1 gpc4012 (
      {stage0_33[492]},
      {stage1_33[190]}
   );
   gpc1_1 gpc4013 (
      {stage0_33[493]},
      {stage1_33[191]}
   );
   gpc1_1 gpc4014 (
      {stage0_33[494]},
      {stage1_33[192]}
   );
   gpc1_1 gpc4015 (
      {stage0_33[495]},
      {stage1_33[193]}
   );
   gpc1_1 gpc4016 (
      {stage0_33[496]},
      {stage1_33[194]}
   );
   gpc1_1 gpc4017 (
      {stage0_33[497]},
      {stage1_33[195]}
   );
   gpc1_1 gpc4018 (
      {stage0_33[498]},
      {stage1_33[196]}
   );
   gpc1_1 gpc4019 (
      {stage0_33[499]},
      {stage1_33[197]}
   );
   gpc1_1 gpc4020 (
      {stage0_33[500]},
      {stage1_33[198]}
   );
   gpc1_1 gpc4021 (
      {stage0_33[501]},
      {stage1_33[199]}
   );
   gpc1_1 gpc4022 (
      {stage0_33[502]},
      {stage1_33[200]}
   );
   gpc1_1 gpc4023 (
      {stage0_33[503]},
      {stage1_33[201]}
   );
   gpc1_1 gpc4024 (
      {stage0_33[504]},
      {stage1_33[202]}
   );
   gpc1_1 gpc4025 (
      {stage0_33[505]},
      {stage1_33[203]}
   );
   gpc1_1 gpc4026 (
      {stage0_33[506]},
      {stage1_33[204]}
   );
   gpc1_1 gpc4027 (
      {stage0_33[507]},
      {stage1_33[205]}
   );
   gpc1_1 gpc4028 (
      {stage0_33[508]},
      {stage1_33[206]}
   );
   gpc1_1 gpc4029 (
      {stage0_33[509]},
      {stage1_33[207]}
   );
   gpc1_1 gpc4030 (
      {stage0_33[510]},
      {stage1_33[208]}
   );
   gpc1_1 gpc4031 (
      {stage0_33[511]},
      {stage1_33[209]}
   );
   gpc1_1 gpc4032 (
      {stage0_34[396]},
      {stage1_34[152]}
   );
   gpc1_1 gpc4033 (
      {stage0_34[397]},
      {stage1_34[153]}
   );
   gpc1_1 gpc4034 (
      {stage0_34[398]},
      {stage1_34[154]}
   );
   gpc1_1 gpc4035 (
      {stage0_34[399]},
      {stage1_34[155]}
   );
   gpc1_1 gpc4036 (
      {stage0_34[400]},
      {stage1_34[156]}
   );
   gpc1_1 gpc4037 (
      {stage0_34[401]},
      {stage1_34[157]}
   );
   gpc1_1 gpc4038 (
      {stage0_34[402]},
      {stage1_34[158]}
   );
   gpc1_1 gpc4039 (
      {stage0_34[403]},
      {stage1_34[159]}
   );
   gpc1_1 gpc4040 (
      {stage0_34[404]},
      {stage1_34[160]}
   );
   gpc1_1 gpc4041 (
      {stage0_34[405]},
      {stage1_34[161]}
   );
   gpc1_1 gpc4042 (
      {stage0_34[406]},
      {stage1_34[162]}
   );
   gpc1_1 gpc4043 (
      {stage0_34[407]},
      {stage1_34[163]}
   );
   gpc1_1 gpc4044 (
      {stage0_34[408]},
      {stage1_34[164]}
   );
   gpc1_1 gpc4045 (
      {stage0_34[409]},
      {stage1_34[165]}
   );
   gpc1_1 gpc4046 (
      {stage0_34[410]},
      {stage1_34[166]}
   );
   gpc1_1 gpc4047 (
      {stage0_34[411]},
      {stage1_34[167]}
   );
   gpc1_1 gpc4048 (
      {stage0_34[412]},
      {stage1_34[168]}
   );
   gpc1_1 gpc4049 (
      {stage0_34[413]},
      {stage1_34[169]}
   );
   gpc1_1 gpc4050 (
      {stage0_34[414]},
      {stage1_34[170]}
   );
   gpc1_1 gpc4051 (
      {stage0_34[415]},
      {stage1_34[171]}
   );
   gpc1_1 gpc4052 (
      {stage0_34[416]},
      {stage1_34[172]}
   );
   gpc1_1 gpc4053 (
      {stage0_34[417]},
      {stage1_34[173]}
   );
   gpc1_1 gpc4054 (
      {stage0_34[418]},
      {stage1_34[174]}
   );
   gpc1_1 gpc4055 (
      {stage0_34[419]},
      {stage1_34[175]}
   );
   gpc1_1 gpc4056 (
      {stage0_34[420]},
      {stage1_34[176]}
   );
   gpc1_1 gpc4057 (
      {stage0_34[421]},
      {stage1_34[177]}
   );
   gpc1_1 gpc4058 (
      {stage0_34[422]},
      {stage1_34[178]}
   );
   gpc1_1 gpc4059 (
      {stage0_34[423]},
      {stage1_34[179]}
   );
   gpc1_1 gpc4060 (
      {stage0_34[424]},
      {stage1_34[180]}
   );
   gpc1_1 gpc4061 (
      {stage0_34[425]},
      {stage1_34[181]}
   );
   gpc1_1 gpc4062 (
      {stage0_34[426]},
      {stage1_34[182]}
   );
   gpc1_1 gpc4063 (
      {stage0_34[427]},
      {stage1_34[183]}
   );
   gpc1_1 gpc4064 (
      {stage0_34[428]},
      {stage1_34[184]}
   );
   gpc1_1 gpc4065 (
      {stage0_34[429]},
      {stage1_34[185]}
   );
   gpc1_1 gpc4066 (
      {stage0_34[430]},
      {stage1_34[186]}
   );
   gpc1_1 gpc4067 (
      {stage0_34[431]},
      {stage1_34[187]}
   );
   gpc1_1 gpc4068 (
      {stage0_34[432]},
      {stage1_34[188]}
   );
   gpc1_1 gpc4069 (
      {stage0_34[433]},
      {stage1_34[189]}
   );
   gpc1_1 gpc4070 (
      {stage0_34[434]},
      {stage1_34[190]}
   );
   gpc1_1 gpc4071 (
      {stage0_34[435]},
      {stage1_34[191]}
   );
   gpc1_1 gpc4072 (
      {stage0_34[436]},
      {stage1_34[192]}
   );
   gpc1_1 gpc4073 (
      {stage0_34[437]},
      {stage1_34[193]}
   );
   gpc1_1 gpc4074 (
      {stage0_34[438]},
      {stage1_34[194]}
   );
   gpc1_1 gpc4075 (
      {stage0_34[439]},
      {stage1_34[195]}
   );
   gpc1_1 gpc4076 (
      {stage0_34[440]},
      {stage1_34[196]}
   );
   gpc1_1 gpc4077 (
      {stage0_34[441]},
      {stage1_34[197]}
   );
   gpc1_1 gpc4078 (
      {stage0_34[442]},
      {stage1_34[198]}
   );
   gpc1_1 gpc4079 (
      {stage0_34[443]},
      {stage1_34[199]}
   );
   gpc1_1 gpc4080 (
      {stage0_34[444]},
      {stage1_34[200]}
   );
   gpc1_1 gpc4081 (
      {stage0_34[445]},
      {stage1_34[201]}
   );
   gpc1_1 gpc4082 (
      {stage0_34[446]},
      {stage1_34[202]}
   );
   gpc1_1 gpc4083 (
      {stage0_34[447]},
      {stage1_34[203]}
   );
   gpc1_1 gpc4084 (
      {stage0_34[448]},
      {stage1_34[204]}
   );
   gpc1_1 gpc4085 (
      {stage0_34[449]},
      {stage1_34[205]}
   );
   gpc1_1 gpc4086 (
      {stage0_34[450]},
      {stage1_34[206]}
   );
   gpc1_1 gpc4087 (
      {stage0_34[451]},
      {stage1_34[207]}
   );
   gpc1_1 gpc4088 (
      {stage0_34[452]},
      {stage1_34[208]}
   );
   gpc1_1 gpc4089 (
      {stage0_34[453]},
      {stage1_34[209]}
   );
   gpc1_1 gpc4090 (
      {stage0_34[454]},
      {stage1_34[210]}
   );
   gpc1_1 gpc4091 (
      {stage0_34[455]},
      {stage1_34[211]}
   );
   gpc1_1 gpc4092 (
      {stage0_34[456]},
      {stage1_34[212]}
   );
   gpc1_1 gpc4093 (
      {stage0_34[457]},
      {stage1_34[213]}
   );
   gpc1_1 gpc4094 (
      {stage0_34[458]},
      {stage1_34[214]}
   );
   gpc1_1 gpc4095 (
      {stage0_34[459]},
      {stage1_34[215]}
   );
   gpc1_1 gpc4096 (
      {stage0_34[460]},
      {stage1_34[216]}
   );
   gpc1_1 gpc4097 (
      {stage0_34[461]},
      {stage1_34[217]}
   );
   gpc1_1 gpc4098 (
      {stage0_34[462]},
      {stage1_34[218]}
   );
   gpc1_1 gpc4099 (
      {stage0_34[463]},
      {stage1_34[219]}
   );
   gpc1_1 gpc4100 (
      {stage0_34[464]},
      {stage1_34[220]}
   );
   gpc1_1 gpc4101 (
      {stage0_34[465]},
      {stage1_34[221]}
   );
   gpc1_1 gpc4102 (
      {stage0_34[466]},
      {stage1_34[222]}
   );
   gpc1_1 gpc4103 (
      {stage0_34[467]},
      {stage1_34[223]}
   );
   gpc1_1 gpc4104 (
      {stage0_34[468]},
      {stage1_34[224]}
   );
   gpc1_1 gpc4105 (
      {stage0_34[469]},
      {stage1_34[225]}
   );
   gpc1_1 gpc4106 (
      {stage0_34[470]},
      {stage1_34[226]}
   );
   gpc1_1 gpc4107 (
      {stage0_34[471]},
      {stage1_34[227]}
   );
   gpc1_1 gpc4108 (
      {stage0_34[472]},
      {stage1_34[228]}
   );
   gpc1_1 gpc4109 (
      {stage0_34[473]},
      {stage1_34[229]}
   );
   gpc1_1 gpc4110 (
      {stage0_34[474]},
      {stage1_34[230]}
   );
   gpc1_1 gpc4111 (
      {stage0_34[475]},
      {stage1_34[231]}
   );
   gpc1_1 gpc4112 (
      {stage0_34[476]},
      {stage1_34[232]}
   );
   gpc1_1 gpc4113 (
      {stage0_34[477]},
      {stage1_34[233]}
   );
   gpc1_1 gpc4114 (
      {stage0_34[478]},
      {stage1_34[234]}
   );
   gpc1_1 gpc4115 (
      {stage0_34[479]},
      {stage1_34[235]}
   );
   gpc1_1 gpc4116 (
      {stage0_34[480]},
      {stage1_34[236]}
   );
   gpc1_1 gpc4117 (
      {stage0_34[481]},
      {stage1_34[237]}
   );
   gpc1_1 gpc4118 (
      {stage0_34[482]},
      {stage1_34[238]}
   );
   gpc1_1 gpc4119 (
      {stage0_34[483]},
      {stage1_34[239]}
   );
   gpc1_1 gpc4120 (
      {stage0_34[484]},
      {stage1_34[240]}
   );
   gpc1_1 gpc4121 (
      {stage0_34[485]},
      {stage1_34[241]}
   );
   gpc1_1 gpc4122 (
      {stage0_34[486]},
      {stage1_34[242]}
   );
   gpc1_1 gpc4123 (
      {stage0_34[487]},
      {stage1_34[243]}
   );
   gpc1_1 gpc4124 (
      {stage0_34[488]},
      {stage1_34[244]}
   );
   gpc1_1 gpc4125 (
      {stage0_34[489]},
      {stage1_34[245]}
   );
   gpc1_1 gpc4126 (
      {stage0_34[490]},
      {stage1_34[246]}
   );
   gpc1_1 gpc4127 (
      {stage0_34[491]},
      {stage1_34[247]}
   );
   gpc1_1 gpc4128 (
      {stage0_34[492]},
      {stage1_34[248]}
   );
   gpc1_1 gpc4129 (
      {stage0_34[493]},
      {stage1_34[249]}
   );
   gpc1_1 gpc4130 (
      {stage0_34[494]},
      {stage1_34[250]}
   );
   gpc1_1 gpc4131 (
      {stage0_34[495]},
      {stage1_34[251]}
   );
   gpc1_1 gpc4132 (
      {stage0_34[496]},
      {stage1_34[252]}
   );
   gpc1_1 gpc4133 (
      {stage0_34[497]},
      {stage1_34[253]}
   );
   gpc1_1 gpc4134 (
      {stage0_34[498]},
      {stage1_34[254]}
   );
   gpc1_1 gpc4135 (
      {stage0_34[499]},
      {stage1_34[255]}
   );
   gpc1_1 gpc4136 (
      {stage0_34[500]},
      {stage1_34[256]}
   );
   gpc1_1 gpc4137 (
      {stage0_34[501]},
      {stage1_34[257]}
   );
   gpc1_1 gpc4138 (
      {stage0_34[502]},
      {stage1_34[258]}
   );
   gpc1_1 gpc4139 (
      {stage0_34[503]},
      {stage1_34[259]}
   );
   gpc1_1 gpc4140 (
      {stage0_34[504]},
      {stage1_34[260]}
   );
   gpc1_1 gpc4141 (
      {stage0_34[505]},
      {stage1_34[261]}
   );
   gpc1_1 gpc4142 (
      {stage0_34[506]},
      {stage1_34[262]}
   );
   gpc1_1 gpc4143 (
      {stage0_34[507]},
      {stage1_34[263]}
   );
   gpc1_1 gpc4144 (
      {stage0_34[508]},
      {stage1_34[264]}
   );
   gpc1_1 gpc4145 (
      {stage0_34[509]},
      {stage1_34[265]}
   );
   gpc1_1 gpc4146 (
      {stage0_34[510]},
      {stage1_34[266]}
   );
   gpc1_1 gpc4147 (
      {stage0_34[511]},
      {stage1_34[267]}
   );
   gpc1_1 gpc4148 (
      {stage0_35[495]},
      {stage1_35[174]}
   );
   gpc1_1 gpc4149 (
      {stage0_35[496]},
      {stage1_35[175]}
   );
   gpc1_1 gpc4150 (
      {stage0_35[497]},
      {stage1_35[176]}
   );
   gpc1_1 gpc4151 (
      {stage0_35[498]},
      {stage1_35[177]}
   );
   gpc1_1 gpc4152 (
      {stage0_35[499]},
      {stage1_35[178]}
   );
   gpc1_1 gpc4153 (
      {stage0_35[500]},
      {stage1_35[179]}
   );
   gpc1_1 gpc4154 (
      {stage0_35[501]},
      {stage1_35[180]}
   );
   gpc1_1 gpc4155 (
      {stage0_35[502]},
      {stage1_35[181]}
   );
   gpc1_1 gpc4156 (
      {stage0_35[503]},
      {stage1_35[182]}
   );
   gpc1_1 gpc4157 (
      {stage0_35[504]},
      {stage1_35[183]}
   );
   gpc1_1 gpc4158 (
      {stage0_35[505]},
      {stage1_35[184]}
   );
   gpc1_1 gpc4159 (
      {stage0_35[506]},
      {stage1_35[185]}
   );
   gpc1_1 gpc4160 (
      {stage0_35[507]},
      {stage1_35[186]}
   );
   gpc1_1 gpc4161 (
      {stage0_35[508]},
      {stage1_35[187]}
   );
   gpc1_1 gpc4162 (
      {stage0_35[509]},
      {stage1_35[188]}
   );
   gpc1_1 gpc4163 (
      {stage0_35[510]},
      {stage1_35[189]}
   );
   gpc1_1 gpc4164 (
      {stage0_35[511]},
      {stage1_35[190]}
   );
   gpc1_1 gpc4165 (
      {stage0_36[367]},
      {stage1_36[186]}
   );
   gpc1_1 gpc4166 (
      {stage0_36[368]},
      {stage1_36[187]}
   );
   gpc1_1 gpc4167 (
      {stage0_36[369]},
      {stage1_36[188]}
   );
   gpc1_1 gpc4168 (
      {stage0_36[370]},
      {stage1_36[189]}
   );
   gpc1_1 gpc4169 (
      {stage0_36[371]},
      {stage1_36[190]}
   );
   gpc1_1 gpc4170 (
      {stage0_36[372]},
      {stage1_36[191]}
   );
   gpc1_1 gpc4171 (
      {stage0_36[373]},
      {stage1_36[192]}
   );
   gpc1_1 gpc4172 (
      {stage0_36[374]},
      {stage1_36[193]}
   );
   gpc1_1 gpc4173 (
      {stage0_36[375]},
      {stage1_36[194]}
   );
   gpc1_1 gpc4174 (
      {stage0_36[376]},
      {stage1_36[195]}
   );
   gpc1_1 gpc4175 (
      {stage0_36[377]},
      {stage1_36[196]}
   );
   gpc1_1 gpc4176 (
      {stage0_36[378]},
      {stage1_36[197]}
   );
   gpc1_1 gpc4177 (
      {stage0_36[379]},
      {stage1_36[198]}
   );
   gpc1_1 gpc4178 (
      {stage0_36[380]},
      {stage1_36[199]}
   );
   gpc1_1 gpc4179 (
      {stage0_36[381]},
      {stage1_36[200]}
   );
   gpc1_1 gpc4180 (
      {stage0_36[382]},
      {stage1_36[201]}
   );
   gpc1_1 gpc4181 (
      {stage0_36[383]},
      {stage1_36[202]}
   );
   gpc1_1 gpc4182 (
      {stage0_36[384]},
      {stage1_36[203]}
   );
   gpc1_1 gpc4183 (
      {stage0_36[385]},
      {stage1_36[204]}
   );
   gpc1_1 gpc4184 (
      {stage0_36[386]},
      {stage1_36[205]}
   );
   gpc1_1 gpc4185 (
      {stage0_36[387]},
      {stage1_36[206]}
   );
   gpc1_1 gpc4186 (
      {stage0_36[388]},
      {stage1_36[207]}
   );
   gpc1_1 gpc4187 (
      {stage0_36[389]},
      {stage1_36[208]}
   );
   gpc1_1 gpc4188 (
      {stage0_36[390]},
      {stage1_36[209]}
   );
   gpc1_1 gpc4189 (
      {stage0_36[391]},
      {stage1_36[210]}
   );
   gpc1_1 gpc4190 (
      {stage0_36[392]},
      {stage1_36[211]}
   );
   gpc1_1 gpc4191 (
      {stage0_36[393]},
      {stage1_36[212]}
   );
   gpc1_1 gpc4192 (
      {stage0_36[394]},
      {stage1_36[213]}
   );
   gpc1_1 gpc4193 (
      {stage0_36[395]},
      {stage1_36[214]}
   );
   gpc1_1 gpc4194 (
      {stage0_36[396]},
      {stage1_36[215]}
   );
   gpc1_1 gpc4195 (
      {stage0_36[397]},
      {stage1_36[216]}
   );
   gpc1_1 gpc4196 (
      {stage0_36[398]},
      {stage1_36[217]}
   );
   gpc1_1 gpc4197 (
      {stage0_36[399]},
      {stage1_36[218]}
   );
   gpc1_1 gpc4198 (
      {stage0_36[400]},
      {stage1_36[219]}
   );
   gpc1_1 gpc4199 (
      {stage0_36[401]},
      {stage1_36[220]}
   );
   gpc1_1 gpc4200 (
      {stage0_36[402]},
      {stage1_36[221]}
   );
   gpc1_1 gpc4201 (
      {stage0_36[403]},
      {stage1_36[222]}
   );
   gpc1_1 gpc4202 (
      {stage0_36[404]},
      {stage1_36[223]}
   );
   gpc1_1 gpc4203 (
      {stage0_36[405]},
      {stage1_36[224]}
   );
   gpc1_1 gpc4204 (
      {stage0_36[406]},
      {stage1_36[225]}
   );
   gpc1_1 gpc4205 (
      {stage0_36[407]},
      {stage1_36[226]}
   );
   gpc1_1 gpc4206 (
      {stage0_36[408]},
      {stage1_36[227]}
   );
   gpc1_1 gpc4207 (
      {stage0_36[409]},
      {stage1_36[228]}
   );
   gpc1_1 gpc4208 (
      {stage0_36[410]},
      {stage1_36[229]}
   );
   gpc1_1 gpc4209 (
      {stage0_36[411]},
      {stage1_36[230]}
   );
   gpc1_1 gpc4210 (
      {stage0_36[412]},
      {stage1_36[231]}
   );
   gpc1_1 gpc4211 (
      {stage0_36[413]},
      {stage1_36[232]}
   );
   gpc1_1 gpc4212 (
      {stage0_36[414]},
      {stage1_36[233]}
   );
   gpc1_1 gpc4213 (
      {stage0_36[415]},
      {stage1_36[234]}
   );
   gpc1_1 gpc4214 (
      {stage0_36[416]},
      {stage1_36[235]}
   );
   gpc1_1 gpc4215 (
      {stage0_36[417]},
      {stage1_36[236]}
   );
   gpc1_1 gpc4216 (
      {stage0_36[418]},
      {stage1_36[237]}
   );
   gpc1_1 gpc4217 (
      {stage0_36[419]},
      {stage1_36[238]}
   );
   gpc1_1 gpc4218 (
      {stage0_36[420]},
      {stage1_36[239]}
   );
   gpc1_1 gpc4219 (
      {stage0_36[421]},
      {stage1_36[240]}
   );
   gpc1_1 gpc4220 (
      {stage0_36[422]},
      {stage1_36[241]}
   );
   gpc1_1 gpc4221 (
      {stage0_36[423]},
      {stage1_36[242]}
   );
   gpc1_1 gpc4222 (
      {stage0_36[424]},
      {stage1_36[243]}
   );
   gpc1_1 gpc4223 (
      {stage0_36[425]},
      {stage1_36[244]}
   );
   gpc1_1 gpc4224 (
      {stage0_36[426]},
      {stage1_36[245]}
   );
   gpc1_1 gpc4225 (
      {stage0_36[427]},
      {stage1_36[246]}
   );
   gpc1_1 gpc4226 (
      {stage0_36[428]},
      {stage1_36[247]}
   );
   gpc1_1 gpc4227 (
      {stage0_36[429]},
      {stage1_36[248]}
   );
   gpc1_1 gpc4228 (
      {stage0_36[430]},
      {stage1_36[249]}
   );
   gpc1_1 gpc4229 (
      {stage0_36[431]},
      {stage1_36[250]}
   );
   gpc1_1 gpc4230 (
      {stage0_36[432]},
      {stage1_36[251]}
   );
   gpc1_1 gpc4231 (
      {stage0_36[433]},
      {stage1_36[252]}
   );
   gpc1_1 gpc4232 (
      {stage0_36[434]},
      {stage1_36[253]}
   );
   gpc1_1 gpc4233 (
      {stage0_36[435]},
      {stage1_36[254]}
   );
   gpc1_1 gpc4234 (
      {stage0_36[436]},
      {stage1_36[255]}
   );
   gpc1_1 gpc4235 (
      {stage0_36[437]},
      {stage1_36[256]}
   );
   gpc1_1 gpc4236 (
      {stage0_36[438]},
      {stage1_36[257]}
   );
   gpc1_1 gpc4237 (
      {stage0_36[439]},
      {stage1_36[258]}
   );
   gpc1_1 gpc4238 (
      {stage0_36[440]},
      {stage1_36[259]}
   );
   gpc1_1 gpc4239 (
      {stage0_36[441]},
      {stage1_36[260]}
   );
   gpc1_1 gpc4240 (
      {stage0_36[442]},
      {stage1_36[261]}
   );
   gpc1_1 gpc4241 (
      {stage0_36[443]},
      {stage1_36[262]}
   );
   gpc1_1 gpc4242 (
      {stage0_36[444]},
      {stage1_36[263]}
   );
   gpc1_1 gpc4243 (
      {stage0_36[445]},
      {stage1_36[264]}
   );
   gpc1_1 gpc4244 (
      {stage0_36[446]},
      {stage1_36[265]}
   );
   gpc1_1 gpc4245 (
      {stage0_36[447]},
      {stage1_36[266]}
   );
   gpc1_1 gpc4246 (
      {stage0_36[448]},
      {stage1_36[267]}
   );
   gpc1_1 gpc4247 (
      {stage0_36[449]},
      {stage1_36[268]}
   );
   gpc1_1 gpc4248 (
      {stage0_36[450]},
      {stage1_36[269]}
   );
   gpc1_1 gpc4249 (
      {stage0_36[451]},
      {stage1_36[270]}
   );
   gpc1_1 gpc4250 (
      {stage0_36[452]},
      {stage1_36[271]}
   );
   gpc1_1 gpc4251 (
      {stage0_36[453]},
      {stage1_36[272]}
   );
   gpc1_1 gpc4252 (
      {stage0_36[454]},
      {stage1_36[273]}
   );
   gpc1_1 gpc4253 (
      {stage0_36[455]},
      {stage1_36[274]}
   );
   gpc1_1 gpc4254 (
      {stage0_36[456]},
      {stage1_36[275]}
   );
   gpc1_1 gpc4255 (
      {stage0_36[457]},
      {stage1_36[276]}
   );
   gpc1_1 gpc4256 (
      {stage0_36[458]},
      {stage1_36[277]}
   );
   gpc1_1 gpc4257 (
      {stage0_36[459]},
      {stage1_36[278]}
   );
   gpc1_1 gpc4258 (
      {stage0_36[460]},
      {stage1_36[279]}
   );
   gpc1_1 gpc4259 (
      {stage0_36[461]},
      {stage1_36[280]}
   );
   gpc1_1 gpc4260 (
      {stage0_36[462]},
      {stage1_36[281]}
   );
   gpc1_1 gpc4261 (
      {stage0_36[463]},
      {stage1_36[282]}
   );
   gpc1_1 gpc4262 (
      {stage0_36[464]},
      {stage1_36[283]}
   );
   gpc1_1 gpc4263 (
      {stage0_36[465]},
      {stage1_36[284]}
   );
   gpc1_1 gpc4264 (
      {stage0_36[466]},
      {stage1_36[285]}
   );
   gpc1_1 gpc4265 (
      {stage0_36[467]},
      {stage1_36[286]}
   );
   gpc1_1 gpc4266 (
      {stage0_36[468]},
      {stage1_36[287]}
   );
   gpc1_1 gpc4267 (
      {stage0_36[469]},
      {stage1_36[288]}
   );
   gpc1_1 gpc4268 (
      {stage0_36[470]},
      {stage1_36[289]}
   );
   gpc1_1 gpc4269 (
      {stage0_36[471]},
      {stage1_36[290]}
   );
   gpc1_1 gpc4270 (
      {stage0_36[472]},
      {stage1_36[291]}
   );
   gpc1_1 gpc4271 (
      {stage0_36[473]},
      {stage1_36[292]}
   );
   gpc1_1 gpc4272 (
      {stage0_36[474]},
      {stage1_36[293]}
   );
   gpc1_1 gpc4273 (
      {stage0_36[475]},
      {stage1_36[294]}
   );
   gpc1_1 gpc4274 (
      {stage0_36[476]},
      {stage1_36[295]}
   );
   gpc1_1 gpc4275 (
      {stage0_36[477]},
      {stage1_36[296]}
   );
   gpc1_1 gpc4276 (
      {stage0_36[478]},
      {stage1_36[297]}
   );
   gpc1_1 gpc4277 (
      {stage0_36[479]},
      {stage1_36[298]}
   );
   gpc1_1 gpc4278 (
      {stage0_36[480]},
      {stage1_36[299]}
   );
   gpc1_1 gpc4279 (
      {stage0_36[481]},
      {stage1_36[300]}
   );
   gpc1_1 gpc4280 (
      {stage0_36[482]},
      {stage1_36[301]}
   );
   gpc1_1 gpc4281 (
      {stage0_36[483]},
      {stage1_36[302]}
   );
   gpc1_1 gpc4282 (
      {stage0_36[484]},
      {stage1_36[303]}
   );
   gpc1_1 gpc4283 (
      {stage0_36[485]},
      {stage1_36[304]}
   );
   gpc1_1 gpc4284 (
      {stage0_36[486]},
      {stage1_36[305]}
   );
   gpc1_1 gpc4285 (
      {stage0_36[487]},
      {stage1_36[306]}
   );
   gpc1_1 gpc4286 (
      {stage0_36[488]},
      {stage1_36[307]}
   );
   gpc1_1 gpc4287 (
      {stage0_36[489]},
      {stage1_36[308]}
   );
   gpc1_1 gpc4288 (
      {stage0_36[490]},
      {stage1_36[309]}
   );
   gpc1_1 gpc4289 (
      {stage0_36[491]},
      {stage1_36[310]}
   );
   gpc1_1 gpc4290 (
      {stage0_36[492]},
      {stage1_36[311]}
   );
   gpc1_1 gpc4291 (
      {stage0_36[493]},
      {stage1_36[312]}
   );
   gpc1_1 gpc4292 (
      {stage0_36[494]},
      {stage1_36[313]}
   );
   gpc1_1 gpc4293 (
      {stage0_36[495]},
      {stage1_36[314]}
   );
   gpc1_1 gpc4294 (
      {stage0_36[496]},
      {stage1_36[315]}
   );
   gpc1_1 gpc4295 (
      {stage0_36[497]},
      {stage1_36[316]}
   );
   gpc1_1 gpc4296 (
      {stage0_36[498]},
      {stage1_36[317]}
   );
   gpc1_1 gpc4297 (
      {stage0_36[499]},
      {stage1_36[318]}
   );
   gpc1_1 gpc4298 (
      {stage0_36[500]},
      {stage1_36[319]}
   );
   gpc1_1 gpc4299 (
      {stage0_36[501]},
      {stage1_36[320]}
   );
   gpc1_1 gpc4300 (
      {stage0_36[502]},
      {stage1_36[321]}
   );
   gpc1_1 gpc4301 (
      {stage0_36[503]},
      {stage1_36[322]}
   );
   gpc1_1 gpc4302 (
      {stage0_36[504]},
      {stage1_36[323]}
   );
   gpc1_1 gpc4303 (
      {stage0_36[505]},
      {stage1_36[324]}
   );
   gpc1_1 gpc4304 (
      {stage0_36[506]},
      {stage1_36[325]}
   );
   gpc1_1 gpc4305 (
      {stage0_36[507]},
      {stage1_36[326]}
   );
   gpc1_1 gpc4306 (
      {stage0_36[508]},
      {stage1_36[327]}
   );
   gpc1_1 gpc4307 (
      {stage0_36[509]},
      {stage1_36[328]}
   );
   gpc1_1 gpc4308 (
      {stage0_36[510]},
      {stage1_36[329]}
   );
   gpc1_1 gpc4309 (
      {stage0_36[511]},
      {stage1_36[330]}
   );
   gpc1_1 gpc4310 (
      {stage0_37[392]},
      {stage1_37[183]}
   );
   gpc1_1 gpc4311 (
      {stage0_37[393]},
      {stage1_37[184]}
   );
   gpc1_1 gpc4312 (
      {stage0_37[394]},
      {stage1_37[185]}
   );
   gpc1_1 gpc4313 (
      {stage0_37[395]},
      {stage1_37[186]}
   );
   gpc1_1 gpc4314 (
      {stage0_37[396]},
      {stage1_37[187]}
   );
   gpc1_1 gpc4315 (
      {stage0_37[397]},
      {stage1_37[188]}
   );
   gpc1_1 gpc4316 (
      {stage0_37[398]},
      {stage1_37[189]}
   );
   gpc1_1 gpc4317 (
      {stage0_37[399]},
      {stage1_37[190]}
   );
   gpc1_1 gpc4318 (
      {stage0_37[400]},
      {stage1_37[191]}
   );
   gpc1_1 gpc4319 (
      {stage0_37[401]},
      {stage1_37[192]}
   );
   gpc1_1 gpc4320 (
      {stage0_37[402]},
      {stage1_37[193]}
   );
   gpc1_1 gpc4321 (
      {stage0_37[403]},
      {stage1_37[194]}
   );
   gpc1_1 gpc4322 (
      {stage0_37[404]},
      {stage1_37[195]}
   );
   gpc1_1 gpc4323 (
      {stage0_37[405]},
      {stage1_37[196]}
   );
   gpc1_1 gpc4324 (
      {stage0_37[406]},
      {stage1_37[197]}
   );
   gpc1_1 gpc4325 (
      {stage0_37[407]},
      {stage1_37[198]}
   );
   gpc1_1 gpc4326 (
      {stage0_37[408]},
      {stage1_37[199]}
   );
   gpc1_1 gpc4327 (
      {stage0_37[409]},
      {stage1_37[200]}
   );
   gpc1_1 gpc4328 (
      {stage0_37[410]},
      {stage1_37[201]}
   );
   gpc1_1 gpc4329 (
      {stage0_37[411]},
      {stage1_37[202]}
   );
   gpc1_1 gpc4330 (
      {stage0_37[412]},
      {stage1_37[203]}
   );
   gpc1_1 gpc4331 (
      {stage0_37[413]},
      {stage1_37[204]}
   );
   gpc1_1 gpc4332 (
      {stage0_37[414]},
      {stage1_37[205]}
   );
   gpc1_1 gpc4333 (
      {stage0_37[415]},
      {stage1_37[206]}
   );
   gpc1_1 gpc4334 (
      {stage0_37[416]},
      {stage1_37[207]}
   );
   gpc1_1 gpc4335 (
      {stage0_37[417]},
      {stage1_37[208]}
   );
   gpc1_1 gpc4336 (
      {stage0_37[418]},
      {stage1_37[209]}
   );
   gpc1_1 gpc4337 (
      {stage0_37[419]},
      {stage1_37[210]}
   );
   gpc1_1 gpc4338 (
      {stage0_37[420]},
      {stage1_37[211]}
   );
   gpc1_1 gpc4339 (
      {stage0_37[421]},
      {stage1_37[212]}
   );
   gpc1_1 gpc4340 (
      {stage0_37[422]},
      {stage1_37[213]}
   );
   gpc1_1 gpc4341 (
      {stage0_37[423]},
      {stage1_37[214]}
   );
   gpc1_1 gpc4342 (
      {stage0_37[424]},
      {stage1_37[215]}
   );
   gpc1_1 gpc4343 (
      {stage0_37[425]},
      {stage1_37[216]}
   );
   gpc1_1 gpc4344 (
      {stage0_37[426]},
      {stage1_37[217]}
   );
   gpc1_1 gpc4345 (
      {stage0_37[427]},
      {stage1_37[218]}
   );
   gpc1_1 gpc4346 (
      {stage0_37[428]},
      {stage1_37[219]}
   );
   gpc1_1 gpc4347 (
      {stage0_37[429]},
      {stage1_37[220]}
   );
   gpc1_1 gpc4348 (
      {stage0_37[430]},
      {stage1_37[221]}
   );
   gpc1_1 gpc4349 (
      {stage0_37[431]},
      {stage1_37[222]}
   );
   gpc1_1 gpc4350 (
      {stage0_37[432]},
      {stage1_37[223]}
   );
   gpc1_1 gpc4351 (
      {stage0_37[433]},
      {stage1_37[224]}
   );
   gpc1_1 gpc4352 (
      {stage0_37[434]},
      {stage1_37[225]}
   );
   gpc1_1 gpc4353 (
      {stage0_37[435]},
      {stage1_37[226]}
   );
   gpc1_1 gpc4354 (
      {stage0_37[436]},
      {stage1_37[227]}
   );
   gpc1_1 gpc4355 (
      {stage0_37[437]},
      {stage1_37[228]}
   );
   gpc1_1 gpc4356 (
      {stage0_37[438]},
      {stage1_37[229]}
   );
   gpc1_1 gpc4357 (
      {stage0_37[439]},
      {stage1_37[230]}
   );
   gpc1_1 gpc4358 (
      {stage0_37[440]},
      {stage1_37[231]}
   );
   gpc1_1 gpc4359 (
      {stage0_37[441]},
      {stage1_37[232]}
   );
   gpc1_1 gpc4360 (
      {stage0_37[442]},
      {stage1_37[233]}
   );
   gpc1_1 gpc4361 (
      {stage0_37[443]},
      {stage1_37[234]}
   );
   gpc1_1 gpc4362 (
      {stage0_37[444]},
      {stage1_37[235]}
   );
   gpc1_1 gpc4363 (
      {stage0_37[445]},
      {stage1_37[236]}
   );
   gpc1_1 gpc4364 (
      {stage0_37[446]},
      {stage1_37[237]}
   );
   gpc1_1 gpc4365 (
      {stage0_37[447]},
      {stage1_37[238]}
   );
   gpc1_1 gpc4366 (
      {stage0_37[448]},
      {stage1_37[239]}
   );
   gpc1_1 gpc4367 (
      {stage0_37[449]},
      {stage1_37[240]}
   );
   gpc1_1 gpc4368 (
      {stage0_37[450]},
      {stage1_37[241]}
   );
   gpc1_1 gpc4369 (
      {stage0_37[451]},
      {stage1_37[242]}
   );
   gpc1_1 gpc4370 (
      {stage0_37[452]},
      {stage1_37[243]}
   );
   gpc1_1 gpc4371 (
      {stage0_37[453]},
      {stage1_37[244]}
   );
   gpc1_1 gpc4372 (
      {stage0_37[454]},
      {stage1_37[245]}
   );
   gpc1_1 gpc4373 (
      {stage0_37[455]},
      {stage1_37[246]}
   );
   gpc1_1 gpc4374 (
      {stage0_37[456]},
      {stage1_37[247]}
   );
   gpc1_1 gpc4375 (
      {stage0_37[457]},
      {stage1_37[248]}
   );
   gpc1_1 gpc4376 (
      {stage0_37[458]},
      {stage1_37[249]}
   );
   gpc1_1 gpc4377 (
      {stage0_37[459]},
      {stage1_37[250]}
   );
   gpc1_1 gpc4378 (
      {stage0_37[460]},
      {stage1_37[251]}
   );
   gpc1_1 gpc4379 (
      {stage0_37[461]},
      {stage1_37[252]}
   );
   gpc1_1 gpc4380 (
      {stage0_37[462]},
      {stage1_37[253]}
   );
   gpc1_1 gpc4381 (
      {stage0_37[463]},
      {stage1_37[254]}
   );
   gpc1_1 gpc4382 (
      {stage0_37[464]},
      {stage1_37[255]}
   );
   gpc1_1 gpc4383 (
      {stage0_37[465]},
      {stage1_37[256]}
   );
   gpc1_1 gpc4384 (
      {stage0_37[466]},
      {stage1_37[257]}
   );
   gpc1_1 gpc4385 (
      {stage0_37[467]},
      {stage1_37[258]}
   );
   gpc1_1 gpc4386 (
      {stage0_37[468]},
      {stage1_37[259]}
   );
   gpc1_1 gpc4387 (
      {stage0_37[469]},
      {stage1_37[260]}
   );
   gpc1_1 gpc4388 (
      {stage0_37[470]},
      {stage1_37[261]}
   );
   gpc1_1 gpc4389 (
      {stage0_37[471]},
      {stage1_37[262]}
   );
   gpc1_1 gpc4390 (
      {stage0_37[472]},
      {stage1_37[263]}
   );
   gpc1_1 gpc4391 (
      {stage0_37[473]},
      {stage1_37[264]}
   );
   gpc1_1 gpc4392 (
      {stage0_37[474]},
      {stage1_37[265]}
   );
   gpc1_1 gpc4393 (
      {stage0_37[475]},
      {stage1_37[266]}
   );
   gpc1_1 gpc4394 (
      {stage0_37[476]},
      {stage1_37[267]}
   );
   gpc1_1 gpc4395 (
      {stage0_37[477]},
      {stage1_37[268]}
   );
   gpc1_1 gpc4396 (
      {stage0_37[478]},
      {stage1_37[269]}
   );
   gpc1_1 gpc4397 (
      {stage0_37[479]},
      {stage1_37[270]}
   );
   gpc1_1 gpc4398 (
      {stage0_37[480]},
      {stage1_37[271]}
   );
   gpc1_1 gpc4399 (
      {stage0_37[481]},
      {stage1_37[272]}
   );
   gpc1_1 gpc4400 (
      {stage0_37[482]},
      {stage1_37[273]}
   );
   gpc1_1 gpc4401 (
      {stage0_37[483]},
      {stage1_37[274]}
   );
   gpc1_1 gpc4402 (
      {stage0_37[484]},
      {stage1_37[275]}
   );
   gpc1_1 gpc4403 (
      {stage0_37[485]},
      {stage1_37[276]}
   );
   gpc1_1 gpc4404 (
      {stage0_37[486]},
      {stage1_37[277]}
   );
   gpc1_1 gpc4405 (
      {stage0_37[487]},
      {stage1_37[278]}
   );
   gpc1_1 gpc4406 (
      {stage0_37[488]},
      {stage1_37[279]}
   );
   gpc1_1 gpc4407 (
      {stage0_37[489]},
      {stage1_37[280]}
   );
   gpc1_1 gpc4408 (
      {stage0_37[490]},
      {stage1_37[281]}
   );
   gpc1_1 gpc4409 (
      {stage0_37[491]},
      {stage1_37[282]}
   );
   gpc1_1 gpc4410 (
      {stage0_37[492]},
      {stage1_37[283]}
   );
   gpc1_1 gpc4411 (
      {stage0_37[493]},
      {stage1_37[284]}
   );
   gpc1_1 gpc4412 (
      {stage0_37[494]},
      {stage1_37[285]}
   );
   gpc1_1 gpc4413 (
      {stage0_37[495]},
      {stage1_37[286]}
   );
   gpc1_1 gpc4414 (
      {stage0_37[496]},
      {stage1_37[287]}
   );
   gpc1_1 gpc4415 (
      {stage0_37[497]},
      {stage1_37[288]}
   );
   gpc1_1 gpc4416 (
      {stage0_37[498]},
      {stage1_37[289]}
   );
   gpc1_1 gpc4417 (
      {stage0_37[499]},
      {stage1_37[290]}
   );
   gpc1_1 gpc4418 (
      {stage0_37[500]},
      {stage1_37[291]}
   );
   gpc1_1 gpc4419 (
      {stage0_37[501]},
      {stage1_37[292]}
   );
   gpc1_1 gpc4420 (
      {stage0_37[502]},
      {stage1_37[293]}
   );
   gpc1_1 gpc4421 (
      {stage0_37[503]},
      {stage1_37[294]}
   );
   gpc1_1 gpc4422 (
      {stage0_37[504]},
      {stage1_37[295]}
   );
   gpc1_1 gpc4423 (
      {stage0_37[505]},
      {stage1_37[296]}
   );
   gpc1_1 gpc4424 (
      {stage0_37[506]},
      {stage1_37[297]}
   );
   gpc1_1 gpc4425 (
      {stage0_37[507]},
      {stage1_37[298]}
   );
   gpc1_1 gpc4426 (
      {stage0_37[508]},
      {stage1_37[299]}
   );
   gpc1_1 gpc4427 (
      {stage0_37[509]},
      {stage1_37[300]}
   );
   gpc1_1 gpc4428 (
      {stage0_37[510]},
      {stage1_37[301]}
   );
   gpc1_1 gpc4429 (
      {stage0_37[511]},
      {stage1_37[302]}
   );
   gpc1_1 gpc4430 (
      {stage0_38[382]},
      {stage1_38[147]}
   );
   gpc1_1 gpc4431 (
      {stage0_38[383]},
      {stage1_38[148]}
   );
   gpc1_1 gpc4432 (
      {stage0_38[384]},
      {stage1_38[149]}
   );
   gpc1_1 gpc4433 (
      {stage0_38[385]},
      {stage1_38[150]}
   );
   gpc1_1 gpc4434 (
      {stage0_38[386]},
      {stage1_38[151]}
   );
   gpc1_1 gpc4435 (
      {stage0_38[387]},
      {stage1_38[152]}
   );
   gpc1_1 gpc4436 (
      {stage0_38[388]},
      {stage1_38[153]}
   );
   gpc1_1 gpc4437 (
      {stage0_38[389]},
      {stage1_38[154]}
   );
   gpc1_1 gpc4438 (
      {stage0_38[390]},
      {stage1_38[155]}
   );
   gpc1_1 gpc4439 (
      {stage0_38[391]},
      {stage1_38[156]}
   );
   gpc1_1 gpc4440 (
      {stage0_38[392]},
      {stage1_38[157]}
   );
   gpc1_1 gpc4441 (
      {stage0_38[393]},
      {stage1_38[158]}
   );
   gpc1_1 gpc4442 (
      {stage0_38[394]},
      {stage1_38[159]}
   );
   gpc1_1 gpc4443 (
      {stage0_38[395]},
      {stage1_38[160]}
   );
   gpc1_1 gpc4444 (
      {stage0_38[396]},
      {stage1_38[161]}
   );
   gpc1_1 gpc4445 (
      {stage0_38[397]},
      {stage1_38[162]}
   );
   gpc1_1 gpc4446 (
      {stage0_38[398]},
      {stage1_38[163]}
   );
   gpc1_1 gpc4447 (
      {stage0_38[399]},
      {stage1_38[164]}
   );
   gpc1_1 gpc4448 (
      {stage0_38[400]},
      {stage1_38[165]}
   );
   gpc1_1 gpc4449 (
      {stage0_38[401]},
      {stage1_38[166]}
   );
   gpc1_1 gpc4450 (
      {stage0_38[402]},
      {stage1_38[167]}
   );
   gpc1_1 gpc4451 (
      {stage0_38[403]},
      {stage1_38[168]}
   );
   gpc1_1 gpc4452 (
      {stage0_38[404]},
      {stage1_38[169]}
   );
   gpc1_1 gpc4453 (
      {stage0_38[405]},
      {stage1_38[170]}
   );
   gpc1_1 gpc4454 (
      {stage0_38[406]},
      {stage1_38[171]}
   );
   gpc1_1 gpc4455 (
      {stage0_38[407]},
      {stage1_38[172]}
   );
   gpc1_1 gpc4456 (
      {stage0_38[408]},
      {stage1_38[173]}
   );
   gpc1_1 gpc4457 (
      {stage0_38[409]},
      {stage1_38[174]}
   );
   gpc1_1 gpc4458 (
      {stage0_38[410]},
      {stage1_38[175]}
   );
   gpc1_1 gpc4459 (
      {stage0_38[411]},
      {stage1_38[176]}
   );
   gpc1_1 gpc4460 (
      {stage0_38[412]},
      {stage1_38[177]}
   );
   gpc1_1 gpc4461 (
      {stage0_38[413]},
      {stage1_38[178]}
   );
   gpc1_1 gpc4462 (
      {stage0_38[414]},
      {stage1_38[179]}
   );
   gpc1_1 gpc4463 (
      {stage0_38[415]},
      {stage1_38[180]}
   );
   gpc1_1 gpc4464 (
      {stage0_38[416]},
      {stage1_38[181]}
   );
   gpc1_1 gpc4465 (
      {stage0_38[417]},
      {stage1_38[182]}
   );
   gpc1_1 gpc4466 (
      {stage0_38[418]},
      {stage1_38[183]}
   );
   gpc1_1 gpc4467 (
      {stage0_38[419]},
      {stage1_38[184]}
   );
   gpc1_1 gpc4468 (
      {stage0_38[420]},
      {stage1_38[185]}
   );
   gpc1_1 gpc4469 (
      {stage0_38[421]},
      {stage1_38[186]}
   );
   gpc1_1 gpc4470 (
      {stage0_38[422]},
      {stage1_38[187]}
   );
   gpc1_1 gpc4471 (
      {stage0_38[423]},
      {stage1_38[188]}
   );
   gpc1_1 gpc4472 (
      {stage0_38[424]},
      {stage1_38[189]}
   );
   gpc1_1 gpc4473 (
      {stage0_38[425]},
      {stage1_38[190]}
   );
   gpc1_1 gpc4474 (
      {stage0_38[426]},
      {stage1_38[191]}
   );
   gpc1_1 gpc4475 (
      {stage0_38[427]},
      {stage1_38[192]}
   );
   gpc1_1 gpc4476 (
      {stage0_38[428]},
      {stage1_38[193]}
   );
   gpc1_1 gpc4477 (
      {stage0_38[429]},
      {stage1_38[194]}
   );
   gpc1_1 gpc4478 (
      {stage0_38[430]},
      {stage1_38[195]}
   );
   gpc1_1 gpc4479 (
      {stage0_38[431]},
      {stage1_38[196]}
   );
   gpc1_1 gpc4480 (
      {stage0_38[432]},
      {stage1_38[197]}
   );
   gpc1_1 gpc4481 (
      {stage0_38[433]},
      {stage1_38[198]}
   );
   gpc1_1 gpc4482 (
      {stage0_38[434]},
      {stage1_38[199]}
   );
   gpc1_1 gpc4483 (
      {stage0_38[435]},
      {stage1_38[200]}
   );
   gpc1_1 gpc4484 (
      {stage0_38[436]},
      {stage1_38[201]}
   );
   gpc1_1 gpc4485 (
      {stage0_38[437]},
      {stage1_38[202]}
   );
   gpc1_1 gpc4486 (
      {stage0_38[438]},
      {stage1_38[203]}
   );
   gpc1_1 gpc4487 (
      {stage0_38[439]},
      {stage1_38[204]}
   );
   gpc1_1 gpc4488 (
      {stage0_38[440]},
      {stage1_38[205]}
   );
   gpc1_1 gpc4489 (
      {stage0_38[441]},
      {stage1_38[206]}
   );
   gpc1_1 gpc4490 (
      {stage0_38[442]},
      {stage1_38[207]}
   );
   gpc1_1 gpc4491 (
      {stage0_38[443]},
      {stage1_38[208]}
   );
   gpc1_1 gpc4492 (
      {stage0_38[444]},
      {stage1_38[209]}
   );
   gpc1_1 gpc4493 (
      {stage0_38[445]},
      {stage1_38[210]}
   );
   gpc1_1 gpc4494 (
      {stage0_38[446]},
      {stage1_38[211]}
   );
   gpc1_1 gpc4495 (
      {stage0_38[447]},
      {stage1_38[212]}
   );
   gpc1_1 gpc4496 (
      {stage0_38[448]},
      {stage1_38[213]}
   );
   gpc1_1 gpc4497 (
      {stage0_38[449]},
      {stage1_38[214]}
   );
   gpc1_1 gpc4498 (
      {stage0_38[450]},
      {stage1_38[215]}
   );
   gpc1_1 gpc4499 (
      {stage0_38[451]},
      {stage1_38[216]}
   );
   gpc1_1 gpc4500 (
      {stage0_38[452]},
      {stage1_38[217]}
   );
   gpc1_1 gpc4501 (
      {stage0_38[453]},
      {stage1_38[218]}
   );
   gpc1_1 gpc4502 (
      {stage0_38[454]},
      {stage1_38[219]}
   );
   gpc1_1 gpc4503 (
      {stage0_38[455]},
      {stage1_38[220]}
   );
   gpc1_1 gpc4504 (
      {stage0_38[456]},
      {stage1_38[221]}
   );
   gpc1_1 gpc4505 (
      {stage0_38[457]},
      {stage1_38[222]}
   );
   gpc1_1 gpc4506 (
      {stage0_38[458]},
      {stage1_38[223]}
   );
   gpc1_1 gpc4507 (
      {stage0_38[459]},
      {stage1_38[224]}
   );
   gpc1_1 gpc4508 (
      {stage0_38[460]},
      {stage1_38[225]}
   );
   gpc1_1 gpc4509 (
      {stage0_38[461]},
      {stage1_38[226]}
   );
   gpc1_1 gpc4510 (
      {stage0_38[462]},
      {stage1_38[227]}
   );
   gpc1_1 gpc4511 (
      {stage0_38[463]},
      {stage1_38[228]}
   );
   gpc1_1 gpc4512 (
      {stage0_38[464]},
      {stage1_38[229]}
   );
   gpc1_1 gpc4513 (
      {stage0_38[465]},
      {stage1_38[230]}
   );
   gpc1_1 gpc4514 (
      {stage0_38[466]},
      {stage1_38[231]}
   );
   gpc1_1 gpc4515 (
      {stage0_38[467]},
      {stage1_38[232]}
   );
   gpc1_1 gpc4516 (
      {stage0_38[468]},
      {stage1_38[233]}
   );
   gpc1_1 gpc4517 (
      {stage0_38[469]},
      {stage1_38[234]}
   );
   gpc1_1 gpc4518 (
      {stage0_38[470]},
      {stage1_38[235]}
   );
   gpc1_1 gpc4519 (
      {stage0_38[471]},
      {stage1_38[236]}
   );
   gpc1_1 gpc4520 (
      {stage0_38[472]},
      {stage1_38[237]}
   );
   gpc1_1 gpc4521 (
      {stage0_38[473]},
      {stage1_38[238]}
   );
   gpc1_1 gpc4522 (
      {stage0_38[474]},
      {stage1_38[239]}
   );
   gpc1_1 gpc4523 (
      {stage0_38[475]},
      {stage1_38[240]}
   );
   gpc1_1 gpc4524 (
      {stage0_38[476]},
      {stage1_38[241]}
   );
   gpc1_1 gpc4525 (
      {stage0_38[477]},
      {stage1_38[242]}
   );
   gpc1_1 gpc4526 (
      {stage0_38[478]},
      {stage1_38[243]}
   );
   gpc1_1 gpc4527 (
      {stage0_38[479]},
      {stage1_38[244]}
   );
   gpc1_1 gpc4528 (
      {stage0_38[480]},
      {stage1_38[245]}
   );
   gpc1_1 gpc4529 (
      {stage0_38[481]},
      {stage1_38[246]}
   );
   gpc1_1 gpc4530 (
      {stage0_38[482]},
      {stage1_38[247]}
   );
   gpc1_1 gpc4531 (
      {stage0_38[483]},
      {stage1_38[248]}
   );
   gpc1_1 gpc4532 (
      {stage0_38[484]},
      {stage1_38[249]}
   );
   gpc1_1 gpc4533 (
      {stage0_38[485]},
      {stage1_38[250]}
   );
   gpc1_1 gpc4534 (
      {stage0_38[486]},
      {stage1_38[251]}
   );
   gpc1_1 gpc4535 (
      {stage0_38[487]},
      {stage1_38[252]}
   );
   gpc1_1 gpc4536 (
      {stage0_38[488]},
      {stage1_38[253]}
   );
   gpc1_1 gpc4537 (
      {stage0_38[489]},
      {stage1_38[254]}
   );
   gpc1_1 gpc4538 (
      {stage0_38[490]},
      {stage1_38[255]}
   );
   gpc1_1 gpc4539 (
      {stage0_38[491]},
      {stage1_38[256]}
   );
   gpc1_1 gpc4540 (
      {stage0_38[492]},
      {stage1_38[257]}
   );
   gpc1_1 gpc4541 (
      {stage0_38[493]},
      {stage1_38[258]}
   );
   gpc1_1 gpc4542 (
      {stage0_38[494]},
      {stage1_38[259]}
   );
   gpc1_1 gpc4543 (
      {stage0_38[495]},
      {stage1_38[260]}
   );
   gpc1_1 gpc4544 (
      {stage0_38[496]},
      {stage1_38[261]}
   );
   gpc1_1 gpc4545 (
      {stage0_38[497]},
      {stage1_38[262]}
   );
   gpc1_1 gpc4546 (
      {stage0_38[498]},
      {stage1_38[263]}
   );
   gpc1_1 gpc4547 (
      {stage0_38[499]},
      {stage1_38[264]}
   );
   gpc1_1 gpc4548 (
      {stage0_38[500]},
      {stage1_38[265]}
   );
   gpc1_1 gpc4549 (
      {stage0_38[501]},
      {stage1_38[266]}
   );
   gpc1_1 gpc4550 (
      {stage0_38[502]},
      {stage1_38[267]}
   );
   gpc1_1 gpc4551 (
      {stage0_38[503]},
      {stage1_38[268]}
   );
   gpc1_1 gpc4552 (
      {stage0_38[504]},
      {stage1_38[269]}
   );
   gpc1_1 gpc4553 (
      {stage0_38[505]},
      {stage1_38[270]}
   );
   gpc1_1 gpc4554 (
      {stage0_38[506]},
      {stage1_38[271]}
   );
   gpc1_1 gpc4555 (
      {stage0_38[507]},
      {stage1_38[272]}
   );
   gpc1_1 gpc4556 (
      {stage0_38[508]},
      {stage1_38[273]}
   );
   gpc1_1 gpc4557 (
      {stage0_38[509]},
      {stage1_38[274]}
   );
   gpc1_1 gpc4558 (
      {stage0_38[510]},
      {stage1_38[275]}
   );
   gpc1_1 gpc4559 (
      {stage0_38[511]},
      {stage1_38[276]}
   );
   gpc1_1 gpc4560 (
      {stage0_39[491]},
      {stage1_39[176]}
   );
   gpc1_1 gpc4561 (
      {stage0_39[492]},
      {stage1_39[177]}
   );
   gpc1_1 gpc4562 (
      {stage0_39[493]},
      {stage1_39[178]}
   );
   gpc1_1 gpc4563 (
      {stage0_39[494]},
      {stage1_39[179]}
   );
   gpc1_1 gpc4564 (
      {stage0_39[495]},
      {stage1_39[180]}
   );
   gpc1_1 gpc4565 (
      {stage0_39[496]},
      {stage1_39[181]}
   );
   gpc1_1 gpc4566 (
      {stage0_39[497]},
      {stage1_39[182]}
   );
   gpc1_1 gpc4567 (
      {stage0_39[498]},
      {stage1_39[183]}
   );
   gpc1_1 gpc4568 (
      {stage0_39[499]},
      {stage1_39[184]}
   );
   gpc1_1 gpc4569 (
      {stage0_39[500]},
      {stage1_39[185]}
   );
   gpc1_1 gpc4570 (
      {stage0_39[501]},
      {stage1_39[186]}
   );
   gpc1_1 gpc4571 (
      {stage0_39[502]},
      {stage1_39[187]}
   );
   gpc1_1 gpc4572 (
      {stage0_39[503]},
      {stage1_39[188]}
   );
   gpc1_1 gpc4573 (
      {stage0_39[504]},
      {stage1_39[189]}
   );
   gpc1_1 gpc4574 (
      {stage0_39[505]},
      {stage1_39[190]}
   );
   gpc1_1 gpc4575 (
      {stage0_39[506]},
      {stage1_39[191]}
   );
   gpc1_1 gpc4576 (
      {stage0_39[507]},
      {stage1_39[192]}
   );
   gpc1_1 gpc4577 (
      {stage0_39[508]},
      {stage1_39[193]}
   );
   gpc1_1 gpc4578 (
      {stage0_39[509]},
      {stage1_39[194]}
   );
   gpc1_1 gpc4579 (
      {stage0_39[510]},
      {stage1_39[195]}
   );
   gpc1_1 gpc4580 (
      {stage0_39[511]},
      {stage1_39[196]}
   );
   gpc1_1 gpc4581 (
      {stage0_40[489]},
      {stage1_40[207]}
   );
   gpc1_1 gpc4582 (
      {stage0_40[490]},
      {stage1_40[208]}
   );
   gpc1_1 gpc4583 (
      {stage0_40[491]},
      {stage1_40[209]}
   );
   gpc1_1 gpc4584 (
      {stage0_40[492]},
      {stage1_40[210]}
   );
   gpc1_1 gpc4585 (
      {stage0_40[493]},
      {stage1_40[211]}
   );
   gpc1_1 gpc4586 (
      {stage0_40[494]},
      {stage1_40[212]}
   );
   gpc1_1 gpc4587 (
      {stage0_40[495]},
      {stage1_40[213]}
   );
   gpc1_1 gpc4588 (
      {stage0_40[496]},
      {stage1_40[214]}
   );
   gpc1_1 gpc4589 (
      {stage0_40[497]},
      {stage1_40[215]}
   );
   gpc1_1 gpc4590 (
      {stage0_40[498]},
      {stage1_40[216]}
   );
   gpc1_1 gpc4591 (
      {stage0_40[499]},
      {stage1_40[217]}
   );
   gpc1_1 gpc4592 (
      {stage0_40[500]},
      {stage1_40[218]}
   );
   gpc1_1 gpc4593 (
      {stage0_40[501]},
      {stage1_40[219]}
   );
   gpc1_1 gpc4594 (
      {stage0_40[502]},
      {stage1_40[220]}
   );
   gpc1_1 gpc4595 (
      {stage0_40[503]},
      {stage1_40[221]}
   );
   gpc1_1 gpc4596 (
      {stage0_40[504]},
      {stage1_40[222]}
   );
   gpc1_1 gpc4597 (
      {stage0_40[505]},
      {stage1_40[223]}
   );
   gpc1_1 gpc4598 (
      {stage0_40[506]},
      {stage1_40[224]}
   );
   gpc1_1 gpc4599 (
      {stage0_40[507]},
      {stage1_40[225]}
   );
   gpc1_1 gpc4600 (
      {stage0_40[508]},
      {stage1_40[226]}
   );
   gpc1_1 gpc4601 (
      {stage0_40[509]},
      {stage1_40[227]}
   );
   gpc1_1 gpc4602 (
      {stage0_40[510]},
      {stage1_40[228]}
   );
   gpc1_1 gpc4603 (
      {stage0_40[511]},
      {stage1_40[229]}
   );
   gpc1_1 gpc4604 (
      {stage0_41[420]},
      {stage1_41[185]}
   );
   gpc1_1 gpc4605 (
      {stage0_41[421]},
      {stage1_41[186]}
   );
   gpc1_1 gpc4606 (
      {stage0_41[422]},
      {stage1_41[187]}
   );
   gpc1_1 gpc4607 (
      {stage0_41[423]},
      {stage1_41[188]}
   );
   gpc1_1 gpc4608 (
      {stage0_41[424]},
      {stage1_41[189]}
   );
   gpc1_1 gpc4609 (
      {stage0_41[425]},
      {stage1_41[190]}
   );
   gpc1_1 gpc4610 (
      {stage0_41[426]},
      {stage1_41[191]}
   );
   gpc1_1 gpc4611 (
      {stage0_41[427]},
      {stage1_41[192]}
   );
   gpc1_1 gpc4612 (
      {stage0_41[428]},
      {stage1_41[193]}
   );
   gpc1_1 gpc4613 (
      {stage0_41[429]},
      {stage1_41[194]}
   );
   gpc1_1 gpc4614 (
      {stage0_41[430]},
      {stage1_41[195]}
   );
   gpc1_1 gpc4615 (
      {stage0_41[431]},
      {stage1_41[196]}
   );
   gpc1_1 gpc4616 (
      {stage0_41[432]},
      {stage1_41[197]}
   );
   gpc1_1 gpc4617 (
      {stage0_41[433]},
      {stage1_41[198]}
   );
   gpc1_1 gpc4618 (
      {stage0_41[434]},
      {stage1_41[199]}
   );
   gpc1_1 gpc4619 (
      {stage0_41[435]},
      {stage1_41[200]}
   );
   gpc1_1 gpc4620 (
      {stage0_41[436]},
      {stage1_41[201]}
   );
   gpc1_1 gpc4621 (
      {stage0_41[437]},
      {stage1_41[202]}
   );
   gpc1_1 gpc4622 (
      {stage0_41[438]},
      {stage1_41[203]}
   );
   gpc1_1 gpc4623 (
      {stage0_41[439]},
      {stage1_41[204]}
   );
   gpc1_1 gpc4624 (
      {stage0_41[440]},
      {stage1_41[205]}
   );
   gpc1_1 gpc4625 (
      {stage0_41[441]},
      {stage1_41[206]}
   );
   gpc1_1 gpc4626 (
      {stage0_41[442]},
      {stage1_41[207]}
   );
   gpc1_1 gpc4627 (
      {stage0_41[443]},
      {stage1_41[208]}
   );
   gpc1_1 gpc4628 (
      {stage0_41[444]},
      {stage1_41[209]}
   );
   gpc1_1 gpc4629 (
      {stage0_41[445]},
      {stage1_41[210]}
   );
   gpc1_1 gpc4630 (
      {stage0_41[446]},
      {stage1_41[211]}
   );
   gpc1_1 gpc4631 (
      {stage0_41[447]},
      {stage1_41[212]}
   );
   gpc1_1 gpc4632 (
      {stage0_41[448]},
      {stage1_41[213]}
   );
   gpc1_1 gpc4633 (
      {stage0_41[449]},
      {stage1_41[214]}
   );
   gpc1_1 gpc4634 (
      {stage0_41[450]},
      {stage1_41[215]}
   );
   gpc1_1 gpc4635 (
      {stage0_41[451]},
      {stage1_41[216]}
   );
   gpc1_1 gpc4636 (
      {stage0_41[452]},
      {stage1_41[217]}
   );
   gpc1_1 gpc4637 (
      {stage0_41[453]},
      {stage1_41[218]}
   );
   gpc1_1 gpc4638 (
      {stage0_41[454]},
      {stage1_41[219]}
   );
   gpc1_1 gpc4639 (
      {stage0_41[455]},
      {stage1_41[220]}
   );
   gpc1_1 gpc4640 (
      {stage0_41[456]},
      {stage1_41[221]}
   );
   gpc1_1 gpc4641 (
      {stage0_41[457]},
      {stage1_41[222]}
   );
   gpc1_1 gpc4642 (
      {stage0_41[458]},
      {stage1_41[223]}
   );
   gpc1_1 gpc4643 (
      {stage0_41[459]},
      {stage1_41[224]}
   );
   gpc1_1 gpc4644 (
      {stage0_41[460]},
      {stage1_41[225]}
   );
   gpc1_1 gpc4645 (
      {stage0_41[461]},
      {stage1_41[226]}
   );
   gpc1_1 gpc4646 (
      {stage0_41[462]},
      {stage1_41[227]}
   );
   gpc1_1 gpc4647 (
      {stage0_41[463]},
      {stage1_41[228]}
   );
   gpc1_1 gpc4648 (
      {stage0_41[464]},
      {stage1_41[229]}
   );
   gpc1_1 gpc4649 (
      {stage0_41[465]},
      {stage1_41[230]}
   );
   gpc1_1 gpc4650 (
      {stage0_41[466]},
      {stage1_41[231]}
   );
   gpc1_1 gpc4651 (
      {stage0_41[467]},
      {stage1_41[232]}
   );
   gpc1_1 gpc4652 (
      {stage0_41[468]},
      {stage1_41[233]}
   );
   gpc1_1 gpc4653 (
      {stage0_41[469]},
      {stage1_41[234]}
   );
   gpc1_1 gpc4654 (
      {stage0_41[470]},
      {stage1_41[235]}
   );
   gpc1_1 gpc4655 (
      {stage0_41[471]},
      {stage1_41[236]}
   );
   gpc1_1 gpc4656 (
      {stage0_41[472]},
      {stage1_41[237]}
   );
   gpc1_1 gpc4657 (
      {stage0_41[473]},
      {stage1_41[238]}
   );
   gpc1_1 gpc4658 (
      {stage0_41[474]},
      {stage1_41[239]}
   );
   gpc1_1 gpc4659 (
      {stage0_41[475]},
      {stage1_41[240]}
   );
   gpc1_1 gpc4660 (
      {stage0_41[476]},
      {stage1_41[241]}
   );
   gpc1_1 gpc4661 (
      {stage0_41[477]},
      {stage1_41[242]}
   );
   gpc1_1 gpc4662 (
      {stage0_41[478]},
      {stage1_41[243]}
   );
   gpc1_1 gpc4663 (
      {stage0_41[479]},
      {stage1_41[244]}
   );
   gpc1_1 gpc4664 (
      {stage0_41[480]},
      {stage1_41[245]}
   );
   gpc1_1 gpc4665 (
      {stage0_41[481]},
      {stage1_41[246]}
   );
   gpc1_1 gpc4666 (
      {stage0_41[482]},
      {stage1_41[247]}
   );
   gpc1_1 gpc4667 (
      {stage0_41[483]},
      {stage1_41[248]}
   );
   gpc1_1 gpc4668 (
      {stage0_41[484]},
      {stage1_41[249]}
   );
   gpc1_1 gpc4669 (
      {stage0_41[485]},
      {stage1_41[250]}
   );
   gpc1_1 gpc4670 (
      {stage0_41[486]},
      {stage1_41[251]}
   );
   gpc1_1 gpc4671 (
      {stage0_41[487]},
      {stage1_41[252]}
   );
   gpc1_1 gpc4672 (
      {stage0_41[488]},
      {stage1_41[253]}
   );
   gpc1_1 gpc4673 (
      {stage0_41[489]},
      {stage1_41[254]}
   );
   gpc1_1 gpc4674 (
      {stage0_41[490]},
      {stage1_41[255]}
   );
   gpc1_1 gpc4675 (
      {stage0_41[491]},
      {stage1_41[256]}
   );
   gpc1_1 gpc4676 (
      {stage0_41[492]},
      {stage1_41[257]}
   );
   gpc1_1 gpc4677 (
      {stage0_41[493]},
      {stage1_41[258]}
   );
   gpc1_1 gpc4678 (
      {stage0_41[494]},
      {stage1_41[259]}
   );
   gpc1_1 gpc4679 (
      {stage0_41[495]},
      {stage1_41[260]}
   );
   gpc1_1 gpc4680 (
      {stage0_41[496]},
      {stage1_41[261]}
   );
   gpc1_1 gpc4681 (
      {stage0_41[497]},
      {stage1_41[262]}
   );
   gpc1_1 gpc4682 (
      {stage0_41[498]},
      {stage1_41[263]}
   );
   gpc1_1 gpc4683 (
      {stage0_41[499]},
      {stage1_41[264]}
   );
   gpc1_1 gpc4684 (
      {stage0_41[500]},
      {stage1_41[265]}
   );
   gpc1_1 gpc4685 (
      {stage0_41[501]},
      {stage1_41[266]}
   );
   gpc1_1 gpc4686 (
      {stage0_41[502]},
      {stage1_41[267]}
   );
   gpc1_1 gpc4687 (
      {stage0_41[503]},
      {stage1_41[268]}
   );
   gpc1_1 gpc4688 (
      {stage0_41[504]},
      {stage1_41[269]}
   );
   gpc1_1 gpc4689 (
      {stage0_41[505]},
      {stage1_41[270]}
   );
   gpc1_1 gpc4690 (
      {stage0_41[506]},
      {stage1_41[271]}
   );
   gpc1_1 gpc4691 (
      {stage0_41[507]},
      {stage1_41[272]}
   );
   gpc1_1 gpc4692 (
      {stage0_41[508]},
      {stage1_41[273]}
   );
   gpc1_1 gpc4693 (
      {stage0_41[509]},
      {stage1_41[274]}
   );
   gpc1_1 gpc4694 (
      {stage0_41[510]},
      {stage1_41[275]}
   );
   gpc1_1 gpc4695 (
      {stage0_41[511]},
      {stage1_41[276]}
   );
   gpc1_1 gpc4696 (
      {stage0_42[451]},
      {stage1_42[168]}
   );
   gpc1_1 gpc4697 (
      {stage0_42[452]},
      {stage1_42[169]}
   );
   gpc1_1 gpc4698 (
      {stage0_42[453]},
      {stage1_42[170]}
   );
   gpc1_1 gpc4699 (
      {stage0_42[454]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4700 (
      {stage0_42[455]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4701 (
      {stage0_42[456]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4702 (
      {stage0_42[457]},
      {stage1_42[174]}
   );
   gpc1_1 gpc4703 (
      {stage0_42[458]},
      {stage1_42[175]}
   );
   gpc1_1 gpc4704 (
      {stage0_42[459]},
      {stage1_42[176]}
   );
   gpc1_1 gpc4705 (
      {stage0_42[460]},
      {stage1_42[177]}
   );
   gpc1_1 gpc4706 (
      {stage0_42[461]},
      {stage1_42[178]}
   );
   gpc1_1 gpc4707 (
      {stage0_42[462]},
      {stage1_42[179]}
   );
   gpc1_1 gpc4708 (
      {stage0_42[463]},
      {stage1_42[180]}
   );
   gpc1_1 gpc4709 (
      {stage0_42[464]},
      {stage1_42[181]}
   );
   gpc1_1 gpc4710 (
      {stage0_42[465]},
      {stage1_42[182]}
   );
   gpc1_1 gpc4711 (
      {stage0_42[466]},
      {stage1_42[183]}
   );
   gpc1_1 gpc4712 (
      {stage0_42[467]},
      {stage1_42[184]}
   );
   gpc1_1 gpc4713 (
      {stage0_42[468]},
      {stage1_42[185]}
   );
   gpc1_1 gpc4714 (
      {stage0_42[469]},
      {stage1_42[186]}
   );
   gpc1_1 gpc4715 (
      {stage0_42[470]},
      {stage1_42[187]}
   );
   gpc1_1 gpc4716 (
      {stage0_42[471]},
      {stage1_42[188]}
   );
   gpc1_1 gpc4717 (
      {stage0_42[472]},
      {stage1_42[189]}
   );
   gpc1_1 gpc4718 (
      {stage0_42[473]},
      {stage1_42[190]}
   );
   gpc1_1 gpc4719 (
      {stage0_42[474]},
      {stage1_42[191]}
   );
   gpc1_1 gpc4720 (
      {stage0_42[475]},
      {stage1_42[192]}
   );
   gpc1_1 gpc4721 (
      {stage0_42[476]},
      {stage1_42[193]}
   );
   gpc1_1 gpc4722 (
      {stage0_42[477]},
      {stage1_42[194]}
   );
   gpc1_1 gpc4723 (
      {stage0_42[478]},
      {stage1_42[195]}
   );
   gpc1_1 gpc4724 (
      {stage0_42[479]},
      {stage1_42[196]}
   );
   gpc1_1 gpc4725 (
      {stage0_42[480]},
      {stage1_42[197]}
   );
   gpc1_1 gpc4726 (
      {stage0_42[481]},
      {stage1_42[198]}
   );
   gpc1_1 gpc4727 (
      {stage0_42[482]},
      {stage1_42[199]}
   );
   gpc1_1 gpc4728 (
      {stage0_42[483]},
      {stage1_42[200]}
   );
   gpc1_1 gpc4729 (
      {stage0_42[484]},
      {stage1_42[201]}
   );
   gpc1_1 gpc4730 (
      {stage0_42[485]},
      {stage1_42[202]}
   );
   gpc1_1 gpc4731 (
      {stage0_42[486]},
      {stage1_42[203]}
   );
   gpc1_1 gpc4732 (
      {stage0_42[487]},
      {stage1_42[204]}
   );
   gpc1_1 gpc4733 (
      {stage0_42[488]},
      {stage1_42[205]}
   );
   gpc1_1 gpc4734 (
      {stage0_42[489]},
      {stage1_42[206]}
   );
   gpc1_1 gpc4735 (
      {stage0_42[490]},
      {stage1_42[207]}
   );
   gpc1_1 gpc4736 (
      {stage0_42[491]},
      {stage1_42[208]}
   );
   gpc1_1 gpc4737 (
      {stage0_42[492]},
      {stage1_42[209]}
   );
   gpc1_1 gpc4738 (
      {stage0_42[493]},
      {stage1_42[210]}
   );
   gpc1_1 gpc4739 (
      {stage0_42[494]},
      {stage1_42[211]}
   );
   gpc1_1 gpc4740 (
      {stage0_42[495]},
      {stage1_42[212]}
   );
   gpc1_1 gpc4741 (
      {stage0_42[496]},
      {stage1_42[213]}
   );
   gpc1_1 gpc4742 (
      {stage0_42[497]},
      {stage1_42[214]}
   );
   gpc1_1 gpc4743 (
      {stage0_42[498]},
      {stage1_42[215]}
   );
   gpc1_1 gpc4744 (
      {stage0_42[499]},
      {stage1_42[216]}
   );
   gpc1_1 gpc4745 (
      {stage0_42[500]},
      {stage1_42[217]}
   );
   gpc1_1 gpc4746 (
      {stage0_42[501]},
      {stage1_42[218]}
   );
   gpc1_1 gpc4747 (
      {stage0_42[502]},
      {stage1_42[219]}
   );
   gpc1_1 gpc4748 (
      {stage0_42[503]},
      {stage1_42[220]}
   );
   gpc1_1 gpc4749 (
      {stage0_42[504]},
      {stage1_42[221]}
   );
   gpc1_1 gpc4750 (
      {stage0_42[505]},
      {stage1_42[222]}
   );
   gpc1_1 gpc4751 (
      {stage0_42[506]},
      {stage1_42[223]}
   );
   gpc1_1 gpc4752 (
      {stage0_42[507]},
      {stage1_42[224]}
   );
   gpc1_1 gpc4753 (
      {stage0_42[508]},
      {stage1_42[225]}
   );
   gpc1_1 gpc4754 (
      {stage0_42[509]},
      {stage1_42[226]}
   );
   gpc1_1 gpc4755 (
      {stage0_42[510]},
      {stage1_42[227]}
   );
   gpc1_1 gpc4756 (
      {stage0_42[511]},
      {stage1_42[228]}
   );
   gpc1_1 gpc4757 (
      {stage0_43[475]},
      {stage1_43[207]}
   );
   gpc1_1 gpc4758 (
      {stage0_43[476]},
      {stage1_43[208]}
   );
   gpc1_1 gpc4759 (
      {stage0_43[477]},
      {stage1_43[209]}
   );
   gpc1_1 gpc4760 (
      {stage0_43[478]},
      {stage1_43[210]}
   );
   gpc1_1 gpc4761 (
      {stage0_43[479]},
      {stage1_43[211]}
   );
   gpc1_1 gpc4762 (
      {stage0_43[480]},
      {stage1_43[212]}
   );
   gpc1_1 gpc4763 (
      {stage0_43[481]},
      {stage1_43[213]}
   );
   gpc1_1 gpc4764 (
      {stage0_43[482]},
      {stage1_43[214]}
   );
   gpc1_1 gpc4765 (
      {stage0_43[483]},
      {stage1_43[215]}
   );
   gpc1_1 gpc4766 (
      {stage0_43[484]},
      {stage1_43[216]}
   );
   gpc1_1 gpc4767 (
      {stage0_43[485]},
      {stage1_43[217]}
   );
   gpc1_1 gpc4768 (
      {stage0_43[486]},
      {stage1_43[218]}
   );
   gpc1_1 gpc4769 (
      {stage0_43[487]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4770 (
      {stage0_43[488]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4771 (
      {stage0_43[489]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4772 (
      {stage0_43[490]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4773 (
      {stage0_43[491]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4774 (
      {stage0_43[492]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4775 (
      {stage0_43[493]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4776 (
      {stage0_43[494]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4777 (
      {stage0_43[495]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4778 (
      {stage0_43[496]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4779 (
      {stage0_43[497]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4780 (
      {stage0_43[498]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4781 (
      {stage0_43[499]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4782 (
      {stage0_43[500]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4783 (
      {stage0_43[501]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4784 (
      {stage0_43[502]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4785 (
      {stage0_43[503]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4786 (
      {stage0_43[504]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4787 (
      {stage0_43[505]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4788 (
      {stage0_43[506]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4789 (
      {stage0_43[507]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4790 (
      {stage0_43[508]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4791 (
      {stage0_43[509]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4792 (
      {stage0_43[510]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4793 (
      {stage0_43[511]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4794 (
      {stage0_44[448]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4795 (
      {stage0_44[449]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4796 (
      {stage0_44[450]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4797 (
      {stage0_44[451]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4798 (
      {stage0_44[452]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4799 (
      {stage0_44[453]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4800 (
      {stage0_44[454]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4801 (
      {stage0_44[455]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4802 (
      {stage0_44[456]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4803 (
      {stage0_44[457]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4804 (
      {stage0_44[458]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4805 (
      {stage0_44[459]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4806 (
      {stage0_44[460]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4807 (
      {stage0_44[461]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4808 (
      {stage0_44[462]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4809 (
      {stage0_44[463]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4810 (
      {stage0_44[464]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4811 (
      {stage0_44[465]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4812 (
      {stage0_44[466]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4813 (
      {stage0_44[467]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4814 (
      {stage0_44[468]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4815 (
      {stage0_44[469]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4816 (
      {stage0_44[470]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4817 (
      {stage0_44[471]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4818 (
      {stage0_44[472]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4819 (
      {stage0_44[473]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4820 (
      {stage0_44[474]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4821 (
      {stage0_44[475]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4822 (
      {stage0_44[476]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4823 (
      {stage0_44[477]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4824 (
      {stage0_44[478]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4825 (
      {stage0_44[479]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4826 (
      {stage0_44[480]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4827 (
      {stage0_44[481]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4828 (
      {stage0_44[482]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4829 (
      {stage0_44[483]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4830 (
      {stage0_44[484]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4831 (
      {stage0_44[485]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4832 (
      {stage0_44[486]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4833 (
      {stage0_44[487]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4834 (
      {stage0_44[488]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4835 (
      {stage0_44[489]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4836 (
      {stage0_44[490]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4837 (
      {stage0_44[491]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4838 (
      {stage0_44[492]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4839 (
      {stage0_44[493]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4840 (
      {stage0_44[494]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4841 (
      {stage0_44[495]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4842 (
      {stage0_44[496]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4843 (
      {stage0_44[497]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4844 (
      {stage0_44[498]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4845 (
      {stage0_44[499]},
      {stage1_44[256]}
   );
   gpc1_1 gpc4846 (
      {stage0_44[500]},
      {stage1_44[257]}
   );
   gpc1_1 gpc4847 (
      {stage0_44[501]},
      {stage1_44[258]}
   );
   gpc1_1 gpc4848 (
      {stage0_44[502]},
      {stage1_44[259]}
   );
   gpc1_1 gpc4849 (
      {stage0_44[503]},
      {stage1_44[260]}
   );
   gpc1_1 gpc4850 (
      {stage0_44[504]},
      {stage1_44[261]}
   );
   gpc1_1 gpc4851 (
      {stage0_44[505]},
      {stage1_44[262]}
   );
   gpc1_1 gpc4852 (
      {stage0_44[506]},
      {stage1_44[263]}
   );
   gpc1_1 gpc4853 (
      {stage0_44[507]},
      {stage1_44[264]}
   );
   gpc1_1 gpc4854 (
      {stage0_44[508]},
      {stage1_44[265]}
   );
   gpc1_1 gpc4855 (
      {stage0_44[509]},
      {stage1_44[266]}
   );
   gpc1_1 gpc4856 (
      {stage0_44[510]},
      {stage1_44[267]}
   );
   gpc1_1 gpc4857 (
      {stage0_44[511]},
      {stage1_44[268]}
   );
   gpc1_1 gpc4858 (
      {stage0_45[498]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4859 (
      {stage0_45[499]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4860 (
      {stage0_45[500]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4861 (
      {stage0_45[501]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4862 (
      {stage0_45[502]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4863 (
      {stage0_45[503]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4864 (
      {stage0_45[504]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4865 (
      {stage0_45[505]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4866 (
      {stage0_45[506]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4867 (
      {stage0_45[507]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4868 (
      {stage0_45[508]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4869 (
      {stage0_45[509]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4870 (
      {stage0_45[510]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4871 (
      {stage0_45[511]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4872 (
      {stage0_46[388]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4873 (
      {stage0_46[389]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4874 (
      {stage0_46[390]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4875 (
      {stage0_46[391]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4876 (
      {stage0_46[392]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4877 (
      {stage0_46[393]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4878 (
      {stage0_46[394]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4879 (
      {stage0_46[395]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4880 (
      {stage0_46[396]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4881 (
      {stage0_46[397]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4882 (
      {stage0_46[398]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4883 (
      {stage0_46[399]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4884 (
      {stage0_46[400]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4885 (
      {stage0_46[401]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4886 (
      {stage0_46[402]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4887 (
      {stage0_46[403]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4888 (
      {stage0_46[404]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4889 (
      {stage0_46[405]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4890 (
      {stage0_46[406]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4891 (
      {stage0_46[407]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4892 (
      {stage0_46[408]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4893 (
      {stage0_46[409]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4894 (
      {stage0_46[410]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4895 (
      {stage0_46[411]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4896 (
      {stage0_46[412]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4897 (
      {stage0_46[413]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4898 (
      {stage0_46[414]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4899 (
      {stage0_46[415]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4900 (
      {stage0_46[416]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4901 (
      {stage0_46[417]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4902 (
      {stage0_46[418]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4903 (
      {stage0_46[419]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4904 (
      {stage0_46[420]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4905 (
      {stage0_46[421]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4906 (
      {stage0_46[422]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4907 (
      {stage0_46[423]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4908 (
      {stage0_46[424]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4909 (
      {stage0_46[425]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4910 (
      {stage0_46[426]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4911 (
      {stage0_46[427]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4912 (
      {stage0_46[428]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4913 (
      {stage0_46[429]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4914 (
      {stage0_46[430]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4915 (
      {stage0_46[431]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4916 (
      {stage0_46[432]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4917 (
      {stage0_46[433]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4918 (
      {stage0_46[434]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4919 (
      {stage0_46[435]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4920 (
      {stage0_46[436]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4921 (
      {stage0_46[437]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4922 (
      {stage0_46[438]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4923 (
      {stage0_46[439]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4924 (
      {stage0_46[440]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4925 (
      {stage0_46[441]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4926 (
      {stage0_46[442]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4927 (
      {stage0_46[443]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4928 (
      {stage0_46[444]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4929 (
      {stage0_46[445]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4930 (
      {stage0_46[446]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4931 (
      {stage0_46[447]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4932 (
      {stage0_46[448]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4933 (
      {stage0_46[449]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4934 (
      {stage0_46[450]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4935 (
      {stage0_46[451]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4936 (
      {stage0_46[452]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4937 (
      {stage0_46[453]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4938 (
      {stage0_46[454]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4939 (
      {stage0_46[455]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4940 (
      {stage0_46[456]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4941 (
      {stage0_46[457]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4942 (
      {stage0_46[458]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4943 (
      {stage0_46[459]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4944 (
      {stage0_46[460]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4945 (
      {stage0_46[461]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4946 (
      {stage0_46[462]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4947 (
      {stage0_46[463]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4948 (
      {stage0_46[464]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4949 (
      {stage0_46[465]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4950 (
      {stage0_46[466]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4951 (
      {stage0_46[467]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4952 (
      {stage0_46[468]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4953 (
      {stage0_46[469]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4954 (
      {stage0_46[470]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4955 (
      {stage0_46[471]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4956 (
      {stage0_46[472]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4957 (
      {stage0_46[473]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4958 (
      {stage0_46[474]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4959 (
      {stage0_46[475]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4960 (
      {stage0_46[476]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4961 (
      {stage0_46[477]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4962 (
      {stage0_46[478]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4963 (
      {stage0_46[479]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4964 (
      {stage0_46[480]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4965 (
      {stage0_46[481]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4966 (
      {stage0_46[482]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4967 (
      {stage0_46[483]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4968 (
      {stage0_46[484]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4969 (
      {stage0_46[485]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4970 (
      {stage0_46[486]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4971 (
      {stage0_46[487]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4972 (
      {stage0_46[488]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4973 (
      {stage0_46[489]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4974 (
      {stage0_46[490]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4975 (
      {stage0_46[491]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4976 (
      {stage0_46[492]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4977 (
      {stage0_46[493]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4978 (
      {stage0_46[494]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4979 (
      {stage0_46[495]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4980 (
      {stage0_46[496]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4981 (
      {stage0_46[497]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4982 (
      {stage0_46[498]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4983 (
      {stage0_46[499]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4984 (
      {stage0_46[500]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4985 (
      {stage0_46[501]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4986 (
      {stage0_46[502]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4987 (
      {stage0_46[503]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4988 (
      {stage0_46[504]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4989 (
      {stage0_46[505]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4990 (
      {stage0_46[506]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4991 (
      {stage0_46[507]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4992 (
      {stage0_46[508]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4993 (
      {stage0_46[509]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4994 (
      {stage0_46[510]},
      {stage1_46[298]}
   );
   gpc1_1 gpc4995 (
      {stage0_46[511]},
      {stage1_46[299]}
   );
   gpc1_1 gpc4996 (
      {stage0_47[437]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4997 (
      {stage0_47[438]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4998 (
      {stage0_47[439]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4999 (
      {stage0_47[440]},
      {stage1_47[206]}
   );
   gpc1_1 gpc5000 (
      {stage0_47[441]},
      {stage1_47[207]}
   );
   gpc1_1 gpc5001 (
      {stage0_47[442]},
      {stage1_47[208]}
   );
   gpc1_1 gpc5002 (
      {stage0_47[443]},
      {stage1_47[209]}
   );
   gpc1_1 gpc5003 (
      {stage0_47[444]},
      {stage1_47[210]}
   );
   gpc1_1 gpc5004 (
      {stage0_47[445]},
      {stage1_47[211]}
   );
   gpc1_1 gpc5005 (
      {stage0_47[446]},
      {stage1_47[212]}
   );
   gpc1_1 gpc5006 (
      {stage0_47[447]},
      {stage1_47[213]}
   );
   gpc1_1 gpc5007 (
      {stage0_47[448]},
      {stage1_47[214]}
   );
   gpc1_1 gpc5008 (
      {stage0_47[449]},
      {stage1_47[215]}
   );
   gpc1_1 gpc5009 (
      {stage0_47[450]},
      {stage1_47[216]}
   );
   gpc1_1 gpc5010 (
      {stage0_47[451]},
      {stage1_47[217]}
   );
   gpc1_1 gpc5011 (
      {stage0_47[452]},
      {stage1_47[218]}
   );
   gpc1_1 gpc5012 (
      {stage0_47[453]},
      {stage1_47[219]}
   );
   gpc1_1 gpc5013 (
      {stage0_47[454]},
      {stage1_47[220]}
   );
   gpc1_1 gpc5014 (
      {stage0_47[455]},
      {stage1_47[221]}
   );
   gpc1_1 gpc5015 (
      {stage0_47[456]},
      {stage1_47[222]}
   );
   gpc1_1 gpc5016 (
      {stage0_47[457]},
      {stage1_47[223]}
   );
   gpc1_1 gpc5017 (
      {stage0_47[458]},
      {stage1_47[224]}
   );
   gpc1_1 gpc5018 (
      {stage0_47[459]},
      {stage1_47[225]}
   );
   gpc1_1 gpc5019 (
      {stage0_47[460]},
      {stage1_47[226]}
   );
   gpc1_1 gpc5020 (
      {stage0_47[461]},
      {stage1_47[227]}
   );
   gpc1_1 gpc5021 (
      {stage0_47[462]},
      {stage1_47[228]}
   );
   gpc1_1 gpc5022 (
      {stage0_47[463]},
      {stage1_47[229]}
   );
   gpc1_1 gpc5023 (
      {stage0_47[464]},
      {stage1_47[230]}
   );
   gpc1_1 gpc5024 (
      {stage0_47[465]},
      {stage1_47[231]}
   );
   gpc1_1 gpc5025 (
      {stage0_47[466]},
      {stage1_47[232]}
   );
   gpc1_1 gpc5026 (
      {stage0_47[467]},
      {stage1_47[233]}
   );
   gpc1_1 gpc5027 (
      {stage0_47[468]},
      {stage1_47[234]}
   );
   gpc1_1 gpc5028 (
      {stage0_47[469]},
      {stage1_47[235]}
   );
   gpc1_1 gpc5029 (
      {stage0_47[470]},
      {stage1_47[236]}
   );
   gpc1_1 gpc5030 (
      {stage0_47[471]},
      {stage1_47[237]}
   );
   gpc1_1 gpc5031 (
      {stage0_47[472]},
      {stage1_47[238]}
   );
   gpc1_1 gpc5032 (
      {stage0_47[473]},
      {stage1_47[239]}
   );
   gpc1_1 gpc5033 (
      {stage0_47[474]},
      {stage1_47[240]}
   );
   gpc1_1 gpc5034 (
      {stage0_47[475]},
      {stage1_47[241]}
   );
   gpc1_1 gpc5035 (
      {stage0_47[476]},
      {stage1_47[242]}
   );
   gpc1_1 gpc5036 (
      {stage0_47[477]},
      {stage1_47[243]}
   );
   gpc1_1 gpc5037 (
      {stage0_47[478]},
      {stage1_47[244]}
   );
   gpc1_1 gpc5038 (
      {stage0_47[479]},
      {stage1_47[245]}
   );
   gpc1_1 gpc5039 (
      {stage0_47[480]},
      {stage1_47[246]}
   );
   gpc1_1 gpc5040 (
      {stage0_47[481]},
      {stage1_47[247]}
   );
   gpc1_1 gpc5041 (
      {stage0_47[482]},
      {stage1_47[248]}
   );
   gpc1_1 gpc5042 (
      {stage0_47[483]},
      {stage1_47[249]}
   );
   gpc1_1 gpc5043 (
      {stage0_47[484]},
      {stage1_47[250]}
   );
   gpc1_1 gpc5044 (
      {stage0_47[485]},
      {stage1_47[251]}
   );
   gpc1_1 gpc5045 (
      {stage0_47[486]},
      {stage1_47[252]}
   );
   gpc1_1 gpc5046 (
      {stage0_47[487]},
      {stage1_47[253]}
   );
   gpc1_1 gpc5047 (
      {stage0_47[488]},
      {stage1_47[254]}
   );
   gpc1_1 gpc5048 (
      {stage0_47[489]},
      {stage1_47[255]}
   );
   gpc1_1 gpc5049 (
      {stage0_47[490]},
      {stage1_47[256]}
   );
   gpc1_1 gpc5050 (
      {stage0_47[491]},
      {stage1_47[257]}
   );
   gpc1_1 gpc5051 (
      {stage0_47[492]},
      {stage1_47[258]}
   );
   gpc1_1 gpc5052 (
      {stage0_47[493]},
      {stage1_47[259]}
   );
   gpc1_1 gpc5053 (
      {stage0_47[494]},
      {stage1_47[260]}
   );
   gpc1_1 gpc5054 (
      {stage0_47[495]},
      {stage1_47[261]}
   );
   gpc1_1 gpc5055 (
      {stage0_47[496]},
      {stage1_47[262]}
   );
   gpc1_1 gpc5056 (
      {stage0_47[497]},
      {stage1_47[263]}
   );
   gpc1_1 gpc5057 (
      {stage0_47[498]},
      {stage1_47[264]}
   );
   gpc1_1 gpc5058 (
      {stage0_47[499]},
      {stage1_47[265]}
   );
   gpc1_1 gpc5059 (
      {stage0_47[500]},
      {stage1_47[266]}
   );
   gpc1_1 gpc5060 (
      {stage0_47[501]},
      {stage1_47[267]}
   );
   gpc1_1 gpc5061 (
      {stage0_47[502]},
      {stage1_47[268]}
   );
   gpc1_1 gpc5062 (
      {stage0_47[503]},
      {stage1_47[269]}
   );
   gpc1_1 gpc5063 (
      {stage0_47[504]},
      {stage1_47[270]}
   );
   gpc1_1 gpc5064 (
      {stage0_47[505]},
      {stage1_47[271]}
   );
   gpc1_1 gpc5065 (
      {stage0_47[506]},
      {stage1_47[272]}
   );
   gpc1_1 gpc5066 (
      {stage0_47[507]},
      {stage1_47[273]}
   );
   gpc1_1 gpc5067 (
      {stage0_47[508]},
      {stage1_47[274]}
   );
   gpc1_1 gpc5068 (
      {stage0_47[509]},
      {stage1_47[275]}
   );
   gpc1_1 gpc5069 (
      {stage0_47[510]},
      {stage1_47[276]}
   );
   gpc1_1 gpc5070 (
      {stage0_47[511]},
      {stage1_47[277]}
   );
   gpc1_1 gpc5071 (
      {stage0_48[495]},
      {stage1_48[194]}
   );
   gpc1_1 gpc5072 (
      {stage0_48[496]},
      {stage1_48[195]}
   );
   gpc1_1 gpc5073 (
      {stage0_48[497]},
      {stage1_48[196]}
   );
   gpc1_1 gpc5074 (
      {stage0_48[498]},
      {stage1_48[197]}
   );
   gpc1_1 gpc5075 (
      {stage0_48[499]},
      {stage1_48[198]}
   );
   gpc1_1 gpc5076 (
      {stage0_48[500]},
      {stage1_48[199]}
   );
   gpc1_1 gpc5077 (
      {stage0_48[501]},
      {stage1_48[200]}
   );
   gpc1_1 gpc5078 (
      {stage0_48[502]},
      {stage1_48[201]}
   );
   gpc1_1 gpc5079 (
      {stage0_48[503]},
      {stage1_48[202]}
   );
   gpc1_1 gpc5080 (
      {stage0_48[504]},
      {stage1_48[203]}
   );
   gpc1_1 gpc5081 (
      {stage0_48[505]},
      {stage1_48[204]}
   );
   gpc1_1 gpc5082 (
      {stage0_48[506]},
      {stage1_48[205]}
   );
   gpc1_1 gpc5083 (
      {stage0_48[507]},
      {stage1_48[206]}
   );
   gpc1_1 gpc5084 (
      {stage0_48[508]},
      {stage1_48[207]}
   );
   gpc1_1 gpc5085 (
      {stage0_48[509]},
      {stage1_48[208]}
   );
   gpc1_1 gpc5086 (
      {stage0_48[510]},
      {stage1_48[209]}
   );
   gpc1_1 gpc5087 (
      {stage0_48[511]},
      {stage1_48[210]}
   );
   gpc1_1 gpc5088 (
      {stage0_49[444]},
      {stage1_49[174]}
   );
   gpc1_1 gpc5089 (
      {stage0_49[445]},
      {stage1_49[175]}
   );
   gpc1_1 gpc5090 (
      {stage0_49[446]},
      {stage1_49[176]}
   );
   gpc1_1 gpc5091 (
      {stage0_49[447]},
      {stage1_49[177]}
   );
   gpc1_1 gpc5092 (
      {stage0_49[448]},
      {stage1_49[178]}
   );
   gpc1_1 gpc5093 (
      {stage0_49[449]},
      {stage1_49[179]}
   );
   gpc1_1 gpc5094 (
      {stage0_49[450]},
      {stage1_49[180]}
   );
   gpc1_1 gpc5095 (
      {stage0_49[451]},
      {stage1_49[181]}
   );
   gpc1_1 gpc5096 (
      {stage0_49[452]},
      {stage1_49[182]}
   );
   gpc1_1 gpc5097 (
      {stage0_49[453]},
      {stage1_49[183]}
   );
   gpc1_1 gpc5098 (
      {stage0_49[454]},
      {stage1_49[184]}
   );
   gpc1_1 gpc5099 (
      {stage0_49[455]},
      {stage1_49[185]}
   );
   gpc1_1 gpc5100 (
      {stage0_49[456]},
      {stage1_49[186]}
   );
   gpc1_1 gpc5101 (
      {stage0_49[457]},
      {stage1_49[187]}
   );
   gpc1_1 gpc5102 (
      {stage0_49[458]},
      {stage1_49[188]}
   );
   gpc1_1 gpc5103 (
      {stage0_49[459]},
      {stage1_49[189]}
   );
   gpc1_1 gpc5104 (
      {stage0_49[460]},
      {stage1_49[190]}
   );
   gpc1_1 gpc5105 (
      {stage0_49[461]},
      {stage1_49[191]}
   );
   gpc1_1 gpc5106 (
      {stage0_49[462]},
      {stage1_49[192]}
   );
   gpc1_1 gpc5107 (
      {stage0_49[463]},
      {stage1_49[193]}
   );
   gpc1_1 gpc5108 (
      {stage0_49[464]},
      {stage1_49[194]}
   );
   gpc1_1 gpc5109 (
      {stage0_49[465]},
      {stage1_49[195]}
   );
   gpc1_1 gpc5110 (
      {stage0_49[466]},
      {stage1_49[196]}
   );
   gpc1_1 gpc5111 (
      {stage0_49[467]},
      {stage1_49[197]}
   );
   gpc1_1 gpc5112 (
      {stage0_49[468]},
      {stage1_49[198]}
   );
   gpc1_1 gpc5113 (
      {stage0_49[469]},
      {stage1_49[199]}
   );
   gpc1_1 gpc5114 (
      {stage0_49[470]},
      {stage1_49[200]}
   );
   gpc1_1 gpc5115 (
      {stage0_49[471]},
      {stage1_49[201]}
   );
   gpc1_1 gpc5116 (
      {stage0_49[472]},
      {stage1_49[202]}
   );
   gpc1_1 gpc5117 (
      {stage0_49[473]},
      {stage1_49[203]}
   );
   gpc1_1 gpc5118 (
      {stage0_49[474]},
      {stage1_49[204]}
   );
   gpc1_1 gpc5119 (
      {stage0_49[475]},
      {stage1_49[205]}
   );
   gpc1_1 gpc5120 (
      {stage0_49[476]},
      {stage1_49[206]}
   );
   gpc1_1 gpc5121 (
      {stage0_49[477]},
      {stage1_49[207]}
   );
   gpc1_1 gpc5122 (
      {stage0_49[478]},
      {stage1_49[208]}
   );
   gpc1_1 gpc5123 (
      {stage0_49[479]},
      {stage1_49[209]}
   );
   gpc1_1 gpc5124 (
      {stage0_49[480]},
      {stage1_49[210]}
   );
   gpc1_1 gpc5125 (
      {stage0_49[481]},
      {stage1_49[211]}
   );
   gpc1_1 gpc5126 (
      {stage0_49[482]},
      {stage1_49[212]}
   );
   gpc1_1 gpc5127 (
      {stage0_49[483]},
      {stage1_49[213]}
   );
   gpc1_1 gpc5128 (
      {stage0_49[484]},
      {stage1_49[214]}
   );
   gpc1_1 gpc5129 (
      {stage0_49[485]},
      {stage1_49[215]}
   );
   gpc1_1 gpc5130 (
      {stage0_49[486]},
      {stage1_49[216]}
   );
   gpc1_1 gpc5131 (
      {stage0_49[487]},
      {stage1_49[217]}
   );
   gpc1_1 gpc5132 (
      {stage0_49[488]},
      {stage1_49[218]}
   );
   gpc1_1 gpc5133 (
      {stage0_49[489]},
      {stage1_49[219]}
   );
   gpc1_1 gpc5134 (
      {stage0_49[490]},
      {stage1_49[220]}
   );
   gpc1_1 gpc5135 (
      {stage0_49[491]},
      {stage1_49[221]}
   );
   gpc1_1 gpc5136 (
      {stage0_49[492]},
      {stage1_49[222]}
   );
   gpc1_1 gpc5137 (
      {stage0_49[493]},
      {stage1_49[223]}
   );
   gpc1_1 gpc5138 (
      {stage0_49[494]},
      {stage1_49[224]}
   );
   gpc1_1 gpc5139 (
      {stage0_49[495]},
      {stage1_49[225]}
   );
   gpc1_1 gpc5140 (
      {stage0_49[496]},
      {stage1_49[226]}
   );
   gpc1_1 gpc5141 (
      {stage0_49[497]},
      {stage1_49[227]}
   );
   gpc1_1 gpc5142 (
      {stage0_49[498]},
      {stage1_49[228]}
   );
   gpc1_1 gpc5143 (
      {stage0_49[499]},
      {stage1_49[229]}
   );
   gpc1_1 gpc5144 (
      {stage0_49[500]},
      {stage1_49[230]}
   );
   gpc1_1 gpc5145 (
      {stage0_49[501]},
      {stage1_49[231]}
   );
   gpc1_1 gpc5146 (
      {stage0_49[502]},
      {stage1_49[232]}
   );
   gpc1_1 gpc5147 (
      {stage0_49[503]},
      {stage1_49[233]}
   );
   gpc1_1 gpc5148 (
      {stage0_49[504]},
      {stage1_49[234]}
   );
   gpc1_1 gpc5149 (
      {stage0_49[505]},
      {stage1_49[235]}
   );
   gpc1_1 gpc5150 (
      {stage0_49[506]},
      {stage1_49[236]}
   );
   gpc1_1 gpc5151 (
      {stage0_49[507]},
      {stage1_49[237]}
   );
   gpc1_1 gpc5152 (
      {stage0_49[508]},
      {stage1_49[238]}
   );
   gpc1_1 gpc5153 (
      {stage0_49[509]},
      {stage1_49[239]}
   );
   gpc1_1 gpc5154 (
      {stage0_49[510]},
      {stage1_49[240]}
   );
   gpc1_1 gpc5155 (
      {stage0_49[511]},
      {stage1_49[241]}
   );
   gpc1_1 gpc5156 (
      {stage0_50[474]},
      {stage1_50[179]}
   );
   gpc1_1 gpc5157 (
      {stage0_50[475]},
      {stage1_50[180]}
   );
   gpc1_1 gpc5158 (
      {stage0_50[476]},
      {stage1_50[181]}
   );
   gpc1_1 gpc5159 (
      {stage0_50[477]},
      {stage1_50[182]}
   );
   gpc1_1 gpc5160 (
      {stage0_50[478]},
      {stage1_50[183]}
   );
   gpc1_1 gpc5161 (
      {stage0_50[479]},
      {stage1_50[184]}
   );
   gpc1_1 gpc5162 (
      {stage0_50[480]},
      {stage1_50[185]}
   );
   gpc1_1 gpc5163 (
      {stage0_50[481]},
      {stage1_50[186]}
   );
   gpc1_1 gpc5164 (
      {stage0_50[482]},
      {stage1_50[187]}
   );
   gpc1_1 gpc5165 (
      {stage0_50[483]},
      {stage1_50[188]}
   );
   gpc1_1 gpc5166 (
      {stage0_50[484]},
      {stage1_50[189]}
   );
   gpc1_1 gpc5167 (
      {stage0_50[485]},
      {stage1_50[190]}
   );
   gpc1_1 gpc5168 (
      {stage0_50[486]},
      {stage1_50[191]}
   );
   gpc1_1 gpc5169 (
      {stage0_50[487]},
      {stage1_50[192]}
   );
   gpc1_1 gpc5170 (
      {stage0_50[488]},
      {stage1_50[193]}
   );
   gpc1_1 gpc5171 (
      {stage0_50[489]},
      {stage1_50[194]}
   );
   gpc1_1 gpc5172 (
      {stage0_50[490]},
      {stage1_50[195]}
   );
   gpc1_1 gpc5173 (
      {stage0_50[491]},
      {stage1_50[196]}
   );
   gpc1_1 gpc5174 (
      {stage0_50[492]},
      {stage1_50[197]}
   );
   gpc1_1 gpc5175 (
      {stage0_50[493]},
      {stage1_50[198]}
   );
   gpc1_1 gpc5176 (
      {stage0_50[494]},
      {stage1_50[199]}
   );
   gpc1_1 gpc5177 (
      {stage0_50[495]},
      {stage1_50[200]}
   );
   gpc1_1 gpc5178 (
      {stage0_50[496]},
      {stage1_50[201]}
   );
   gpc1_1 gpc5179 (
      {stage0_50[497]},
      {stage1_50[202]}
   );
   gpc1_1 gpc5180 (
      {stage0_50[498]},
      {stage1_50[203]}
   );
   gpc1_1 gpc5181 (
      {stage0_50[499]},
      {stage1_50[204]}
   );
   gpc1_1 gpc5182 (
      {stage0_50[500]},
      {stage1_50[205]}
   );
   gpc1_1 gpc5183 (
      {stage0_50[501]},
      {stage1_50[206]}
   );
   gpc1_1 gpc5184 (
      {stage0_50[502]},
      {stage1_50[207]}
   );
   gpc1_1 gpc5185 (
      {stage0_50[503]},
      {stage1_50[208]}
   );
   gpc1_1 gpc5186 (
      {stage0_50[504]},
      {stage1_50[209]}
   );
   gpc1_1 gpc5187 (
      {stage0_50[505]},
      {stage1_50[210]}
   );
   gpc1_1 gpc5188 (
      {stage0_50[506]},
      {stage1_50[211]}
   );
   gpc1_1 gpc5189 (
      {stage0_50[507]},
      {stage1_50[212]}
   );
   gpc1_1 gpc5190 (
      {stage0_50[508]},
      {stage1_50[213]}
   );
   gpc1_1 gpc5191 (
      {stage0_50[509]},
      {stage1_50[214]}
   );
   gpc1_1 gpc5192 (
      {stage0_50[510]},
      {stage1_50[215]}
   );
   gpc1_1 gpc5193 (
      {stage0_50[511]},
      {stage1_50[216]}
   );
   gpc1_1 gpc5194 (
      {stage0_51[501]},
      {stage1_51[216]}
   );
   gpc1_1 gpc5195 (
      {stage0_51[502]},
      {stage1_51[217]}
   );
   gpc1_1 gpc5196 (
      {stage0_51[503]},
      {stage1_51[218]}
   );
   gpc1_1 gpc5197 (
      {stage0_51[504]},
      {stage1_51[219]}
   );
   gpc1_1 gpc5198 (
      {stage0_51[505]},
      {stage1_51[220]}
   );
   gpc1_1 gpc5199 (
      {stage0_51[506]},
      {stage1_51[221]}
   );
   gpc1_1 gpc5200 (
      {stage0_51[507]},
      {stage1_51[222]}
   );
   gpc1_1 gpc5201 (
      {stage0_51[508]},
      {stage1_51[223]}
   );
   gpc1_1 gpc5202 (
      {stage0_51[509]},
      {stage1_51[224]}
   );
   gpc1_1 gpc5203 (
      {stage0_51[510]},
      {stage1_51[225]}
   );
   gpc1_1 gpc5204 (
      {stage0_51[511]},
      {stage1_51[226]}
   );
   gpc1_1 gpc5205 (
      {stage0_52[410]},
      {stage1_52[202]}
   );
   gpc1_1 gpc5206 (
      {stage0_52[411]},
      {stage1_52[203]}
   );
   gpc1_1 gpc5207 (
      {stage0_52[412]},
      {stage1_52[204]}
   );
   gpc1_1 gpc5208 (
      {stage0_52[413]},
      {stage1_52[205]}
   );
   gpc1_1 gpc5209 (
      {stage0_52[414]},
      {stage1_52[206]}
   );
   gpc1_1 gpc5210 (
      {stage0_52[415]},
      {stage1_52[207]}
   );
   gpc1_1 gpc5211 (
      {stage0_52[416]},
      {stage1_52[208]}
   );
   gpc1_1 gpc5212 (
      {stage0_52[417]},
      {stage1_52[209]}
   );
   gpc1_1 gpc5213 (
      {stage0_52[418]},
      {stage1_52[210]}
   );
   gpc1_1 gpc5214 (
      {stage0_52[419]},
      {stage1_52[211]}
   );
   gpc1_1 gpc5215 (
      {stage0_52[420]},
      {stage1_52[212]}
   );
   gpc1_1 gpc5216 (
      {stage0_52[421]},
      {stage1_52[213]}
   );
   gpc1_1 gpc5217 (
      {stage0_52[422]},
      {stage1_52[214]}
   );
   gpc1_1 gpc5218 (
      {stage0_52[423]},
      {stage1_52[215]}
   );
   gpc1_1 gpc5219 (
      {stage0_52[424]},
      {stage1_52[216]}
   );
   gpc1_1 gpc5220 (
      {stage0_52[425]},
      {stage1_52[217]}
   );
   gpc1_1 gpc5221 (
      {stage0_52[426]},
      {stage1_52[218]}
   );
   gpc1_1 gpc5222 (
      {stage0_52[427]},
      {stage1_52[219]}
   );
   gpc1_1 gpc5223 (
      {stage0_52[428]},
      {stage1_52[220]}
   );
   gpc1_1 gpc5224 (
      {stage0_52[429]},
      {stage1_52[221]}
   );
   gpc1_1 gpc5225 (
      {stage0_52[430]},
      {stage1_52[222]}
   );
   gpc1_1 gpc5226 (
      {stage0_52[431]},
      {stage1_52[223]}
   );
   gpc1_1 gpc5227 (
      {stage0_52[432]},
      {stage1_52[224]}
   );
   gpc1_1 gpc5228 (
      {stage0_52[433]},
      {stage1_52[225]}
   );
   gpc1_1 gpc5229 (
      {stage0_52[434]},
      {stage1_52[226]}
   );
   gpc1_1 gpc5230 (
      {stage0_52[435]},
      {stage1_52[227]}
   );
   gpc1_1 gpc5231 (
      {stage0_52[436]},
      {stage1_52[228]}
   );
   gpc1_1 gpc5232 (
      {stage0_52[437]},
      {stage1_52[229]}
   );
   gpc1_1 gpc5233 (
      {stage0_52[438]},
      {stage1_52[230]}
   );
   gpc1_1 gpc5234 (
      {stage0_52[439]},
      {stage1_52[231]}
   );
   gpc1_1 gpc5235 (
      {stage0_52[440]},
      {stage1_52[232]}
   );
   gpc1_1 gpc5236 (
      {stage0_52[441]},
      {stage1_52[233]}
   );
   gpc1_1 gpc5237 (
      {stage0_52[442]},
      {stage1_52[234]}
   );
   gpc1_1 gpc5238 (
      {stage0_52[443]},
      {stage1_52[235]}
   );
   gpc1_1 gpc5239 (
      {stage0_52[444]},
      {stage1_52[236]}
   );
   gpc1_1 gpc5240 (
      {stage0_52[445]},
      {stage1_52[237]}
   );
   gpc1_1 gpc5241 (
      {stage0_52[446]},
      {stage1_52[238]}
   );
   gpc1_1 gpc5242 (
      {stage0_52[447]},
      {stage1_52[239]}
   );
   gpc1_1 gpc5243 (
      {stage0_52[448]},
      {stage1_52[240]}
   );
   gpc1_1 gpc5244 (
      {stage0_52[449]},
      {stage1_52[241]}
   );
   gpc1_1 gpc5245 (
      {stage0_52[450]},
      {stage1_52[242]}
   );
   gpc1_1 gpc5246 (
      {stage0_52[451]},
      {stage1_52[243]}
   );
   gpc1_1 gpc5247 (
      {stage0_52[452]},
      {stage1_52[244]}
   );
   gpc1_1 gpc5248 (
      {stage0_52[453]},
      {stage1_52[245]}
   );
   gpc1_1 gpc5249 (
      {stage0_52[454]},
      {stage1_52[246]}
   );
   gpc1_1 gpc5250 (
      {stage0_52[455]},
      {stage1_52[247]}
   );
   gpc1_1 gpc5251 (
      {stage0_52[456]},
      {stage1_52[248]}
   );
   gpc1_1 gpc5252 (
      {stage0_52[457]},
      {stage1_52[249]}
   );
   gpc1_1 gpc5253 (
      {stage0_52[458]},
      {stage1_52[250]}
   );
   gpc1_1 gpc5254 (
      {stage0_52[459]},
      {stage1_52[251]}
   );
   gpc1_1 gpc5255 (
      {stage0_52[460]},
      {stage1_52[252]}
   );
   gpc1_1 gpc5256 (
      {stage0_52[461]},
      {stage1_52[253]}
   );
   gpc1_1 gpc5257 (
      {stage0_52[462]},
      {stage1_52[254]}
   );
   gpc1_1 gpc5258 (
      {stage0_52[463]},
      {stage1_52[255]}
   );
   gpc1_1 gpc5259 (
      {stage0_52[464]},
      {stage1_52[256]}
   );
   gpc1_1 gpc5260 (
      {stage0_52[465]},
      {stage1_52[257]}
   );
   gpc1_1 gpc5261 (
      {stage0_52[466]},
      {stage1_52[258]}
   );
   gpc1_1 gpc5262 (
      {stage0_52[467]},
      {stage1_52[259]}
   );
   gpc1_1 gpc5263 (
      {stage0_52[468]},
      {stage1_52[260]}
   );
   gpc1_1 gpc5264 (
      {stage0_52[469]},
      {stage1_52[261]}
   );
   gpc1_1 gpc5265 (
      {stage0_52[470]},
      {stage1_52[262]}
   );
   gpc1_1 gpc5266 (
      {stage0_52[471]},
      {stage1_52[263]}
   );
   gpc1_1 gpc5267 (
      {stage0_52[472]},
      {stage1_52[264]}
   );
   gpc1_1 gpc5268 (
      {stage0_52[473]},
      {stage1_52[265]}
   );
   gpc1_1 gpc5269 (
      {stage0_52[474]},
      {stage1_52[266]}
   );
   gpc1_1 gpc5270 (
      {stage0_52[475]},
      {stage1_52[267]}
   );
   gpc1_1 gpc5271 (
      {stage0_52[476]},
      {stage1_52[268]}
   );
   gpc1_1 gpc5272 (
      {stage0_52[477]},
      {stage1_52[269]}
   );
   gpc1_1 gpc5273 (
      {stage0_52[478]},
      {stage1_52[270]}
   );
   gpc1_1 gpc5274 (
      {stage0_52[479]},
      {stage1_52[271]}
   );
   gpc1_1 gpc5275 (
      {stage0_52[480]},
      {stage1_52[272]}
   );
   gpc1_1 gpc5276 (
      {stage0_52[481]},
      {stage1_52[273]}
   );
   gpc1_1 gpc5277 (
      {stage0_52[482]},
      {stage1_52[274]}
   );
   gpc1_1 gpc5278 (
      {stage0_52[483]},
      {stage1_52[275]}
   );
   gpc1_1 gpc5279 (
      {stage0_52[484]},
      {stage1_52[276]}
   );
   gpc1_1 gpc5280 (
      {stage0_52[485]},
      {stage1_52[277]}
   );
   gpc1_1 gpc5281 (
      {stage0_52[486]},
      {stage1_52[278]}
   );
   gpc1_1 gpc5282 (
      {stage0_52[487]},
      {stage1_52[279]}
   );
   gpc1_1 gpc5283 (
      {stage0_52[488]},
      {stage1_52[280]}
   );
   gpc1_1 gpc5284 (
      {stage0_52[489]},
      {stage1_52[281]}
   );
   gpc1_1 gpc5285 (
      {stage0_52[490]},
      {stage1_52[282]}
   );
   gpc1_1 gpc5286 (
      {stage0_52[491]},
      {stage1_52[283]}
   );
   gpc1_1 gpc5287 (
      {stage0_52[492]},
      {stage1_52[284]}
   );
   gpc1_1 gpc5288 (
      {stage0_52[493]},
      {stage1_52[285]}
   );
   gpc1_1 gpc5289 (
      {stage0_52[494]},
      {stage1_52[286]}
   );
   gpc1_1 gpc5290 (
      {stage0_52[495]},
      {stage1_52[287]}
   );
   gpc1_1 gpc5291 (
      {stage0_52[496]},
      {stage1_52[288]}
   );
   gpc1_1 gpc5292 (
      {stage0_52[497]},
      {stage1_52[289]}
   );
   gpc1_1 gpc5293 (
      {stage0_52[498]},
      {stage1_52[290]}
   );
   gpc1_1 gpc5294 (
      {stage0_52[499]},
      {stage1_52[291]}
   );
   gpc1_1 gpc5295 (
      {stage0_52[500]},
      {stage1_52[292]}
   );
   gpc1_1 gpc5296 (
      {stage0_52[501]},
      {stage1_52[293]}
   );
   gpc1_1 gpc5297 (
      {stage0_52[502]},
      {stage1_52[294]}
   );
   gpc1_1 gpc5298 (
      {stage0_52[503]},
      {stage1_52[295]}
   );
   gpc1_1 gpc5299 (
      {stage0_52[504]},
      {stage1_52[296]}
   );
   gpc1_1 gpc5300 (
      {stage0_52[505]},
      {stage1_52[297]}
   );
   gpc1_1 gpc5301 (
      {stage0_52[506]},
      {stage1_52[298]}
   );
   gpc1_1 gpc5302 (
      {stage0_52[507]},
      {stage1_52[299]}
   );
   gpc1_1 gpc5303 (
      {stage0_52[508]},
      {stage1_52[300]}
   );
   gpc1_1 gpc5304 (
      {stage0_52[509]},
      {stage1_52[301]}
   );
   gpc1_1 gpc5305 (
      {stage0_52[510]},
      {stage1_52[302]}
   );
   gpc1_1 gpc5306 (
      {stage0_52[511]},
      {stage1_52[303]}
   );
   gpc1_1 gpc5307 (
      {stage0_53[497]},
      {stage1_53[172]}
   );
   gpc1_1 gpc5308 (
      {stage0_53[498]},
      {stage1_53[173]}
   );
   gpc1_1 gpc5309 (
      {stage0_53[499]},
      {stage1_53[174]}
   );
   gpc1_1 gpc5310 (
      {stage0_53[500]},
      {stage1_53[175]}
   );
   gpc1_1 gpc5311 (
      {stage0_53[501]},
      {stage1_53[176]}
   );
   gpc1_1 gpc5312 (
      {stage0_53[502]},
      {stage1_53[177]}
   );
   gpc1_1 gpc5313 (
      {stage0_53[503]},
      {stage1_53[178]}
   );
   gpc1_1 gpc5314 (
      {stage0_53[504]},
      {stage1_53[179]}
   );
   gpc1_1 gpc5315 (
      {stage0_53[505]},
      {stage1_53[180]}
   );
   gpc1_1 gpc5316 (
      {stage0_53[506]},
      {stage1_53[181]}
   );
   gpc1_1 gpc5317 (
      {stage0_53[507]},
      {stage1_53[182]}
   );
   gpc1_1 gpc5318 (
      {stage0_53[508]},
      {stage1_53[183]}
   );
   gpc1_1 gpc5319 (
      {stage0_53[509]},
      {stage1_53[184]}
   );
   gpc1_1 gpc5320 (
      {stage0_53[510]},
      {stage1_53[185]}
   );
   gpc1_1 gpc5321 (
      {stage0_53[511]},
      {stage1_53[186]}
   );
   gpc1_1 gpc5322 (
      {stage0_54[441]},
      {stage1_54[192]}
   );
   gpc1_1 gpc5323 (
      {stage0_54[442]},
      {stage1_54[193]}
   );
   gpc1_1 gpc5324 (
      {stage0_54[443]},
      {stage1_54[194]}
   );
   gpc1_1 gpc5325 (
      {stage0_54[444]},
      {stage1_54[195]}
   );
   gpc1_1 gpc5326 (
      {stage0_54[445]},
      {stage1_54[196]}
   );
   gpc1_1 gpc5327 (
      {stage0_54[446]},
      {stage1_54[197]}
   );
   gpc1_1 gpc5328 (
      {stage0_54[447]},
      {stage1_54[198]}
   );
   gpc1_1 gpc5329 (
      {stage0_54[448]},
      {stage1_54[199]}
   );
   gpc1_1 gpc5330 (
      {stage0_54[449]},
      {stage1_54[200]}
   );
   gpc1_1 gpc5331 (
      {stage0_54[450]},
      {stage1_54[201]}
   );
   gpc1_1 gpc5332 (
      {stage0_54[451]},
      {stage1_54[202]}
   );
   gpc1_1 gpc5333 (
      {stage0_54[452]},
      {stage1_54[203]}
   );
   gpc1_1 gpc5334 (
      {stage0_54[453]},
      {stage1_54[204]}
   );
   gpc1_1 gpc5335 (
      {stage0_54[454]},
      {stage1_54[205]}
   );
   gpc1_1 gpc5336 (
      {stage0_54[455]},
      {stage1_54[206]}
   );
   gpc1_1 gpc5337 (
      {stage0_54[456]},
      {stage1_54[207]}
   );
   gpc1_1 gpc5338 (
      {stage0_54[457]},
      {stage1_54[208]}
   );
   gpc1_1 gpc5339 (
      {stage0_54[458]},
      {stage1_54[209]}
   );
   gpc1_1 gpc5340 (
      {stage0_54[459]},
      {stage1_54[210]}
   );
   gpc1_1 gpc5341 (
      {stage0_54[460]},
      {stage1_54[211]}
   );
   gpc1_1 gpc5342 (
      {stage0_54[461]},
      {stage1_54[212]}
   );
   gpc1_1 gpc5343 (
      {stage0_54[462]},
      {stage1_54[213]}
   );
   gpc1_1 gpc5344 (
      {stage0_54[463]},
      {stage1_54[214]}
   );
   gpc1_1 gpc5345 (
      {stage0_54[464]},
      {stage1_54[215]}
   );
   gpc1_1 gpc5346 (
      {stage0_54[465]},
      {stage1_54[216]}
   );
   gpc1_1 gpc5347 (
      {stage0_54[466]},
      {stage1_54[217]}
   );
   gpc1_1 gpc5348 (
      {stage0_54[467]},
      {stage1_54[218]}
   );
   gpc1_1 gpc5349 (
      {stage0_54[468]},
      {stage1_54[219]}
   );
   gpc1_1 gpc5350 (
      {stage0_54[469]},
      {stage1_54[220]}
   );
   gpc1_1 gpc5351 (
      {stage0_54[470]},
      {stage1_54[221]}
   );
   gpc1_1 gpc5352 (
      {stage0_54[471]},
      {stage1_54[222]}
   );
   gpc1_1 gpc5353 (
      {stage0_54[472]},
      {stage1_54[223]}
   );
   gpc1_1 gpc5354 (
      {stage0_54[473]},
      {stage1_54[224]}
   );
   gpc1_1 gpc5355 (
      {stage0_54[474]},
      {stage1_54[225]}
   );
   gpc1_1 gpc5356 (
      {stage0_54[475]},
      {stage1_54[226]}
   );
   gpc1_1 gpc5357 (
      {stage0_54[476]},
      {stage1_54[227]}
   );
   gpc1_1 gpc5358 (
      {stage0_54[477]},
      {stage1_54[228]}
   );
   gpc1_1 gpc5359 (
      {stage0_54[478]},
      {stage1_54[229]}
   );
   gpc1_1 gpc5360 (
      {stage0_54[479]},
      {stage1_54[230]}
   );
   gpc1_1 gpc5361 (
      {stage0_54[480]},
      {stage1_54[231]}
   );
   gpc1_1 gpc5362 (
      {stage0_54[481]},
      {stage1_54[232]}
   );
   gpc1_1 gpc5363 (
      {stage0_54[482]},
      {stage1_54[233]}
   );
   gpc1_1 gpc5364 (
      {stage0_54[483]},
      {stage1_54[234]}
   );
   gpc1_1 gpc5365 (
      {stage0_54[484]},
      {stage1_54[235]}
   );
   gpc1_1 gpc5366 (
      {stage0_54[485]},
      {stage1_54[236]}
   );
   gpc1_1 gpc5367 (
      {stage0_54[486]},
      {stage1_54[237]}
   );
   gpc1_1 gpc5368 (
      {stage0_54[487]},
      {stage1_54[238]}
   );
   gpc1_1 gpc5369 (
      {stage0_54[488]},
      {stage1_54[239]}
   );
   gpc1_1 gpc5370 (
      {stage0_54[489]},
      {stage1_54[240]}
   );
   gpc1_1 gpc5371 (
      {stage0_54[490]},
      {stage1_54[241]}
   );
   gpc1_1 gpc5372 (
      {stage0_54[491]},
      {stage1_54[242]}
   );
   gpc1_1 gpc5373 (
      {stage0_54[492]},
      {stage1_54[243]}
   );
   gpc1_1 gpc5374 (
      {stage0_54[493]},
      {stage1_54[244]}
   );
   gpc1_1 gpc5375 (
      {stage0_54[494]},
      {stage1_54[245]}
   );
   gpc1_1 gpc5376 (
      {stage0_54[495]},
      {stage1_54[246]}
   );
   gpc1_1 gpc5377 (
      {stage0_54[496]},
      {stage1_54[247]}
   );
   gpc1_1 gpc5378 (
      {stage0_54[497]},
      {stage1_54[248]}
   );
   gpc1_1 gpc5379 (
      {stage0_54[498]},
      {stage1_54[249]}
   );
   gpc1_1 gpc5380 (
      {stage0_54[499]},
      {stage1_54[250]}
   );
   gpc1_1 gpc5381 (
      {stage0_54[500]},
      {stage1_54[251]}
   );
   gpc1_1 gpc5382 (
      {stage0_54[501]},
      {stage1_54[252]}
   );
   gpc1_1 gpc5383 (
      {stage0_54[502]},
      {stage1_54[253]}
   );
   gpc1_1 gpc5384 (
      {stage0_54[503]},
      {stage1_54[254]}
   );
   gpc1_1 gpc5385 (
      {stage0_54[504]},
      {stage1_54[255]}
   );
   gpc1_1 gpc5386 (
      {stage0_54[505]},
      {stage1_54[256]}
   );
   gpc1_1 gpc5387 (
      {stage0_54[506]},
      {stage1_54[257]}
   );
   gpc1_1 gpc5388 (
      {stage0_54[507]},
      {stage1_54[258]}
   );
   gpc1_1 gpc5389 (
      {stage0_54[508]},
      {stage1_54[259]}
   );
   gpc1_1 gpc5390 (
      {stage0_54[509]},
      {stage1_54[260]}
   );
   gpc1_1 gpc5391 (
      {stage0_54[510]},
      {stage1_54[261]}
   );
   gpc1_1 gpc5392 (
      {stage0_54[511]},
      {stage1_54[262]}
   );
   gpc1_1 gpc5393 (
      {stage0_55[508]},
      {stage1_55[222]}
   );
   gpc1_1 gpc5394 (
      {stage0_55[509]},
      {stage1_55[223]}
   );
   gpc1_1 gpc5395 (
      {stage0_55[510]},
      {stage1_55[224]}
   );
   gpc1_1 gpc5396 (
      {stage0_55[511]},
      {stage1_55[225]}
   );
   gpc1_1 gpc5397 (
      {stage0_56[444]},
      {stage1_56[189]}
   );
   gpc1_1 gpc5398 (
      {stage0_56[445]},
      {stage1_56[190]}
   );
   gpc1_1 gpc5399 (
      {stage0_56[446]},
      {stage1_56[191]}
   );
   gpc1_1 gpc5400 (
      {stage0_56[447]},
      {stage1_56[192]}
   );
   gpc1_1 gpc5401 (
      {stage0_56[448]},
      {stage1_56[193]}
   );
   gpc1_1 gpc5402 (
      {stage0_56[449]},
      {stage1_56[194]}
   );
   gpc1_1 gpc5403 (
      {stage0_56[450]},
      {stage1_56[195]}
   );
   gpc1_1 gpc5404 (
      {stage0_56[451]},
      {stage1_56[196]}
   );
   gpc1_1 gpc5405 (
      {stage0_56[452]},
      {stage1_56[197]}
   );
   gpc1_1 gpc5406 (
      {stage0_56[453]},
      {stage1_56[198]}
   );
   gpc1_1 gpc5407 (
      {stage0_56[454]},
      {stage1_56[199]}
   );
   gpc1_1 gpc5408 (
      {stage0_56[455]},
      {stage1_56[200]}
   );
   gpc1_1 gpc5409 (
      {stage0_56[456]},
      {stage1_56[201]}
   );
   gpc1_1 gpc5410 (
      {stage0_56[457]},
      {stage1_56[202]}
   );
   gpc1_1 gpc5411 (
      {stage0_56[458]},
      {stage1_56[203]}
   );
   gpc1_1 gpc5412 (
      {stage0_56[459]},
      {stage1_56[204]}
   );
   gpc1_1 gpc5413 (
      {stage0_56[460]},
      {stage1_56[205]}
   );
   gpc1_1 gpc5414 (
      {stage0_56[461]},
      {stage1_56[206]}
   );
   gpc1_1 gpc5415 (
      {stage0_56[462]},
      {stage1_56[207]}
   );
   gpc1_1 gpc5416 (
      {stage0_56[463]},
      {stage1_56[208]}
   );
   gpc1_1 gpc5417 (
      {stage0_56[464]},
      {stage1_56[209]}
   );
   gpc1_1 gpc5418 (
      {stage0_56[465]},
      {stage1_56[210]}
   );
   gpc1_1 gpc5419 (
      {stage0_56[466]},
      {stage1_56[211]}
   );
   gpc1_1 gpc5420 (
      {stage0_56[467]},
      {stage1_56[212]}
   );
   gpc1_1 gpc5421 (
      {stage0_56[468]},
      {stage1_56[213]}
   );
   gpc1_1 gpc5422 (
      {stage0_56[469]},
      {stage1_56[214]}
   );
   gpc1_1 gpc5423 (
      {stage0_56[470]},
      {stage1_56[215]}
   );
   gpc1_1 gpc5424 (
      {stage0_56[471]},
      {stage1_56[216]}
   );
   gpc1_1 gpc5425 (
      {stage0_56[472]},
      {stage1_56[217]}
   );
   gpc1_1 gpc5426 (
      {stage0_56[473]},
      {stage1_56[218]}
   );
   gpc1_1 gpc5427 (
      {stage0_56[474]},
      {stage1_56[219]}
   );
   gpc1_1 gpc5428 (
      {stage0_56[475]},
      {stage1_56[220]}
   );
   gpc1_1 gpc5429 (
      {stage0_56[476]},
      {stage1_56[221]}
   );
   gpc1_1 gpc5430 (
      {stage0_56[477]},
      {stage1_56[222]}
   );
   gpc1_1 gpc5431 (
      {stage0_56[478]},
      {stage1_56[223]}
   );
   gpc1_1 gpc5432 (
      {stage0_56[479]},
      {stage1_56[224]}
   );
   gpc1_1 gpc5433 (
      {stage0_56[480]},
      {stage1_56[225]}
   );
   gpc1_1 gpc5434 (
      {stage0_56[481]},
      {stage1_56[226]}
   );
   gpc1_1 gpc5435 (
      {stage0_56[482]},
      {stage1_56[227]}
   );
   gpc1_1 gpc5436 (
      {stage0_56[483]},
      {stage1_56[228]}
   );
   gpc1_1 gpc5437 (
      {stage0_56[484]},
      {stage1_56[229]}
   );
   gpc1_1 gpc5438 (
      {stage0_56[485]},
      {stage1_56[230]}
   );
   gpc1_1 gpc5439 (
      {stage0_56[486]},
      {stage1_56[231]}
   );
   gpc1_1 gpc5440 (
      {stage0_56[487]},
      {stage1_56[232]}
   );
   gpc1_1 gpc5441 (
      {stage0_56[488]},
      {stage1_56[233]}
   );
   gpc1_1 gpc5442 (
      {stage0_56[489]},
      {stage1_56[234]}
   );
   gpc1_1 gpc5443 (
      {stage0_56[490]},
      {stage1_56[235]}
   );
   gpc1_1 gpc5444 (
      {stage0_56[491]},
      {stage1_56[236]}
   );
   gpc1_1 gpc5445 (
      {stage0_56[492]},
      {stage1_56[237]}
   );
   gpc1_1 gpc5446 (
      {stage0_56[493]},
      {stage1_56[238]}
   );
   gpc1_1 gpc5447 (
      {stage0_56[494]},
      {stage1_56[239]}
   );
   gpc1_1 gpc5448 (
      {stage0_56[495]},
      {stage1_56[240]}
   );
   gpc1_1 gpc5449 (
      {stage0_56[496]},
      {stage1_56[241]}
   );
   gpc1_1 gpc5450 (
      {stage0_56[497]},
      {stage1_56[242]}
   );
   gpc1_1 gpc5451 (
      {stage0_56[498]},
      {stage1_56[243]}
   );
   gpc1_1 gpc5452 (
      {stage0_56[499]},
      {stage1_56[244]}
   );
   gpc1_1 gpc5453 (
      {stage0_56[500]},
      {stage1_56[245]}
   );
   gpc1_1 gpc5454 (
      {stage0_56[501]},
      {stage1_56[246]}
   );
   gpc1_1 gpc5455 (
      {stage0_56[502]},
      {stage1_56[247]}
   );
   gpc1_1 gpc5456 (
      {stage0_56[503]},
      {stage1_56[248]}
   );
   gpc1_1 gpc5457 (
      {stage0_56[504]},
      {stage1_56[249]}
   );
   gpc1_1 gpc5458 (
      {stage0_56[505]},
      {stage1_56[250]}
   );
   gpc1_1 gpc5459 (
      {stage0_56[506]},
      {stage1_56[251]}
   );
   gpc1_1 gpc5460 (
      {stage0_56[507]},
      {stage1_56[252]}
   );
   gpc1_1 gpc5461 (
      {stage0_56[508]},
      {stage1_56[253]}
   );
   gpc1_1 gpc5462 (
      {stage0_56[509]},
      {stage1_56[254]}
   );
   gpc1_1 gpc5463 (
      {stage0_56[510]},
      {stage1_56[255]}
   );
   gpc1_1 gpc5464 (
      {stage0_56[511]},
      {stage1_56[256]}
   );
   gpc1_1 gpc5465 (
      {stage0_57[510]},
      {stage1_57[178]}
   );
   gpc1_1 gpc5466 (
      {stage0_57[511]},
      {stage1_57[179]}
   );
   gpc1_1 gpc5467 (
      {stage0_58[493]},
      {stage1_58[224]}
   );
   gpc1_1 gpc5468 (
      {stage0_58[494]},
      {stage1_58[225]}
   );
   gpc1_1 gpc5469 (
      {stage0_58[495]},
      {stage1_58[226]}
   );
   gpc1_1 gpc5470 (
      {stage0_58[496]},
      {stage1_58[227]}
   );
   gpc1_1 gpc5471 (
      {stage0_58[497]},
      {stage1_58[228]}
   );
   gpc1_1 gpc5472 (
      {stage0_58[498]},
      {stage1_58[229]}
   );
   gpc1_1 gpc5473 (
      {stage0_58[499]},
      {stage1_58[230]}
   );
   gpc1_1 gpc5474 (
      {stage0_58[500]},
      {stage1_58[231]}
   );
   gpc1_1 gpc5475 (
      {stage0_58[501]},
      {stage1_58[232]}
   );
   gpc1_1 gpc5476 (
      {stage0_58[502]},
      {stage1_58[233]}
   );
   gpc1_1 gpc5477 (
      {stage0_58[503]},
      {stage1_58[234]}
   );
   gpc1_1 gpc5478 (
      {stage0_58[504]},
      {stage1_58[235]}
   );
   gpc1_1 gpc5479 (
      {stage0_58[505]},
      {stage1_58[236]}
   );
   gpc1_1 gpc5480 (
      {stage0_58[506]},
      {stage1_58[237]}
   );
   gpc1_1 gpc5481 (
      {stage0_58[507]},
      {stage1_58[238]}
   );
   gpc1_1 gpc5482 (
      {stage0_58[508]},
      {stage1_58[239]}
   );
   gpc1_1 gpc5483 (
      {stage0_58[509]},
      {stage1_58[240]}
   );
   gpc1_1 gpc5484 (
      {stage0_58[510]},
      {stage1_58[241]}
   );
   gpc1_1 gpc5485 (
      {stage0_58[511]},
      {stage1_58[242]}
   );
   gpc1_1 gpc5486 (
      {stage0_59[412]},
      {stage1_59[194]}
   );
   gpc1_1 gpc5487 (
      {stage0_59[413]},
      {stage1_59[195]}
   );
   gpc1_1 gpc5488 (
      {stage0_59[414]},
      {stage1_59[196]}
   );
   gpc1_1 gpc5489 (
      {stage0_59[415]},
      {stage1_59[197]}
   );
   gpc1_1 gpc5490 (
      {stage0_59[416]},
      {stage1_59[198]}
   );
   gpc1_1 gpc5491 (
      {stage0_59[417]},
      {stage1_59[199]}
   );
   gpc1_1 gpc5492 (
      {stage0_59[418]},
      {stage1_59[200]}
   );
   gpc1_1 gpc5493 (
      {stage0_59[419]},
      {stage1_59[201]}
   );
   gpc1_1 gpc5494 (
      {stage0_59[420]},
      {stage1_59[202]}
   );
   gpc1_1 gpc5495 (
      {stage0_59[421]},
      {stage1_59[203]}
   );
   gpc1_1 gpc5496 (
      {stage0_59[422]},
      {stage1_59[204]}
   );
   gpc1_1 gpc5497 (
      {stage0_59[423]},
      {stage1_59[205]}
   );
   gpc1_1 gpc5498 (
      {stage0_59[424]},
      {stage1_59[206]}
   );
   gpc1_1 gpc5499 (
      {stage0_59[425]},
      {stage1_59[207]}
   );
   gpc1_1 gpc5500 (
      {stage0_59[426]},
      {stage1_59[208]}
   );
   gpc1_1 gpc5501 (
      {stage0_59[427]},
      {stage1_59[209]}
   );
   gpc1_1 gpc5502 (
      {stage0_59[428]},
      {stage1_59[210]}
   );
   gpc1_1 gpc5503 (
      {stage0_59[429]},
      {stage1_59[211]}
   );
   gpc1_1 gpc5504 (
      {stage0_59[430]},
      {stage1_59[212]}
   );
   gpc1_1 gpc5505 (
      {stage0_59[431]},
      {stage1_59[213]}
   );
   gpc1_1 gpc5506 (
      {stage0_59[432]},
      {stage1_59[214]}
   );
   gpc1_1 gpc5507 (
      {stage0_59[433]},
      {stage1_59[215]}
   );
   gpc1_1 gpc5508 (
      {stage0_59[434]},
      {stage1_59[216]}
   );
   gpc1_1 gpc5509 (
      {stage0_59[435]},
      {stage1_59[217]}
   );
   gpc1_1 gpc5510 (
      {stage0_59[436]},
      {stage1_59[218]}
   );
   gpc1_1 gpc5511 (
      {stage0_59[437]},
      {stage1_59[219]}
   );
   gpc1_1 gpc5512 (
      {stage0_59[438]},
      {stage1_59[220]}
   );
   gpc1_1 gpc5513 (
      {stage0_59[439]},
      {stage1_59[221]}
   );
   gpc1_1 gpc5514 (
      {stage0_59[440]},
      {stage1_59[222]}
   );
   gpc1_1 gpc5515 (
      {stage0_59[441]},
      {stage1_59[223]}
   );
   gpc1_1 gpc5516 (
      {stage0_59[442]},
      {stage1_59[224]}
   );
   gpc1_1 gpc5517 (
      {stage0_59[443]},
      {stage1_59[225]}
   );
   gpc1_1 gpc5518 (
      {stage0_59[444]},
      {stage1_59[226]}
   );
   gpc1_1 gpc5519 (
      {stage0_59[445]},
      {stage1_59[227]}
   );
   gpc1_1 gpc5520 (
      {stage0_59[446]},
      {stage1_59[228]}
   );
   gpc1_1 gpc5521 (
      {stage0_59[447]},
      {stage1_59[229]}
   );
   gpc1_1 gpc5522 (
      {stage0_59[448]},
      {stage1_59[230]}
   );
   gpc1_1 gpc5523 (
      {stage0_59[449]},
      {stage1_59[231]}
   );
   gpc1_1 gpc5524 (
      {stage0_59[450]},
      {stage1_59[232]}
   );
   gpc1_1 gpc5525 (
      {stage0_59[451]},
      {stage1_59[233]}
   );
   gpc1_1 gpc5526 (
      {stage0_59[452]},
      {stage1_59[234]}
   );
   gpc1_1 gpc5527 (
      {stage0_59[453]},
      {stage1_59[235]}
   );
   gpc1_1 gpc5528 (
      {stage0_59[454]},
      {stage1_59[236]}
   );
   gpc1_1 gpc5529 (
      {stage0_59[455]},
      {stage1_59[237]}
   );
   gpc1_1 gpc5530 (
      {stage0_59[456]},
      {stage1_59[238]}
   );
   gpc1_1 gpc5531 (
      {stage0_59[457]},
      {stage1_59[239]}
   );
   gpc1_1 gpc5532 (
      {stage0_59[458]},
      {stage1_59[240]}
   );
   gpc1_1 gpc5533 (
      {stage0_59[459]},
      {stage1_59[241]}
   );
   gpc1_1 gpc5534 (
      {stage0_59[460]},
      {stage1_59[242]}
   );
   gpc1_1 gpc5535 (
      {stage0_59[461]},
      {stage1_59[243]}
   );
   gpc1_1 gpc5536 (
      {stage0_59[462]},
      {stage1_59[244]}
   );
   gpc1_1 gpc5537 (
      {stage0_59[463]},
      {stage1_59[245]}
   );
   gpc1_1 gpc5538 (
      {stage0_59[464]},
      {stage1_59[246]}
   );
   gpc1_1 gpc5539 (
      {stage0_59[465]},
      {stage1_59[247]}
   );
   gpc1_1 gpc5540 (
      {stage0_59[466]},
      {stage1_59[248]}
   );
   gpc1_1 gpc5541 (
      {stage0_59[467]},
      {stage1_59[249]}
   );
   gpc1_1 gpc5542 (
      {stage0_59[468]},
      {stage1_59[250]}
   );
   gpc1_1 gpc5543 (
      {stage0_59[469]},
      {stage1_59[251]}
   );
   gpc1_1 gpc5544 (
      {stage0_59[470]},
      {stage1_59[252]}
   );
   gpc1_1 gpc5545 (
      {stage0_59[471]},
      {stage1_59[253]}
   );
   gpc1_1 gpc5546 (
      {stage0_59[472]},
      {stage1_59[254]}
   );
   gpc1_1 gpc5547 (
      {stage0_59[473]},
      {stage1_59[255]}
   );
   gpc1_1 gpc5548 (
      {stage0_59[474]},
      {stage1_59[256]}
   );
   gpc1_1 gpc5549 (
      {stage0_59[475]},
      {stage1_59[257]}
   );
   gpc1_1 gpc5550 (
      {stage0_59[476]},
      {stage1_59[258]}
   );
   gpc1_1 gpc5551 (
      {stage0_59[477]},
      {stage1_59[259]}
   );
   gpc1_1 gpc5552 (
      {stage0_59[478]},
      {stage1_59[260]}
   );
   gpc1_1 gpc5553 (
      {stage0_59[479]},
      {stage1_59[261]}
   );
   gpc1_1 gpc5554 (
      {stage0_59[480]},
      {stage1_59[262]}
   );
   gpc1_1 gpc5555 (
      {stage0_59[481]},
      {stage1_59[263]}
   );
   gpc1_1 gpc5556 (
      {stage0_59[482]},
      {stage1_59[264]}
   );
   gpc1_1 gpc5557 (
      {stage0_59[483]},
      {stage1_59[265]}
   );
   gpc1_1 gpc5558 (
      {stage0_59[484]},
      {stage1_59[266]}
   );
   gpc1_1 gpc5559 (
      {stage0_59[485]},
      {stage1_59[267]}
   );
   gpc1_1 gpc5560 (
      {stage0_59[486]},
      {stage1_59[268]}
   );
   gpc1_1 gpc5561 (
      {stage0_59[487]},
      {stage1_59[269]}
   );
   gpc1_1 gpc5562 (
      {stage0_59[488]},
      {stage1_59[270]}
   );
   gpc1_1 gpc5563 (
      {stage0_59[489]},
      {stage1_59[271]}
   );
   gpc1_1 gpc5564 (
      {stage0_59[490]},
      {stage1_59[272]}
   );
   gpc1_1 gpc5565 (
      {stage0_59[491]},
      {stage1_59[273]}
   );
   gpc1_1 gpc5566 (
      {stage0_59[492]},
      {stage1_59[274]}
   );
   gpc1_1 gpc5567 (
      {stage0_59[493]},
      {stage1_59[275]}
   );
   gpc1_1 gpc5568 (
      {stage0_59[494]},
      {stage1_59[276]}
   );
   gpc1_1 gpc5569 (
      {stage0_59[495]},
      {stage1_59[277]}
   );
   gpc1_1 gpc5570 (
      {stage0_59[496]},
      {stage1_59[278]}
   );
   gpc1_1 gpc5571 (
      {stage0_59[497]},
      {stage1_59[279]}
   );
   gpc1_1 gpc5572 (
      {stage0_59[498]},
      {stage1_59[280]}
   );
   gpc1_1 gpc5573 (
      {stage0_59[499]},
      {stage1_59[281]}
   );
   gpc1_1 gpc5574 (
      {stage0_59[500]},
      {stage1_59[282]}
   );
   gpc1_1 gpc5575 (
      {stage0_59[501]},
      {stage1_59[283]}
   );
   gpc1_1 gpc5576 (
      {stage0_59[502]},
      {stage1_59[284]}
   );
   gpc1_1 gpc5577 (
      {stage0_59[503]},
      {stage1_59[285]}
   );
   gpc1_1 gpc5578 (
      {stage0_59[504]},
      {stage1_59[286]}
   );
   gpc1_1 gpc5579 (
      {stage0_59[505]},
      {stage1_59[287]}
   );
   gpc1_1 gpc5580 (
      {stage0_59[506]},
      {stage1_59[288]}
   );
   gpc1_1 gpc5581 (
      {stage0_59[507]},
      {stage1_59[289]}
   );
   gpc1_1 gpc5582 (
      {stage0_59[508]},
      {stage1_59[290]}
   );
   gpc1_1 gpc5583 (
      {stage0_59[509]},
      {stage1_59[291]}
   );
   gpc1_1 gpc5584 (
      {stage0_59[510]},
      {stage1_59[292]}
   );
   gpc1_1 gpc5585 (
      {stage0_59[511]},
      {stage1_59[293]}
   );
   gpc1_1 gpc5586 (
      {stage0_60[502]},
      {stage1_60[190]}
   );
   gpc1_1 gpc5587 (
      {stage0_60[503]},
      {stage1_60[191]}
   );
   gpc1_1 gpc5588 (
      {stage0_60[504]},
      {stage1_60[192]}
   );
   gpc1_1 gpc5589 (
      {stage0_60[505]},
      {stage1_60[193]}
   );
   gpc1_1 gpc5590 (
      {stage0_60[506]},
      {stage1_60[194]}
   );
   gpc1_1 gpc5591 (
      {stage0_60[507]},
      {stage1_60[195]}
   );
   gpc1_1 gpc5592 (
      {stage0_60[508]},
      {stage1_60[196]}
   );
   gpc1_1 gpc5593 (
      {stage0_60[509]},
      {stage1_60[197]}
   );
   gpc1_1 gpc5594 (
      {stage0_60[510]},
      {stage1_60[198]}
   );
   gpc1_1 gpc5595 (
      {stage0_60[511]},
      {stage1_60[199]}
   );
   gpc1_1 gpc5596 (
      {stage0_62[330]},
      {stage1_62[191]}
   );
   gpc1_1 gpc5597 (
      {stage0_62[331]},
      {stage1_62[192]}
   );
   gpc1_1 gpc5598 (
      {stage0_62[332]},
      {stage1_62[193]}
   );
   gpc1_1 gpc5599 (
      {stage0_62[333]},
      {stage1_62[194]}
   );
   gpc1_1 gpc5600 (
      {stage0_62[334]},
      {stage1_62[195]}
   );
   gpc1_1 gpc5601 (
      {stage0_62[335]},
      {stage1_62[196]}
   );
   gpc1_1 gpc5602 (
      {stage0_62[336]},
      {stage1_62[197]}
   );
   gpc1_1 gpc5603 (
      {stage0_62[337]},
      {stage1_62[198]}
   );
   gpc1_1 gpc5604 (
      {stage0_62[338]},
      {stage1_62[199]}
   );
   gpc1_1 gpc5605 (
      {stage0_62[339]},
      {stage1_62[200]}
   );
   gpc1_1 gpc5606 (
      {stage0_62[340]},
      {stage1_62[201]}
   );
   gpc1_1 gpc5607 (
      {stage0_62[341]},
      {stage1_62[202]}
   );
   gpc1_1 gpc5608 (
      {stage0_62[342]},
      {stage1_62[203]}
   );
   gpc1_1 gpc5609 (
      {stage0_62[343]},
      {stage1_62[204]}
   );
   gpc1_1 gpc5610 (
      {stage0_62[344]},
      {stage1_62[205]}
   );
   gpc1_1 gpc5611 (
      {stage0_62[345]},
      {stage1_62[206]}
   );
   gpc1_1 gpc5612 (
      {stage0_62[346]},
      {stage1_62[207]}
   );
   gpc1_1 gpc5613 (
      {stage0_62[347]},
      {stage1_62[208]}
   );
   gpc1_1 gpc5614 (
      {stage0_62[348]},
      {stage1_62[209]}
   );
   gpc1_1 gpc5615 (
      {stage0_62[349]},
      {stage1_62[210]}
   );
   gpc1_1 gpc5616 (
      {stage0_62[350]},
      {stage1_62[211]}
   );
   gpc1_1 gpc5617 (
      {stage0_62[351]},
      {stage1_62[212]}
   );
   gpc1_1 gpc5618 (
      {stage0_62[352]},
      {stage1_62[213]}
   );
   gpc1_1 gpc5619 (
      {stage0_62[353]},
      {stage1_62[214]}
   );
   gpc1_1 gpc5620 (
      {stage0_62[354]},
      {stage1_62[215]}
   );
   gpc1_1 gpc5621 (
      {stage0_62[355]},
      {stage1_62[216]}
   );
   gpc1_1 gpc5622 (
      {stage0_62[356]},
      {stage1_62[217]}
   );
   gpc1_1 gpc5623 (
      {stage0_62[357]},
      {stage1_62[218]}
   );
   gpc1_1 gpc5624 (
      {stage0_62[358]},
      {stage1_62[219]}
   );
   gpc1_1 gpc5625 (
      {stage0_62[359]},
      {stage1_62[220]}
   );
   gpc1_1 gpc5626 (
      {stage0_62[360]},
      {stage1_62[221]}
   );
   gpc1_1 gpc5627 (
      {stage0_62[361]},
      {stage1_62[222]}
   );
   gpc1_1 gpc5628 (
      {stage0_62[362]},
      {stage1_62[223]}
   );
   gpc1_1 gpc5629 (
      {stage0_62[363]},
      {stage1_62[224]}
   );
   gpc1_1 gpc5630 (
      {stage0_62[364]},
      {stage1_62[225]}
   );
   gpc1_1 gpc5631 (
      {stage0_62[365]},
      {stage1_62[226]}
   );
   gpc1_1 gpc5632 (
      {stage0_62[366]},
      {stage1_62[227]}
   );
   gpc1_1 gpc5633 (
      {stage0_62[367]},
      {stage1_62[228]}
   );
   gpc1_1 gpc5634 (
      {stage0_62[368]},
      {stage1_62[229]}
   );
   gpc1_1 gpc5635 (
      {stage0_62[369]},
      {stage1_62[230]}
   );
   gpc1_1 gpc5636 (
      {stage0_62[370]},
      {stage1_62[231]}
   );
   gpc1_1 gpc5637 (
      {stage0_62[371]},
      {stage1_62[232]}
   );
   gpc1_1 gpc5638 (
      {stage0_62[372]},
      {stage1_62[233]}
   );
   gpc1_1 gpc5639 (
      {stage0_62[373]},
      {stage1_62[234]}
   );
   gpc1_1 gpc5640 (
      {stage0_62[374]},
      {stage1_62[235]}
   );
   gpc1_1 gpc5641 (
      {stage0_62[375]},
      {stage1_62[236]}
   );
   gpc1_1 gpc5642 (
      {stage0_62[376]},
      {stage1_62[237]}
   );
   gpc1_1 gpc5643 (
      {stage0_62[377]},
      {stage1_62[238]}
   );
   gpc1_1 gpc5644 (
      {stage0_62[378]},
      {stage1_62[239]}
   );
   gpc1_1 gpc5645 (
      {stage0_62[379]},
      {stage1_62[240]}
   );
   gpc1_1 gpc5646 (
      {stage0_62[380]},
      {stage1_62[241]}
   );
   gpc1_1 gpc5647 (
      {stage0_62[381]},
      {stage1_62[242]}
   );
   gpc1_1 gpc5648 (
      {stage0_62[382]},
      {stage1_62[243]}
   );
   gpc1_1 gpc5649 (
      {stage0_62[383]},
      {stage1_62[244]}
   );
   gpc1_1 gpc5650 (
      {stage0_62[384]},
      {stage1_62[245]}
   );
   gpc1_1 gpc5651 (
      {stage0_62[385]},
      {stage1_62[246]}
   );
   gpc1_1 gpc5652 (
      {stage0_62[386]},
      {stage1_62[247]}
   );
   gpc1_1 gpc5653 (
      {stage0_62[387]},
      {stage1_62[248]}
   );
   gpc1_1 gpc5654 (
      {stage0_62[388]},
      {stage1_62[249]}
   );
   gpc1_1 gpc5655 (
      {stage0_62[389]},
      {stage1_62[250]}
   );
   gpc1_1 gpc5656 (
      {stage0_62[390]},
      {stage1_62[251]}
   );
   gpc1_1 gpc5657 (
      {stage0_62[391]},
      {stage1_62[252]}
   );
   gpc1_1 gpc5658 (
      {stage0_62[392]},
      {stage1_62[253]}
   );
   gpc1_1 gpc5659 (
      {stage0_62[393]},
      {stage1_62[254]}
   );
   gpc1_1 gpc5660 (
      {stage0_62[394]},
      {stage1_62[255]}
   );
   gpc1_1 gpc5661 (
      {stage0_62[395]},
      {stage1_62[256]}
   );
   gpc1_1 gpc5662 (
      {stage0_62[396]},
      {stage1_62[257]}
   );
   gpc1_1 gpc5663 (
      {stage0_62[397]},
      {stage1_62[258]}
   );
   gpc1_1 gpc5664 (
      {stage0_62[398]},
      {stage1_62[259]}
   );
   gpc1_1 gpc5665 (
      {stage0_62[399]},
      {stage1_62[260]}
   );
   gpc1_1 gpc5666 (
      {stage0_62[400]},
      {stage1_62[261]}
   );
   gpc1_1 gpc5667 (
      {stage0_62[401]},
      {stage1_62[262]}
   );
   gpc1_1 gpc5668 (
      {stage0_62[402]},
      {stage1_62[263]}
   );
   gpc1_1 gpc5669 (
      {stage0_62[403]},
      {stage1_62[264]}
   );
   gpc1_1 gpc5670 (
      {stage0_62[404]},
      {stage1_62[265]}
   );
   gpc1_1 gpc5671 (
      {stage0_62[405]},
      {stage1_62[266]}
   );
   gpc1_1 gpc5672 (
      {stage0_62[406]},
      {stage1_62[267]}
   );
   gpc1_1 gpc5673 (
      {stage0_62[407]},
      {stage1_62[268]}
   );
   gpc1_1 gpc5674 (
      {stage0_62[408]},
      {stage1_62[269]}
   );
   gpc1_1 gpc5675 (
      {stage0_62[409]},
      {stage1_62[270]}
   );
   gpc1_1 gpc5676 (
      {stage0_62[410]},
      {stage1_62[271]}
   );
   gpc1_1 gpc5677 (
      {stage0_62[411]},
      {stage1_62[272]}
   );
   gpc1_1 gpc5678 (
      {stage0_62[412]},
      {stage1_62[273]}
   );
   gpc1_1 gpc5679 (
      {stage0_62[413]},
      {stage1_62[274]}
   );
   gpc1_1 gpc5680 (
      {stage0_62[414]},
      {stage1_62[275]}
   );
   gpc1_1 gpc5681 (
      {stage0_62[415]},
      {stage1_62[276]}
   );
   gpc1_1 gpc5682 (
      {stage0_62[416]},
      {stage1_62[277]}
   );
   gpc1_1 gpc5683 (
      {stage0_62[417]},
      {stage1_62[278]}
   );
   gpc1_1 gpc5684 (
      {stage0_62[418]},
      {stage1_62[279]}
   );
   gpc1_1 gpc5685 (
      {stage0_62[419]},
      {stage1_62[280]}
   );
   gpc1_1 gpc5686 (
      {stage0_62[420]},
      {stage1_62[281]}
   );
   gpc1_1 gpc5687 (
      {stage0_62[421]},
      {stage1_62[282]}
   );
   gpc1_1 gpc5688 (
      {stage0_62[422]},
      {stage1_62[283]}
   );
   gpc1_1 gpc5689 (
      {stage0_62[423]},
      {stage1_62[284]}
   );
   gpc1_1 gpc5690 (
      {stage0_62[424]},
      {stage1_62[285]}
   );
   gpc1_1 gpc5691 (
      {stage0_62[425]},
      {stage1_62[286]}
   );
   gpc1_1 gpc5692 (
      {stage0_62[426]},
      {stage1_62[287]}
   );
   gpc1_1 gpc5693 (
      {stage0_62[427]},
      {stage1_62[288]}
   );
   gpc1_1 gpc5694 (
      {stage0_62[428]},
      {stage1_62[289]}
   );
   gpc1_1 gpc5695 (
      {stage0_62[429]},
      {stage1_62[290]}
   );
   gpc1_1 gpc5696 (
      {stage0_62[430]},
      {stage1_62[291]}
   );
   gpc1_1 gpc5697 (
      {stage0_62[431]},
      {stage1_62[292]}
   );
   gpc1_1 gpc5698 (
      {stage0_62[432]},
      {stage1_62[293]}
   );
   gpc1_1 gpc5699 (
      {stage0_62[433]},
      {stage1_62[294]}
   );
   gpc1_1 gpc5700 (
      {stage0_62[434]},
      {stage1_62[295]}
   );
   gpc1_1 gpc5701 (
      {stage0_62[435]},
      {stage1_62[296]}
   );
   gpc1_1 gpc5702 (
      {stage0_62[436]},
      {stage1_62[297]}
   );
   gpc1_1 gpc5703 (
      {stage0_62[437]},
      {stage1_62[298]}
   );
   gpc1_1 gpc5704 (
      {stage0_62[438]},
      {stage1_62[299]}
   );
   gpc1_1 gpc5705 (
      {stage0_62[439]},
      {stage1_62[300]}
   );
   gpc1_1 gpc5706 (
      {stage0_62[440]},
      {stage1_62[301]}
   );
   gpc1_1 gpc5707 (
      {stage0_62[441]},
      {stage1_62[302]}
   );
   gpc1_1 gpc5708 (
      {stage0_62[442]},
      {stage1_62[303]}
   );
   gpc1_1 gpc5709 (
      {stage0_62[443]},
      {stage1_62[304]}
   );
   gpc1_1 gpc5710 (
      {stage0_62[444]},
      {stage1_62[305]}
   );
   gpc1_1 gpc5711 (
      {stage0_62[445]},
      {stage1_62[306]}
   );
   gpc1_1 gpc5712 (
      {stage0_62[446]},
      {stage1_62[307]}
   );
   gpc1_1 gpc5713 (
      {stage0_62[447]},
      {stage1_62[308]}
   );
   gpc1_1 gpc5714 (
      {stage0_62[448]},
      {stage1_62[309]}
   );
   gpc1_1 gpc5715 (
      {stage0_62[449]},
      {stage1_62[310]}
   );
   gpc1_1 gpc5716 (
      {stage0_62[450]},
      {stage1_62[311]}
   );
   gpc1_1 gpc5717 (
      {stage0_62[451]},
      {stage1_62[312]}
   );
   gpc1_1 gpc5718 (
      {stage0_62[452]},
      {stage1_62[313]}
   );
   gpc1_1 gpc5719 (
      {stage0_62[453]},
      {stage1_62[314]}
   );
   gpc1_1 gpc5720 (
      {stage0_62[454]},
      {stage1_62[315]}
   );
   gpc1_1 gpc5721 (
      {stage0_62[455]},
      {stage1_62[316]}
   );
   gpc1_1 gpc5722 (
      {stage0_62[456]},
      {stage1_62[317]}
   );
   gpc1_1 gpc5723 (
      {stage0_62[457]},
      {stage1_62[318]}
   );
   gpc1_1 gpc5724 (
      {stage0_62[458]},
      {stage1_62[319]}
   );
   gpc1_1 gpc5725 (
      {stage0_62[459]},
      {stage1_62[320]}
   );
   gpc1_1 gpc5726 (
      {stage0_62[460]},
      {stage1_62[321]}
   );
   gpc1_1 gpc5727 (
      {stage0_62[461]},
      {stage1_62[322]}
   );
   gpc1_1 gpc5728 (
      {stage0_62[462]},
      {stage1_62[323]}
   );
   gpc1_1 gpc5729 (
      {stage0_62[463]},
      {stage1_62[324]}
   );
   gpc1_1 gpc5730 (
      {stage0_62[464]},
      {stage1_62[325]}
   );
   gpc1_1 gpc5731 (
      {stage0_62[465]},
      {stage1_62[326]}
   );
   gpc1_1 gpc5732 (
      {stage0_62[466]},
      {stage1_62[327]}
   );
   gpc1_1 gpc5733 (
      {stage0_62[467]},
      {stage1_62[328]}
   );
   gpc1_1 gpc5734 (
      {stage0_62[468]},
      {stage1_62[329]}
   );
   gpc1_1 gpc5735 (
      {stage0_62[469]},
      {stage1_62[330]}
   );
   gpc1_1 gpc5736 (
      {stage0_62[470]},
      {stage1_62[331]}
   );
   gpc1_1 gpc5737 (
      {stage0_62[471]},
      {stage1_62[332]}
   );
   gpc1_1 gpc5738 (
      {stage0_62[472]},
      {stage1_62[333]}
   );
   gpc1_1 gpc5739 (
      {stage0_62[473]},
      {stage1_62[334]}
   );
   gpc1_1 gpc5740 (
      {stage0_62[474]},
      {stage1_62[335]}
   );
   gpc1_1 gpc5741 (
      {stage0_62[475]},
      {stage1_62[336]}
   );
   gpc1_1 gpc5742 (
      {stage0_62[476]},
      {stage1_62[337]}
   );
   gpc1_1 gpc5743 (
      {stage0_62[477]},
      {stage1_62[338]}
   );
   gpc1_1 gpc5744 (
      {stage0_62[478]},
      {stage1_62[339]}
   );
   gpc1_1 gpc5745 (
      {stage0_62[479]},
      {stage1_62[340]}
   );
   gpc1_1 gpc5746 (
      {stage0_62[480]},
      {stage1_62[341]}
   );
   gpc1_1 gpc5747 (
      {stage0_62[481]},
      {stage1_62[342]}
   );
   gpc1_1 gpc5748 (
      {stage0_62[482]},
      {stage1_62[343]}
   );
   gpc1_1 gpc5749 (
      {stage0_62[483]},
      {stage1_62[344]}
   );
   gpc1_1 gpc5750 (
      {stage0_62[484]},
      {stage1_62[345]}
   );
   gpc1_1 gpc5751 (
      {stage0_62[485]},
      {stage1_62[346]}
   );
   gpc1_1 gpc5752 (
      {stage0_62[486]},
      {stage1_62[347]}
   );
   gpc1_1 gpc5753 (
      {stage0_62[487]},
      {stage1_62[348]}
   );
   gpc1_1 gpc5754 (
      {stage0_62[488]},
      {stage1_62[349]}
   );
   gpc1_1 gpc5755 (
      {stage0_62[489]},
      {stage1_62[350]}
   );
   gpc1_1 gpc5756 (
      {stage0_62[490]},
      {stage1_62[351]}
   );
   gpc1_1 gpc5757 (
      {stage0_62[491]},
      {stage1_62[352]}
   );
   gpc1_1 gpc5758 (
      {stage0_62[492]},
      {stage1_62[353]}
   );
   gpc1_1 gpc5759 (
      {stage0_62[493]},
      {stage1_62[354]}
   );
   gpc1_1 gpc5760 (
      {stage0_62[494]},
      {stage1_62[355]}
   );
   gpc1_1 gpc5761 (
      {stage0_62[495]},
      {stage1_62[356]}
   );
   gpc1_1 gpc5762 (
      {stage0_62[496]},
      {stage1_62[357]}
   );
   gpc1_1 gpc5763 (
      {stage0_62[497]},
      {stage1_62[358]}
   );
   gpc1_1 gpc5764 (
      {stage0_62[498]},
      {stage1_62[359]}
   );
   gpc1_1 gpc5765 (
      {stage0_62[499]},
      {stage1_62[360]}
   );
   gpc1_1 gpc5766 (
      {stage0_62[500]},
      {stage1_62[361]}
   );
   gpc1_1 gpc5767 (
      {stage0_62[501]},
      {stage1_62[362]}
   );
   gpc1_1 gpc5768 (
      {stage0_62[502]},
      {stage1_62[363]}
   );
   gpc1_1 gpc5769 (
      {stage0_62[503]},
      {stage1_62[364]}
   );
   gpc1_1 gpc5770 (
      {stage0_62[504]},
      {stage1_62[365]}
   );
   gpc1_1 gpc5771 (
      {stage0_62[505]},
      {stage1_62[366]}
   );
   gpc1_1 gpc5772 (
      {stage0_62[506]},
      {stage1_62[367]}
   );
   gpc1_1 gpc5773 (
      {stage0_62[507]},
      {stage1_62[368]}
   );
   gpc1_1 gpc5774 (
      {stage0_62[508]},
      {stage1_62[369]}
   );
   gpc1_1 gpc5775 (
      {stage0_62[509]},
      {stage1_62[370]}
   );
   gpc1_1 gpc5776 (
      {stage0_62[510]},
      {stage1_62[371]}
   );
   gpc1_1 gpc5777 (
      {stage0_62[511]},
      {stage1_62[372]}
   );
   gpc1_1 gpc5778 (
      {stage0_63[342]},
      {stage1_63[125]}
   );
   gpc1_1 gpc5779 (
      {stage0_63[343]},
      {stage1_63[126]}
   );
   gpc1_1 gpc5780 (
      {stage0_63[344]},
      {stage1_63[127]}
   );
   gpc1_1 gpc5781 (
      {stage0_63[345]},
      {stage1_63[128]}
   );
   gpc1_1 gpc5782 (
      {stage0_63[346]},
      {stage1_63[129]}
   );
   gpc1_1 gpc5783 (
      {stage0_63[347]},
      {stage1_63[130]}
   );
   gpc1_1 gpc5784 (
      {stage0_63[348]},
      {stage1_63[131]}
   );
   gpc1_1 gpc5785 (
      {stage0_63[349]},
      {stage1_63[132]}
   );
   gpc1_1 gpc5786 (
      {stage0_63[350]},
      {stage1_63[133]}
   );
   gpc1_1 gpc5787 (
      {stage0_63[351]},
      {stage1_63[134]}
   );
   gpc1_1 gpc5788 (
      {stage0_63[352]},
      {stage1_63[135]}
   );
   gpc1_1 gpc5789 (
      {stage0_63[353]},
      {stage1_63[136]}
   );
   gpc1_1 gpc5790 (
      {stage0_63[354]},
      {stage1_63[137]}
   );
   gpc1_1 gpc5791 (
      {stage0_63[355]},
      {stage1_63[138]}
   );
   gpc1_1 gpc5792 (
      {stage0_63[356]},
      {stage1_63[139]}
   );
   gpc1_1 gpc5793 (
      {stage0_63[357]},
      {stage1_63[140]}
   );
   gpc1_1 gpc5794 (
      {stage0_63[358]},
      {stage1_63[141]}
   );
   gpc1_1 gpc5795 (
      {stage0_63[359]},
      {stage1_63[142]}
   );
   gpc1_1 gpc5796 (
      {stage0_63[360]},
      {stage1_63[143]}
   );
   gpc1_1 gpc5797 (
      {stage0_63[361]},
      {stage1_63[144]}
   );
   gpc1_1 gpc5798 (
      {stage0_63[362]},
      {stage1_63[145]}
   );
   gpc1_1 gpc5799 (
      {stage0_63[363]},
      {stage1_63[146]}
   );
   gpc1_1 gpc5800 (
      {stage0_63[364]},
      {stage1_63[147]}
   );
   gpc1_1 gpc5801 (
      {stage0_63[365]},
      {stage1_63[148]}
   );
   gpc1_1 gpc5802 (
      {stage0_63[366]},
      {stage1_63[149]}
   );
   gpc1_1 gpc5803 (
      {stage0_63[367]},
      {stage1_63[150]}
   );
   gpc1_1 gpc5804 (
      {stage0_63[368]},
      {stage1_63[151]}
   );
   gpc1_1 gpc5805 (
      {stage0_63[369]},
      {stage1_63[152]}
   );
   gpc1_1 gpc5806 (
      {stage0_63[370]},
      {stage1_63[153]}
   );
   gpc1_1 gpc5807 (
      {stage0_63[371]},
      {stage1_63[154]}
   );
   gpc1_1 gpc5808 (
      {stage0_63[372]},
      {stage1_63[155]}
   );
   gpc1_1 gpc5809 (
      {stage0_63[373]},
      {stage1_63[156]}
   );
   gpc1_1 gpc5810 (
      {stage0_63[374]},
      {stage1_63[157]}
   );
   gpc1_1 gpc5811 (
      {stage0_63[375]},
      {stage1_63[158]}
   );
   gpc1_1 gpc5812 (
      {stage0_63[376]},
      {stage1_63[159]}
   );
   gpc1_1 gpc5813 (
      {stage0_63[377]},
      {stage1_63[160]}
   );
   gpc1_1 gpc5814 (
      {stage0_63[378]},
      {stage1_63[161]}
   );
   gpc1_1 gpc5815 (
      {stage0_63[379]},
      {stage1_63[162]}
   );
   gpc1_1 gpc5816 (
      {stage0_63[380]},
      {stage1_63[163]}
   );
   gpc1_1 gpc5817 (
      {stage0_63[381]},
      {stage1_63[164]}
   );
   gpc1_1 gpc5818 (
      {stage0_63[382]},
      {stage1_63[165]}
   );
   gpc1_1 gpc5819 (
      {stage0_63[383]},
      {stage1_63[166]}
   );
   gpc1_1 gpc5820 (
      {stage0_63[384]},
      {stage1_63[167]}
   );
   gpc1_1 gpc5821 (
      {stage0_63[385]},
      {stage1_63[168]}
   );
   gpc1_1 gpc5822 (
      {stage0_63[386]},
      {stage1_63[169]}
   );
   gpc1_1 gpc5823 (
      {stage0_63[387]},
      {stage1_63[170]}
   );
   gpc1_1 gpc5824 (
      {stage0_63[388]},
      {stage1_63[171]}
   );
   gpc1_1 gpc5825 (
      {stage0_63[389]},
      {stage1_63[172]}
   );
   gpc1_1 gpc5826 (
      {stage0_63[390]},
      {stage1_63[173]}
   );
   gpc1_1 gpc5827 (
      {stage0_63[391]},
      {stage1_63[174]}
   );
   gpc1_1 gpc5828 (
      {stage0_63[392]},
      {stage1_63[175]}
   );
   gpc1_1 gpc5829 (
      {stage0_63[393]},
      {stage1_63[176]}
   );
   gpc1_1 gpc5830 (
      {stage0_63[394]},
      {stage1_63[177]}
   );
   gpc1_1 gpc5831 (
      {stage0_63[395]},
      {stage1_63[178]}
   );
   gpc1_1 gpc5832 (
      {stage0_63[396]},
      {stage1_63[179]}
   );
   gpc1_1 gpc5833 (
      {stage0_63[397]},
      {stage1_63[180]}
   );
   gpc1_1 gpc5834 (
      {stage0_63[398]},
      {stage1_63[181]}
   );
   gpc1_1 gpc5835 (
      {stage0_63[399]},
      {stage1_63[182]}
   );
   gpc1_1 gpc5836 (
      {stage0_63[400]},
      {stage1_63[183]}
   );
   gpc1_1 gpc5837 (
      {stage0_63[401]},
      {stage1_63[184]}
   );
   gpc1_1 gpc5838 (
      {stage0_63[402]},
      {stage1_63[185]}
   );
   gpc1_1 gpc5839 (
      {stage0_63[403]},
      {stage1_63[186]}
   );
   gpc1_1 gpc5840 (
      {stage0_63[404]},
      {stage1_63[187]}
   );
   gpc1_1 gpc5841 (
      {stage0_63[405]},
      {stage1_63[188]}
   );
   gpc1_1 gpc5842 (
      {stage0_63[406]},
      {stage1_63[189]}
   );
   gpc1_1 gpc5843 (
      {stage0_63[407]},
      {stage1_63[190]}
   );
   gpc1_1 gpc5844 (
      {stage0_63[408]},
      {stage1_63[191]}
   );
   gpc1_1 gpc5845 (
      {stage0_63[409]},
      {stage1_63[192]}
   );
   gpc1_1 gpc5846 (
      {stage0_63[410]},
      {stage1_63[193]}
   );
   gpc1_1 gpc5847 (
      {stage0_63[411]},
      {stage1_63[194]}
   );
   gpc1_1 gpc5848 (
      {stage0_63[412]},
      {stage1_63[195]}
   );
   gpc1_1 gpc5849 (
      {stage0_63[413]},
      {stage1_63[196]}
   );
   gpc1_1 gpc5850 (
      {stage0_63[414]},
      {stage1_63[197]}
   );
   gpc1_1 gpc5851 (
      {stage0_63[415]},
      {stage1_63[198]}
   );
   gpc1_1 gpc5852 (
      {stage0_63[416]},
      {stage1_63[199]}
   );
   gpc1_1 gpc5853 (
      {stage0_63[417]},
      {stage1_63[200]}
   );
   gpc1_1 gpc5854 (
      {stage0_63[418]},
      {stage1_63[201]}
   );
   gpc1_1 gpc5855 (
      {stage0_63[419]},
      {stage1_63[202]}
   );
   gpc1_1 gpc5856 (
      {stage0_63[420]},
      {stage1_63[203]}
   );
   gpc1_1 gpc5857 (
      {stage0_63[421]},
      {stage1_63[204]}
   );
   gpc1_1 gpc5858 (
      {stage0_63[422]},
      {stage1_63[205]}
   );
   gpc1_1 gpc5859 (
      {stage0_63[423]},
      {stage1_63[206]}
   );
   gpc1_1 gpc5860 (
      {stage0_63[424]},
      {stage1_63[207]}
   );
   gpc1_1 gpc5861 (
      {stage0_63[425]},
      {stage1_63[208]}
   );
   gpc1_1 gpc5862 (
      {stage0_63[426]},
      {stage1_63[209]}
   );
   gpc1_1 gpc5863 (
      {stage0_63[427]},
      {stage1_63[210]}
   );
   gpc1_1 gpc5864 (
      {stage0_63[428]},
      {stage1_63[211]}
   );
   gpc1_1 gpc5865 (
      {stage0_63[429]},
      {stage1_63[212]}
   );
   gpc1_1 gpc5866 (
      {stage0_63[430]},
      {stage1_63[213]}
   );
   gpc1_1 gpc5867 (
      {stage0_63[431]},
      {stage1_63[214]}
   );
   gpc1_1 gpc5868 (
      {stage0_63[432]},
      {stage1_63[215]}
   );
   gpc1_1 gpc5869 (
      {stage0_63[433]},
      {stage1_63[216]}
   );
   gpc1_1 gpc5870 (
      {stage0_63[434]},
      {stage1_63[217]}
   );
   gpc1_1 gpc5871 (
      {stage0_63[435]},
      {stage1_63[218]}
   );
   gpc1_1 gpc5872 (
      {stage0_63[436]},
      {stage1_63[219]}
   );
   gpc1_1 gpc5873 (
      {stage0_63[437]},
      {stage1_63[220]}
   );
   gpc1_1 gpc5874 (
      {stage0_63[438]},
      {stage1_63[221]}
   );
   gpc1_1 gpc5875 (
      {stage0_63[439]},
      {stage1_63[222]}
   );
   gpc1_1 gpc5876 (
      {stage0_63[440]},
      {stage1_63[223]}
   );
   gpc1_1 gpc5877 (
      {stage0_63[441]},
      {stage1_63[224]}
   );
   gpc1_1 gpc5878 (
      {stage0_63[442]},
      {stage1_63[225]}
   );
   gpc1_1 gpc5879 (
      {stage0_63[443]},
      {stage1_63[226]}
   );
   gpc1_1 gpc5880 (
      {stage0_63[444]},
      {stage1_63[227]}
   );
   gpc1_1 gpc5881 (
      {stage0_63[445]},
      {stage1_63[228]}
   );
   gpc1_1 gpc5882 (
      {stage0_63[446]},
      {stage1_63[229]}
   );
   gpc1_1 gpc5883 (
      {stage0_63[447]},
      {stage1_63[230]}
   );
   gpc1_1 gpc5884 (
      {stage0_63[448]},
      {stage1_63[231]}
   );
   gpc1_1 gpc5885 (
      {stage0_63[449]},
      {stage1_63[232]}
   );
   gpc1_1 gpc5886 (
      {stage0_63[450]},
      {stage1_63[233]}
   );
   gpc1_1 gpc5887 (
      {stage0_63[451]},
      {stage1_63[234]}
   );
   gpc1_1 gpc5888 (
      {stage0_63[452]},
      {stage1_63[235]}
   );
   gpc1_1 gpc5889 (
      {stage0_63[453]},
      {stage1_63[236]}
   );
   gpc1_1 gpc5890 (
      {stage0_63[454]},
      {stage1_63[237]}
   );
   gpc1_1 gpc5891 (
      {stage0_63[455]},
      {stage1_63[238]}
   );
   gpc1_1 gpc5892 (
      {stage0_63[456]},
      {stage1_63[239]}
   );
   gpc1_1 gpc5893 (
      {stage0_63[457]},
      {stage1_63[240]}
   );
   gpc1_1 gpc5894 (
      {stage0_63[458]},
      {stage1_63[241]}
   );
   gpc1_1 gpc5895 (
      {stage0_63[459]},
      {stage1_63[242]}
   );
   gpc1_1 gpc5896 (
      {stage0_63[460]},
      {stage1_63[243]}
   );
   gpc1_1 gpc5897 (
      {stage0_63[461]},
      {stage1_63[244]}
   );
   gpc1_1 gpc5898 (
      {stage0_63[462]},
      {stage1_63[245]}
   );
   gpc1_1 gpc5899 (
      {stage0_63[463]},
      {stage1_63[246]}
   );
   gpc1_1 gpc5900 (
      {stage0_63[464]},
      {stage1_63[247]}
   );
   gpc1_1 gpc5901 (
      {stage0_63[465]},
      {stage1_63[248]}
   );
   gpc1_1 gpc5902 (
      {stage0_63[466]},
      {stage1_63[249]}
   );
   gpc1_1 gpc5903 (
      {stage0_63[467]},
      {stage1_63[250]}
   );
   gpc1_1 gpc5904 (
      {stage0_63[468]},
      {stage1_63[251]}
   );
   gpc1_1 gpc5905 (
      {stage0_63[469]},
      {stage1_63[252]}
   );
   gpc1_1 gpc5906 (
      {stage0_63[470]},
      {stage1_63[253]}
   );
   gpc1_1 gpc5907 (
      {stage0_63[471]},
      {stage1_63[254]}
   );
   gpc1_1 gpc5908 (
      {stage0_63[472]},
      {stage1_63[255]}
   );
   gpc1_1 gpc5909 (
      {stage0_63[473]},
      {stage1_63[256]}
   );
   gpc1_1 gpc5910 (
      {stage0_63[474]},
      {stage1_63[257]}
   );
   gpc1_1 gpc5911 (
      {stage0_63[475]},
      {stage1_63[258]}
   );
   gpc1_1 gpc5912 (
      {stage0_63[476]},
      {stage1_63[259]}
   );
   gpc1_1 gpc5913 (
      {stage0_63[477]},
      {stage1_63[260]}
   );
   gpc1_1 gpc5914 (
      {stage0_63[478]},
      {stage1_63[261]}
   );
   gpc1_1 gpc5915 (
      {stage0_63[479]},
      {stage1_63[262]}
   );
   gpc1_1 gpc5916 (
      {stage0_63[480]},
      {stage1_63[263]}
   );
   gpc1_1 gpc5917 (
      {stage0_63[481]},
      {stage1_63[264]}
   );
   gpc1_1 gpc5918 (
      {stage0_63[482]},
      {stage1_63[265]}
   );
   gpc1_1 gpc5919 (
      {stage0_63[483]},
      {stage1_63[266]}
   );
   gpc1_1 gpc5920 (
      {stage0_63[484]},
      {stage1_63[267]}
   );
   gpc1_1 gpc5921 (
      {stage0_63[485]},
      {stage1_63[268]}
   );
   gpc1_1 gpc5922 (
      {stage0_63[486]},
      {stage1_63[269]}
   );
   gpc1_1 gpc5923 (
      {stage0_63[487]},
      {stage1_63[270]}
   );
   gpc1_1 gpc5924 (
      {stage0_63[488]},
      {stage1_63[271]}
   );
   gpc1_1 gpc5925 (
      {stage0_63[489]},
      {stage1_63[272]}
   );
   gpc1_1 gpc5926 (
      {stage0_63[490]},
      {stage1_63[273]}
   );
   gpc1_1 gpc5927 (
      {stage0_63[491]},
      {stage1_63[274]}
   );
   gpc1_1 gpc5928 (
      {stage0_63[492]},
      {stage1_63[275]}
   );
   gpc1_1 gpc5929 (
      {stage0_63[493]},
      {stage1_63[276]}
   );
   gpc1_1 gpc5930 (
      {stage0_63[494]},
      {stage1_63[277]}
   );
   gpc1_1 gpc5931 (
      {stage0_63[495]},
      {stage1_63[278]}
   );
   gpc1_1 gpc5932 (
      {stage0_63[496]},
      {stage1_63[279]}
   );
   gpc1_1 gpc5933 (
      {stage0_63[497]},
      {stage1_63[280]}
   );
   gpc1_1 gpc5934 (
      {stage0_63[498]},
      {stage1_63[281]}
   );
   gpc1_1 gpc5935 (
      {stage0_63[499]},
      {stage1_63[282]}
   );
   gpc1_1 gpc5936 (
      {stage0_63[500]},
      {stage1_63[283]}
   );
   gpc1_1 gpc5937 (
      {stage0_63[501]},
      {stage1_63[284]}
   );
   gpc1_1 gpc5938 (
      {stage0_63[502]},
      {stage1_63[285]}
   );
   gpc1_1 gpc5939 (
      {stage0_63[503]},
      {stage1_63[286]}
   );
   gpc1_1 gpc5940 (
      {stage0_63[504]},
      {stage1_63[287]}
   );
   gpc1_1 gpc5941 (
      {stage0_63[505]},
      {stage1_63[288]}
   );
   gpc1_1 gpc5942 (
      {stage0_63[506]},
      {stage1_63[289]}
   );
   gpc1_1 gpc5943 (
      {stage0_63[507]},
      {stage1_63[290]}
   );
   gpc1_1 gpc5944 (
      {stage0_63[508]},
      {stage1_63[291]}
   );
   gpc1_1 gpc5945 (
      {stage0_63[509]},
      {stage1_63[292]}
   );
   gpc1_1 gpc5946 (
      {stage0_63[510]},
      {stage1_63[293]}
   );
   gpc1_1 gpc5947 (
      {stage0_63[511]},
      {stage1_63[294]}
   );
   gpc1163_5 gpc5948 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc5949 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc5950 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc5951 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc5952 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc5953 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc5954 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc5955 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc5956 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc5957 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc5958 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc5959 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc5960 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc5961 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc5962 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc5963 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc5964 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc5965 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc5966 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc5967 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc5968 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc5969 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc5970 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc5971 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc5972 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc615_5 gpc5973 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106]},
      {stage1_1[96]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc615_5 gpc5974 (
      {stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111]},
      {stage1_1[97]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc5975 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[0],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc5976 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[1],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc5977 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[2],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc5978 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[3],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc5979 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[4],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc5980 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[5],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc5981 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[6],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc5982 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage2_5[7],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc5983 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69]},
      {stage2_5[8],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc5984 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage2_5[9],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc5985 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage2_5[10],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc5986 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], 1'b0},
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87]},
      {stage2_5[11],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc5987 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[12],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc5988 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[13],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc5989 (
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[14],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc5990 (
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[15],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc5991 (
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[16],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc606_5 gpc5992 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[17],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc606_5 gpc5993 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[18],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc606_5 gpc5994 (
      {stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[19],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc5995 (
      {stage1_2[130], stage1_2[131], stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[20],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc5996 (
      {stage1_2[136], stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[21],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc606_5 gpc5997 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[22],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc606_5 gpc5998 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152], stage1_2[153]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[23],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc606_5 gpc5999 (
      {stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157], stage1_2[158], stage1_2[159]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[24],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc606_5 gpc6000 (
      {stage1_2[160], stage1_2[161], stage1_2[162], stage1_2[163], stage1_2[164], stage1_2[165]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[25],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc606_5 gpc6001 (
      {stage1_2[166], stage1_2[167], stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[26],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc606_5 gpc6002 (
      {stage1_2[172], stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[27],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc606_5 gpc6003 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182], stage1_2[183]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[28],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc606_5 gpc6004 (
      {stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187], stage1_2[188], stage1_2[189]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[29],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc606_5 gpc6005 (
      {stage1_2[190], stage1_2[191], stage1_2[192], stage1_2[193], stage1_2[194], stage1_2[195]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[30],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc606_5 gpc6006 (
      {stage1_2[196], stage1_2[197], stage1_2[198], stage1_2[199], stage1_2[200], stage1_2[201]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[31],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc606_5 gpc6007 (
      {stage1_2[202], stage1_2[203], stage1_2[204], stage1_2[205], stage1_2[206], stage1_2[207]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[32],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc1415_5 gpc6008 (
      {stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92]},
      {stage1_4[126]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[21],stage2_5[33],stage2_4[60],stage2_3[60]}
   );
   gpc1415_5 gpc6009 (
      {stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage1_4[127]},
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7]},
      {stage1_6[1]},
      {stage2_7[1],stage2_6[22],stage2_5[34],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc6010 (
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102]},
      {stage1_4[128]},
      {stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13]},
      {stage2_7[2],stage2_6[23],stage2_5[35],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc6011 (
      {stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage1_4[129]},
      {stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19]},
      {stage2_7[3],stage2_6[24],stage2_5[36],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc6012 (
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112]},
      {stage1_4[130]},
      {stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25]},
      {stage2_7[4],stage2_6[25],stage2_5[37],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc6013 (
      {stage1_3[113], stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117]},
      {stage1_4[131]},
      {stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31]},
      {stage2_7[5],stage2_6[26],stage2_5[38],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc6014 (
      {stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122]},
      {stage1_4[132]},
      {stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37]},
      {stage2_7[6],stage2_6[27],stage2_5[39],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc6015 (
      {stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage1_4[133]},
      {stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43]},
      {stage2_7[7],stage2_6[28],stage2_5[40],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc6016 (
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132]},
      {stage1_4[134]},
      {stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49]},
      {stage2_7[8],stage2_6[29],stage2_5[41],stage2_4[68],stage2_3[68]}
   );
   gpc623_5 gpc6017 (
      {stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[135], stage1_4[136]},
      {stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55]},
      {stage2_7[9],stage2_6[30],stage2_5[42],stage2_4[69],stage2_3[69]}
   );
   gpc623_5 gpc6018 (
      {stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[137], stage1_4[138]},
      {stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61]},
      {stage2_7[10],stage2_6[31],stage2_5[43],stage2_4[70],stage2_3[70]}
   );
   gpc606_5 gpc6019 (
      {stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[11],stage2_6[32],stage2_5[44],stage2_4[71]}
   );
   gpc606_5 gpc6020 (
      {stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[12],stage2_6[33],stage2_5[45],stage2_4[72]}
   );
   gpc606_5 gpc6021 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[13],stage2_6[34],stage2_5[46],stage2_4[73]}
   );
   gpc606_5 gpc6022 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162]},
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage2_8[3],stage2_7[14],stage2_6[35],stage2_5[47],stage2_4[74]}
   );
   gpc606_5 gpc6023 (
      {stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168]},
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage2_8[4],stage2_7[15],stage2_6[36],stage2_5[48],stage2_4[75]}
   );
   gpc606_5 gpc6024 (
      {stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174]},
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36], stage1_6[37]},
      {stage2_8[5],stage2_7[16],stage2_6[37],stage2_5[49],stage2_4[76]}
   );
   gpc606_5 gpc6025 (
      {stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42], stage1_6[43]},
      {stage2_8[6],stage2_7[17],stage2_6[38],stage2_5[50],stage2_4[77]}
   );
   gpc606_5 gpc6026 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49]},
      {stage2_8[7],stage2_7[18],stage2_6[39],stage2_5[51],stage2_4[78]}
   );
   gpc606_5 gpc6027 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192]},
      {stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage2_8[8],stage2_7[19],stage2_6[40],stage2_5[52],stage2_4[79]}
   );
   gpc606_5 gpc6028 (
      {stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198]},
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage2_8[9],stage2_7[20],stage2_6[41],stage2_5[53],stage2_4[80]}
   );
   gpc606_5 gpc6029 (
      {stage1_4[199], stage1_4[200], stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204]},
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66], stage1_6[67]},
      {stage2_8[10],stage2_7[21],stage2_6[42],stage2_5[54],stage2_4[81]}
   );
   gpc606_5 gpc6030 (
      {stage1_4[205], stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72], stage1_6[73]},
      {stage2_8[11],stage2_7[22],stage2_6[43],stage2_5[55],stage2_4[82]}
   );
   gpc606_5 gpc6031 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79]},
      {stage2_8[12],stage2_7[23],stage2_6[44],stage2_5[56],stage2_4[83]}
   );
   gpc606_5 gpc6032 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221], stage1_4[222]},
      {stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage2_8[13],stage2_7[24],stage2_6[45],stage2_5[57],stage2_4[84]}
   );
   gpc606_5 gpc6033 (
      {stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227], stage1_4[228]},
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage2_8[14],stage2_7[25],stage2_6[46],stage2_5[58],stage2_4[85]}
   );
   gpc606_5 gpc6034 (
      {stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233], stage1_4[234]},
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96], stage1_6[97]},
      {stage2_8[15],stage2_7[26],stage2_6[47],stage2_5[59],stage2_4[86]}
   );
   gpc606_5 gpc6035 (
      {stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239], stage1_4[240]},
      {stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102], stage1_6[103]},
      {stage2_8[16],stage2_7[27],stage2_6[48],stage2_5[60],stage2_4[87]}
   );
   gpc606_5 gpc6036 (
      {stage1_4[241], stage1_4[242], stage1_4[243], stage1_4[244], stage1_4[245], stage1_4[246]},
      {stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108], stage1_6[109]},
      {stage2_8[17],stage2_7[28],stage2_6[49],stage2_5[61],stage2_4[88]}
   );
   gpc606_5 gpc6037 (
      {stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[18],stage2_7[29],stage2_6[50],stage2_5[62]}
   );
   gpc606_5 gpc6038 (
      {stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[19],stage2_7[30],stage2_6[51],stage2_5[63]}
   );
   gpc606_5 gpc6039 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[20],stage2_7[31],stage2_6[52],stage2_5[64]}
   );
   gpc606_5 gpc6040 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[21],stage2_7[32],stage2_6[53],stage2_5[65]}
   );
   gpc606_5 gpc6041 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[22],stage2_7[33],stage2_6[54],stage2_5[66]}
   );
   gpc606_5 gpc6042 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[23],stage2_7[34],stage2_6[55],stage2_5[67]}
   );
   gpc606_5 gpc6043 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[24],stage2_7[35],stage2_6[56],stage2_5[68]}
   );
   gpc606_5 gpc6044 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[25],stage2_7[36],stage2_6[57],stage2_5[69]}
   );
   gpc606_5 gpc6045 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[26],stage2_7[37],stage2_6[58],stage2_5[70]}
   );
   gpc606_5 gpc6046 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[27],stage2_7[38],stage2_6[59],stage2_5[71]}
   );
   gpc606_5 gpc6047 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[28],stage2_7[39],stage2_6[60],stage2_5[72]}
   );
   gpc606_5 gpc6048 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[29],stage2_7[40],stage2_6[61],stage2_5[73]}
   );
   gpc606_5 gpc6049 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[30],stage2_7[41],stage2_6[62],stage2_5[74]}
   );
   gpc606_5 gpc6050 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[31],stage2_7[42],stage2_6[63],stage2_5[75]}
   );
   gpc606_5 gpc6051 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[32],stage2_7[43],stage2_6[64],stage2_5[76]}
   );
   gpc606_5 gpc6052 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[33],stage2_7[44],stage2_6[65],stage2_5[77]}
   );
   gpc606_5 gpc6053 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[34],stage2_7[45],stage2_6[66],stage2_5[78]}
   );
   gpc606_5 gpc6054 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[35],stage2_7[46],stage2_6[67],stage2_5[79]}
   );
   gpc606_5 gpc6055 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[36],stage2_7[47],stage2_6[68],stage2_5[80]}
   );
   gpc606_5 gpc6056 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[114], stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage2_9[19],stage2_8[37],stage2_7[48],stage2_6[69],stage2_5[81]}
   );
   gpc606_5 gpc6057 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage2_9[20],stage2_8[38],stage2_7[49],stage2_6[70],stage2_5[82]}
   );
   gpc615_5 gpc6058 (
      {stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_7[126]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[21],stage2_8[39],stage2_7[50],stage2_6[71]}
   );
   gpc615_5 gpc6059 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_7[127]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[22],stage2_8[40],stage2_7[51],stage2_6[72]}
   );
   gpc615_5 gpc6060 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124]},
      {stage1_7[128]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[23],stage2_8[41],stage2_7[52],stage2_6[73]}
   );
   gpc615_5 gpc6061 (
      {stage1_6[125], stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129]},
      {stage1_7[129]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[24],stage2_8[42],stage2_7[53],stage2_6[74]}
   );
   gpc615_5 gpc6062 (
      {stage1_6[130], stage1_6[131], stage1_6[132], stage1_6[133], stage1_6[134]},
      {stage1_7[130]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[25],stage2_8[43],stage2_7[54],stage2_6[75]}
   );
   gpc615_5 gpc6063 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[26],stage2_8[44],stage2_7[55]}
   );
   gpc615_5 gpc6064 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[27],stage2_8[45],stage2_7[56]}
   );
   gpc615_5 gpc6065 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[28],stage2_8[46],stage2_7[57]}
   );
   gpc615_5 gpc6066 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[29],stage2_8[47],stage2_7[58]}
   );
   gpc615_5 gpc6067 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[30],stage2_8[48],stage2_7[59]}
   );
   gpc615_5 gpc6068 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[31],stage2_8[49],stage2_7[60]}
   );
   gpc615_5 gpc6069 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[36]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[32],stage2_8[50],stage2_7[61]}
   );
   gpc615_5 gpc6070 (
      {stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170]},
      {stage1_8[37]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[33],stage2_8[51],stage2_7[62]}
   );
   gpc615_5 gpc6071 (
      {stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175]},
      {stage1_8[38]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[34],stage2_8[52],stage2_7[63]}
   );
   gpc615_5 gpc6072 (
      {stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_8[39]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[35],stage2_8[53],stage2_7[64]}
   );
   gpc615_5 gpc6073 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185]},
      {stage1_8[40]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[36],stage2_8[54],stage2_7[65]}
   );
   gpc615_5 gpc6074 (
      {stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190]},
      {stage1_8[41]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[37],stage2_8[55],stage2_7[66]}
   );
   gpc615_5 gpc6075 (
      {stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195]},
      {stage1_8[42]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[38],stage2_8[56],stage2_7[67]}
   );
   gpc615_5 gpc6076 (
      {stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200]},
      {stage1_8[43]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[39],stage2_8[57],stage2_7[68]}
   );
   gpc615_5 gpc6077 (
      {stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205]},
      {stage1_8[44]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[40],stage2_8[58],stage2_7[69]}
   );
   gpc615_5 gpc6078 (
      {stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_8[45]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[41],stage2_8[59],stage2_7[70]}
   );
   gpc615_5 gpc6079 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215]},
      {stage1_8[46]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[42],stage2_8[60],stage2_7[71]}
   );
   gpc615_5 gpc6080 (
      {stage1_7[216], stage1_7[217], stage1_7[218], stage1_7[219], stage1_7[220]},
      {stage1_8[47]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[43],stage2_8[61],stage2_7[72]}
   );
   gpc615_5 gpc6081 (
      {stage1_7[221], stage1_7[222], stage1_7[223], stage1_7[224], stage1_7[225]},
      {stage1_8[48]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[44],stage2_8[62],stage2_7[73]}
   );
   gpc615_5 gpc6082 (
      {stage1_7[226], stage1_7[227], stage1_7[228], stage1_7[229], stage1_7[230]},
      {stage1_8[49]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[45],stage2_8[63],stage2_7[74]}
   );
   gpc615_5 gpc6083 (
      {stage1_7[231], stage1_7[232], stage1_7[233], stage1_7[234], stage1_7[235]},
      {stage1_8[50]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[46],stage2_8[64],stage2_7[75]}
   );
   gpc615_5 gpc6084 (
      {stage1_7[236], stage1_7[237], stage1_7[238], stage1_7[239], stage1_7[240]},
      {stage1_8[51]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[26],stage2_9[47],stage2_8[65],stage2_7[76]}
   );
   gpc615_5 gpc6085 (
      {stage1_7[241], stage1_7[242], stage1_7[243], stage1_7[244], stage1_7[245]},
      {stage1_8[52]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[27],stage2_9[48],stage2_8[66],stage2_7[77]}
   );
   gpc615_5 gpc6086 (
      {stage1_7[246], stage1_7[247], stage1_7[248], stage1_7[249], stage1_7[250]},
      {stage1_8[53]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[28],stage2_9[49],stage2_8[67],stage2_7[78]}
   );
   gpc615_5 gpc6087 (
      {stage1_7[251], stage1_7[252], stage1_7[253], stage1_7[254], stage1_7[255]},
      {stage1_8[54]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[29],stage2_9[50],stage2_8[68],stage2_7[79]}
   );
   gpc615_5 gpc6088 (
      {stage1_7[256], stage1_7[257], stage1_7[258], stage1_7[259], stage1_7[260]},
      {stage1_8[55]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[30],stage2_9[51],stage2_8[69],stage2_7[80]}
   );
   gpc615_5 gpc6089 (
      {stage1_7[261], stage1_7[262], stage1_7[263], stage1_7[264], stage1_7[265]},
      {stage1_8[56]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[31],stage2_9[52],stage2_8[70],stage2_7[81]}
   );
   gpc615_5 gpc6090 (
      {stage1_7[266], stage1_7[267], stage1_7[268], stage1_7[269], stage1_7[270]},
      {stage1_8[57]},
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage2_11[27],stage2_10[32],stage2_9[53],stage2_8[71],stage2_7[82]}
   );
   gpc615_5 gpc6091 (
      {stage1_7[271], stage1_7[272], stage1_7[273], stage1_7[274], stage1_7[275]},
      {stage1_8[58]},
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage2_11[28],stage2_10[33],stage2_9[54],stage2_8[72],stage2_7[83]}
   );
   gpc615_5 gpc6092 (
      {stage1_7[276], stage1_7[277], stage1_7[278], stage1_7[279], stage1_7[280]},
      {stage1_8[59]},
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage2_11[29],stage2_10[34],stage2_9[55],stage2_8[73],stage2_7[84]}
   );
   gpc615_5 gpc6093 (
      {stage1_7[281], stage1_7[282], stage1_7[283], stage1_7[284], stage1_7[285]},
      {stage1_8[60]},
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage2_11[30],stage2_10[35],stage2_9[56],stage2_8[74],stage2_7[85]}
   );
   gpc615_5 gpc6094 (
      {stage1_7[286], stage1_7[287], stage1_7[288], stage1_7[289], stage1_7[290]},
      {stage1_8[61]},
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage2_11[31],stage2_10[36],stage2_9[57],stage2_8[75],stage2_7[86]}
   );
   gpc615_5 gpc6095 (
      {stage1_7[291], stage1_7[292], stage1_7[293], stage1_7[294], stage1_7[295]},
      {stage1_8[62]},
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage2_11[32],stage2_10[37],stage2_9[58],stage2_8[76],stage2_7[87]}
   );
   gpc615_5 gpc6096 (
      {stage1_7[296], stage1_7[297], stage1_7[298], stage1_7[299], stage1_7[300]},
      {stage1_8[63]},
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage2_11[33],stage2_10[38],stage2_9[59],stage2_8[77],stage2_7[88]}
   );
   gpc615_5 gpc6097 (
      {stage1_7[301], stage1_7[302], stage1_7[303], stage1_7[304], stage1_7[305]},
      {stage1_8[64]},
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage2_11[34],stage2_10[39],stage2_9[60],stage2_8[78],stage2_7[89]}
   );
   gpc615_5 gpc6098 (
      {stage1_7[306], stage1_7[307], stage1_7[308], stage1_7[309], stage1_7[310]},
      {stage1_8[65]},
      {stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213], stage1_9[214], stage1_9[215]},
      {stage2_11[35],stage2_10[40],stage2_9[61],stage2_8[79],stage2_7[90]}
   );
   gpc615_5 gpc6099 (
      {stage1_7[311], stage1_7[312], stage1_7[313], stage1_7[314], stage1_7[315]},
      {stage1_8[66]},
      {stage1_9[216], stage1_9[217], stage1_9[218], stage1_9[219], stage1_9[220], stage1_9[221]},
      {stage2_11[36],stage2_10[41],stage2_9[62],stage2_8[80],stage2_7[91]}
   );
   gpc615_5 gpc6100 (
      {stage1_7[316], stage1_7[317], stage1_7[318], stage1_7[319], stage1_7[320]},
      {stage1_8[67]},
      {stage1_9[222], stage1_9[223], stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227]},
      {stage2_11[37],stage2_10[42],stage2_9[63],stage2_8[81],stage2_7[92]}
   );
   gpc615_5 gpc6101 (
      {stage1_7[321], stage1_7[322], stage1_7[323], stage1_7[324], stage1_7[325]},
      {stage1_8[68]},
      {stage1_9[228], stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage2_11[38],stage2_10[43],stage2_9[64],stage2_8[82],stage2_7[93]}
   );
   gpc615_5 gpc6102 (
      {stage1_7[326], stage1_7[327], stage1_7[328], stage1_7[329], stage1_7[330]},
      {stage1_8[69]},
      {stage1_9[234], stage1_9[235], stage1_9[236], stage1_9[237], stage1_9[238], stage1_9[239]},
      {stage2_11[39],stage2_10[44],stage2_9[65],stage2_8[83],stage2_7[94]}
   );
   gpc615_5 gpc6103 (
      {stage1_7[331], stage1_7[332], stage1_7[333], stage1_7[334], stage1_7[335]},
      {stage1_8[70]},
      {stage1_9[240], stage1_9[241], stage1_9[242], stage1_9[243], stage1_9[244], stage1_9[245]},
      {stage2_11[40],stage2_10[45],stage2_9[66],stage2_8[84],stage2_7[95]}
   );
   gpc615_5 gpc6104 (
      {stage1_7[336], stage1_7[337], stage1_7[338], stage1_7[339], 1'b0},
      {stage1_8[71]},
      {stage1_9[246], stage1_9[247], stage1_9[248], stage1_9[249], stage1_9[250], stage1_9[251]},
      {stage2_11[41],stage2_10[46],stage2_9[67],stage2_8[85],stage2_7[96]}
   );
   gpc606_5 gpc6105 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[42],stage2_10[47],stage2_9[68],stage2_8[86]}
   );
   gpc606_5 gpc6106 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[43],stage2_10[48],stage2_9[69],stage2_8[87]}
   );
   gpc606_5 gpc6107 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[44],stage2_10[49],stage2_9[70],stage2_8[88]}
   );
   gpc606_5 gpc6108 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[45],stage2_10[50],stage2_9[71],stage2_8[89]}
   );
   gpc606_5 gpc6109 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[46],stage2_10[51],stage2_9[72],stage2_8[90]}
   );
   gpc606_5 gpc6110 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[47],stage2_10[52],stage2_9[73],stage2_8[91]}
   );
   gpc606_5 gpc6111 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[48],stage2_10[53],stage2_9[74],stage2_8[92]}
   );
   gpc606_5 gpc6112 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[49],stage2_10[54],stage2_9[75],stage2_8[93]}
   );
   gpc606_5 gpc6113 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[50],stage2_10[55],stage2_9[76],stage2_8[94]}
   );
   gpc606_5 gpc6114 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[51],stage2_10[56],stage2_9[77],stage2_8[95]}
   );
   gpc606_5 gpc6115 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[52],stage2_10[57],stage2_9[78],stage2_8[96]}
   );
   gpc606_5 gpc6116 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[53],stage2_10[58],stage2_9[79],stage2_8[97]}
   );
   gpc606_5 gpc6117 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[54],stage2_10[59],stage2_9[80],stage2_8[98]}
   );
   gpc606_5 gpc6118 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[55],stage2_10[60],stage2_9[81],stage2_8[99]}
   );
   gpc606_5 gpc6119 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[56],stage2_10[61],stage2_9[82],stage2_8[100]}
   );
   gpc606_5 gpc6120 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[57],stage2_10[62],stage2_9[83],stage2_8[101]}
   );
   gpc606_5 gpc6121 (
      {stage1_9[252], stage1_9[253], stage1_9[254], stage1_9[255], stage1_9[256], stage1_9[257]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[16],stage2_11[58],stage2_10[63],stage2_9[84]}
   );
   gpc606_5 gpc6122 (
      {stage1_9[258], stage1_9[259], stage1_9[260], stage1_9[261], stage1_9[262], stage1_9[263]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[17],stage2_11[59],stage2_10[64],stage2_9[85]}
   );
   gpc606_5 gpc6123 (
      {stage1_9[264], stage1_9[265], stage1_9[266], stage1_9[267], stage1_9[268], stage1_9[269]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[18],stage2_11[60],stage2_10[65],stage2_9[86]}
   );
   gpc606_5 gpc6124 (
      {stage1_9[270], stage1_9[271], stage1_9[272], stage1_9[273], stage1_9[274], stage1_9[275]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[19],stage2_11[61],stage2_10[66],stage2_9[87]}
   );
   gpc606_5 gpc6125 (
      {stage1_9[276], stage1_9[277], stage1_9[278], stage1_9[279], stage1_9[280], stage1_9[281]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[20],stage2_11[62],stage2_10[67],stage2_9[88]}
   );
   gpc606_5 gpc6126 (
      {stage1_9[282], stage1_9[283], stage1_9[284], stage1_9[285], stage1_9[286], stage1_9[287]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[21],stage2_11[63],stage2_10[68],stage2_9[89]}
   );
   gpc606_5 gpc6127 (
      {stage1_9[288], stage1_9[289], stage1_9[290], stage1_9[291], stage1_9[292], stage1_9[293]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[22],stage2_11[64],stage2_10[69],stage2_9[90]}
   );
   gpc606_5 gpc6128 (
      {stage1_9[294], stage1_9[295], stage1_9[296], stage1_9[297], stage1_9[298], stage1_9[299]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[23],stage2_11[65],stage2_10[70],stage2_9[91]}
   );
   gpc606_5 gpc6129 (
      {stage1_9[300], stage1_9[301], stage1_9[302], stage1_9[303], stage1_9[304], stage1_9[305]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[24],stage2_11[66],stage2_10[71],stage2_9[92]}
   );
   gpc606_5 gpc6130 (
      {stage1_9[306], stage1_9[307], stage1_9[308], stage1_9[309], stage1_9[310], stage1_9[311]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[25],stage2_11[67],stage2_10[72],stage2_9[93]}
   );
   gpc606_5 gpc6131 (
      {stage1_9[312], stage1_9[313], stage1_9[314], stage1_9[315], stage1_9[316], stage1_9[317]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[26],stage2_11[68],stage2_10[73],stage2_9[94]}
   );
   gpc606_5 gpc6132 (
      {stage1_9[318], stage1_9[319], stage1_9[320], stage1_9[321], stage1_9[322], stage1_9[323]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[27],stage2_11[69],stage2_10[74],stage2_9[95]}
   );
   gpc606_5 gpc6133 (
      {stage1_9[324], stage1_9[325], stage1_9[326], stage1_9[327], stage1_9[328], stage1_9[329]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[28],stage2_11[70],stage2_10[75],stage2_9[96]}
   );
   gpc606_5 gpc6134 (
      {stage1_9[330], stage1_9[331], stage1_9[332], stage1_9[333], stage1_9[334], stage1_9[335]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[29],stage2_11[71],stage2_10[76],stage2_9[97]}
   );
   gpc606_5 gpc6135 (
      {stage1_9[336], stage1_9[337], stage1_9[338], stage1_9[339], stage1_9[340], stage1_9[341]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[30],stage2_11[72],stage2_10[77],stage2_9[98]}
   );
   gpc606_5 gpc6136 (
      {stage1_9[342], stage1_9[343], stage1_9[344], stage1_9[345], stage1_9[346], stage1_9[347]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[31],stage2_11[73],stage2_10[78],stage2_9[99]}
   );
   gpc606_5 gpc6137 (
      {stage1_9[348], stage1_9[349], stage1_9[350], stage1_9[351], stage1_9[352], stage1_9[353]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[32],stage2_11[74],stage2_10[79],stage2_9[100]}
   );
   gpc606_5 gpc6138 (
      {stage1_9[354], stage1_9[355], stage1_9[356], stage1_9[357], stage1_9[358], stage1_9[359]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[33],stage2_11[75],stage2_10[80],stage2_9[101]}
   );
   gpc615_5 gpc6139 (
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_11[108]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[34],stage2_11[76],stage2_10[81]}
   );
   gpc1163_5 gpc6140 (
      {stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_13[0]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[19],stage2_12[35],stage2_11[77]}
   );
   gpc1163_5 gpc6141 (
      {stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage1_13[1]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[20],stage2_12[36],stage2_11[78]}
   );
   gpc1163_5 gpc6142 (
      {stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage1_13[2]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[21],stage2_12[37],stage2_11[79]}
   );
   gpc1163_5 gpc6143 (
      {stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage1_13[3]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[22],stage2_12[38],stage2_11[80]}
   );
   gpc1163_5 gpc6144 (
      {stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage1_13[4]},
      {stage1_14[4]},
      {stage2_15[4],stage2_14[5],stage2_13[23],stage2_12[39],stage2_11[81]}
   );
   gpc1163_5 gpc6145 (
      {stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[5]},
      {stage1_14[5]},
      {stage2_15[5],stage2_14[6],stage2_13[24],stage2_12[40],stage2_11[82]}
   );
   gpc1163_5 gpc6146 (
      {stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_13[6]},
      {stage1_14[6]},
      {stage2_15[6],stage2_14[7],stage2_13[25],stage2_12[41],stage2_11[83]}
   );
   gpc1163_5 gpc6147 (
      {stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_13[7]},
      {stage1_14[7]},
      {stage2_15[7],stage2_14[8],stage2_13[26],stage2_12[42],stage2_11[84]}
   );
   gpc1163_5 gpc6148 (
      {stage1_11[133], stage1_11[134], stage1_11[135]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[8]},
      {stage1_14[8]},
      {stage2_15[8],stage2_14[9],stage2_13[27],stage2_12[43],stage2_11[85]}
   );
   gpc1163_5 gpc6149 (
      {stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_13[9]},
      {stage1_14[9]},
      {stage2_15[9],stage2_14[10],stage2_13[28],stage2_12[44],stage2_11[86]}
   );
   gpc1163_5 gpc6150 (
      {stage1_11[139], stage1_11[140], stage1_11[141]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage1_13[10]},
      {stage1_14[10]},
      {stage2_15[10],stage2_14[11],stage2_13[29],stage2_12[45],stage2_11[87]}
   );
   gpc1163_5 gpc6151 (
      {stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage1_13[11]},
      {stage1_14[11]},
      {stage2_15[11],stage2_14[12],stage2_13[30],stage2_12[46],stage2_11[88]}
   );
   gpc1163_5 gpc6152 (
      {stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage1_13[12]},
      {stage1_14[12]},
      {stage2_15[12],stage2_14[13],stage2_13[31],stage2_12[47],stage2_11[89]}
   );
   gpc1163_5 gpc6153 (
      {stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[13]},
      {stage1_14[13]},
      {stage2_15[13],stage2_14[14],stage2_13[32],stage2_12[48],stage2_11[90]}
   );
   gpc1163_5 gpc6154 (
      {stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage1_13[14]},
      {stage1_14[14]},
      {stage2_15[14],stage2_14[15],stage2_13[33],stage2_12[49],stage2_11[91]}
   );
   gpc1163_5 gpc6155 (
      {stage1_11[154], stage1_11[155], stage1_11[156]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_13[15]},
      {stage1_14[15]},
      {stage2_15[15],stage2_14[16],stage2_13[34],stage2_12[50],stage2_11[92]}
   );
   gpc1163_5 gpc6156 (
      {stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage1_13[16]},
      {stage1_14[16]},
      {stage2_15[16],stage2_14[17],stage2_13[35],stage2_12[51],stage2_11[93]}
   );
   gpc1163_5 gpc6157 (
      {stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_13[17]},
      {stage1_14[17]},
      {stage2_15[17],stage2_14[18],stage2_13[36],stage2_12[52],stage2_11[94]}
   );
   gpc1163_5 gpc6158 (
      {stage1_11[163], stage1_11[164], stage1_11[165]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[18]},
      {stage1_14[18]},
      {stage2_15[18],stage2_14[19],stage2_13[37],stage2_12[53],stage2_11[95]}
   );
   gpc1163_5 gpc6159 (
      {stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_13[19]},
      {stage1_14[19]},
      {stage2_15[19],stage2_14[20],stage2_13[38],stage2_12[54],stage2_11[96]}
   );
   gpc1163_5 gpc6160 (
      {stage1_11[169], stage1_11[170], stage1_11[171]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_13[20]},
      {stage1_14[20]},
      {stage2_15[20],stage2_14[21],stage2_13[39],stage2_12[55],stage2_11[97]}
   );
   gpc615_5 gpc6161 (
      {stage1_11[172], stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176]},
      {stage1_12[132]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[21],stage2_14[22],stage2_13[40],stage2_12[56],stage2_11[98]}
   );
   gpc615_5 gpc6162 (
      {stage1_11[177], stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181]},
      {stage1_12[133]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[22],stage2_14[23],stage2_13[41],stage2_12[57],stage2_11[99]}
   );
   gpc615_5 gpc6163 (
      {stage1_11[182], stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186]},
      {stage1_12[134]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[23],stage2_14[24],stage2_13[42],stage2_12[58],stage2_11[100]}
   );
   gpc615_5 gpc6164 (
      {stage1_11[187], stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191]},
      {stage1_12[135]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[24],stage2_14[25],stage2_13[43],stage2_12[59],stage2_11[101]}
   );
   gpc615_5 gpc6165 (
      {stage1_11[192], stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196]},
      {stage1_12[136]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[25],stage2_14[26],stage2_13[44],stage2_12[60],stage2_11[102]}
   );
   gpc615_5 gpc6166 (
      {stage1_11[197], stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201]},
      {stage1_12[137]},
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage2_15[26],stage2_14[27],stage2_13[45],stage2_12[61],stage2_11[103]}
   );
   gpc615_5 gpc6167 (
      {stage1_11[202], stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206]},
      {stage1_12[138]},
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage2_15[27],stage2_14[28],stage2_13[46],stage2_12[62],stage2_11[104]}
   );
   gpc615_5 gpc6168 (
      {stage1_11[207], stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211]},
      {stage1_12[139]},
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage2_15[28],stage2_14[29],stage2_13[47],stage2_12[63],stage2_11[105]}
   );
   gpc615_5 gpc6169 (
      {stage1_11[212], stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216]},
      {stage1_12[140]},
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage2_15[29],stage2_14[30],stage2_13[48],stage2_12[64],stage2_11[106]}
   );
   gpc615_5 gpc6170 (
      {stage1_11[217], stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221]},
      {stage1_12[141]},
      {stage1_13[75], stage1_13[76], stage1_13[77], stage1_13[78], stage1_13[79], stage1_13[80]},
      {stage2_15[30],stage2_14[31],stage2_13[49],stage2_12[65],stage2_11[107]}
   );
   gpc615_5 gpc6171 (
      {stage1_11[222], stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226]},
      {stage1_12[142]},
      {stage1_13[81], stage1_13[82], stage1_13[83], stage1_13[84], stage1_13[85], stage1_13[86]},
      {stage2_15[31],stage2_14[32],stage2_13[50],stage2_12[66],stage2_11[108]}
   );
   gpc615_5 gpc6172 (
      {stage1_11[227], stage1_11[228], stage1_11[229], stage1_11[230], stage1_11[231]},
      {stage1_12[143]},
      {stage1_13[87], stage1_13[88], stage1_13[89], stage1_13[90], stage1_13[91], stage1_13[92]},
      {stage2_15[32],stage2_14[33],stage2_13[51],stage2_12[67],stage2_11[109]}
   );
   gpc615_5 gpc6173 (
      {stage1_11[232], stage1_11[233], stage1_11[234], stage1_11[235], stage1_11[236]},
      {stage1_12[144]},
      {stage1_13[93], stage1_13[94], stage1_13[95], stage1_13[96], stage1_13[97], stage1_13[98]},
      {stage2_15[33],stage2_14[34],stage2_13[52],stage2_12[68],stage2_11[110]}
   );
   gpc615_5 gpc6174 (
      {stage1_11[237], stage1_11[238], stage1_11[239], stage1_11[240], stage1_11[241]},
      {stage1_12[145]},
      {stage1_13[99], stage1_13[100], stage1_13[101], stage1_13[102], stage1_13[103], stage1_13[104]},
      {stage2_15[34],stage2_14[35],stage2_13[53],stage2_12[69],stage2_11[111]}
   );
   gpc615_5 gpc6175 (
      {stage1_11[242], stage1_11[243], stage1_11[244], stage1_11[245], stage1_11[246]},
      {stage1_12[146]},
      {stage1_13[105], stage1_13[106], stage1_13[107], stage1_13[108], stage1_13[109], stage1_13[110]},
      {stage2_15[35],stage2_14[36],stage2_13[54],stage2_12[70],stage2_11[112]}
   );
   gpc615_5 gpc6176 (
      {stage1_11[247], stage1_11[248], stage1_11[249], stage1_11[250], stage1_11[251]},
      {stage1_12[147]},
      {stage1_13[111], stage1_13[112], stage1_13[113], stage1_13[114], stage1_13[115], stage1_13[116]},
      {stage2_15[36],stage2_14[37],stage2_13[55],stage2_12[71],stage2_11[113]}
   );
   gpc615_5 gpc6177 (
      {stage1_11[252], stage1_11[253], stage1_11[254], stage1_11[255], stage1_11[256]},
      {stage1_12[148]},
      {stage1_13[117], stage1_13[118], stage1_13[119], stage1_13[120], stage1_13[121], stage1_13[122]},
      {stage2_15[37],stage2_14[38],stage2_13[56],stage2_12[72],stage2_11[114]}
   );
   gpc615_5 gpc6178 (
      {stage1_11[257], stage1_11[258], stage1_11[259], stage1_11[260], stage1_11[261]},
      {stage1_12[149]},
      {stage1_13[123], stage1_13[124], stage1_13[125], stage1_13[126], stage1_13[127], stage1_13[128]},
      {stage2_15[38],stage2_14[39],stage2_13[57],stage2_12[73],stage2_11[115]}
   );
   gpc615_5 gpc6179 (
      {stage1_11[262], stage1_11[263], stage1_11[264], stage1_11[265], stage1_11[266]},
      {stage1_12[150]},
      {stage1_13[129], stage1_13[130], stage1_13[131], stage1_13[132], stage1_13[133], stage1_13[134]},
      {stage2_15[39],stage2_14[40],stage2_13[58],stage2_12[74],stage2_11[116]}
   );
   gpc615_5 gpc6180 (
      {stage1_11[267], stage1_11[268], stage1_11[269], stage1_11[270], stage1_11[271]},
      {stage1_12[151]},
      {stage1_13[135], stage1_13[136], stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140]},
      {stage2_15[40],stage2_14[41],stage2_13[59],stage2_12[75],stage2_11[117]}
   );
   gpc615_5 gpc6181 (
      {stage1_11[272], stage1_11[273], stage1_11[274], stage1_11[275], stage1_11[276]},
      {stage1_12[152]},
      {stage1_13[141], stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage2_15[41],stage2_14[42],stage2_13[60],stage2_12[76],stage2_11[118]}
   );
   gpc615_5 gpc6182 (
      {stage1_11[277], stage1_11[278], stage1_11[279], stage1_11[280], stage1_11[281]},
      {stage1_12[153]},
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151], stage1_13[152]},
      {stage2_15[42],stage2_14[43],stage2_13[61],stage2_12[77],stage2_11[119]}
   );
   gpc615_5 gpc6183 (
      {stage1_11[282], stage1_11[283], stage1_11[284], stage1_11[285], stage1_11[286]},
      {stage1_12[154]},
      {stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158]},
      {stage2_15[43],stage2_14[44],stage2_13[62],stage2_12[78],stage2_11[120]}
   );
   gpc615_5 gpc6184 (
      {stage1_11[287], stage1_11[288], stage1_11[289], stage1_11[290], stage1_11[291]},
      {stage1_12[155]},
      {stage1_13[159], stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage2_15[44],stage2_14[45],stage2_13[63],stage2_12[79],stage2_11[121]}
   );
   gpc615_5 gpc6185 (
      {stage1_11[292], stage1_11[293], stage1_11[294], stage1_11[295], stage1_11[296]},
      {stage1_12[156]},
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170]},
      {stage2_15[45],stage2_14[46],stage2_13[64],stage2_12[80],stage2_11[122]}
   );
   gpc615_5 gpc6186 (
      {stage1_11[297], stage1_11[298], stage1_11[299], stage1_11[300], stage1_11[301]},
      {stage1_12[157]},
      {stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage2_15[46],stage2_14[47],stage2_13[65],stage2_12[81],stage2_11[123]}
   );
   gpc615_5 gpc6187 (
      {stage1_11[302], stage1_11[303], stage1_11[304], stage1_11[305], stage1_11[306]},
      {stage1_12[158]},
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181], stage1_13[182]},
      {stage2_15[47],stage2_14[48],stage2_13[66],stage2_12[82],stage2_11[124]}
   );
   gpc606_5 gpc6188 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26]},
      {stage2_16[0],stage2_15[48],stage2_14[49],stage2_13[67],stage2_12[83]}
   );
   gpc606_5 gpc6189 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31], stage1_14[32]},
      {stage2_16[1],stage2_15[49],stage2_14[50],stage2_13[68],stage2_12[84]}
   );
   gpc606_5 gpc6190 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37], stage1_14[38]},
      {stage2_16[2],stage2_15[50],stage2_14[51],stage2_13[69],stage2_12[85]}
   );
   gpc1163_5 gpc6191 (
      {stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[0],stage2_16[3],stage2_15[51],stage2_14[52]}
   );
   gpc1163_5 gpc6192 (
      {stage1_14[42], stage1_14[43], stage1_14[44]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[1]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[1],stage2_16[4],stage2_15[52],stage2_14[53]}
   );
   gpc1163_5 gpc6193 (
      {stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[2]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[2],stage2_16[5],stage2_15[53],stage2_14[54]}
   );
   gpc1163_5 gpc6194 (
      {stage1_14[48], stage1_14[49], stage1_14[50]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[3]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[3],stage2_16[6],stage2_15[54],stage2_14[55]}
   );
   gpc1163_5 gpc6195 (
      {stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[4]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[4],stage2_16[7],stage2_15[55],stage2_14[56]}
   );
   gpc1163_5 gpc6196 (
      {stage1_14[54], stage1_14[55], stage1_14[56]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[5]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[5],stage2_16[8],stage2_15[56],stage2_14[57]}
   );
   gpc1163_5 gpc6197 (
      {stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage1_16[6]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[6],stage2_16[9],stage2_15[57],stage2_14[58]}
   );
   gpc1163_5 gpc6198 (
      {stage1_14[60], stage1_14[61], stage1_14[62]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[7]},
      {stage1_17[7]},
      {stage2_18[7],stage2_17[7],stage2_16[10],stage2_15[58],stage2_14[59]}
   );
   gpc1163_5 gpc6199 (
      {stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[8]},
      {stage1_17[8]},
      {stage2_18[8],stage2_17[8],stage2_16[11],stage2_15[59],stage2_14[60]}
   );
   gpc1163_5 gpc6200 (
      {stage1_14[66], stage1_14[67], stage1_14[68]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage1_16[9]},
      {stage1_17[9]},
      {stage2_18[9],stage2_17[9],stage2_16[12],stage2_15[60],stage2_14[61]}
   );
   gpc1163_5 gpc6201 (
      {stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_16[10]},
      {stage1_17[10]},
      {stage2_18[10],stage2_17[10],stage2_16[13],stage2_15[61],stage2_14[62]}
   );
   gpc1163_5 gpc6202 (
      {stage1_14[72], stage1_14[73], stage1_14[74]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage1_16[11]},
      {stage1_17[11]},
      {stage2_18[11],stage2_17[11],stage2_16[14],stage2_15[62],stage2_14[63]}
   );
   gpc1163_5 gpc6203 (
      {stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[12]},
      {stage1_17[12]},
      {stage2_18[12],stage2_17[12],stage2_16[15],stage2_15[63],stage2_14[64]}
   );
   gpc1163_5 gpc6204 (
      {stage1_14[78], stage1_14[79], stage1_14[80]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[13]},
      {stage1_17[13]},
      {stage2_18[13],stage2_17[13],stage2_16[16],stage2_15[64],stage2_14[65]}
   );
   gpc1163_5 gpc6205 (
      {stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage1_16[14]},
      {stage1_17[14]},
      {stage2_18[14],stage2_17[14],stage2_16[17],stage2_15[65],stage2_14[66]}
   );
   gpc1163_5 gpc6206 (
      {stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage1_16[15]},
      {stage1_17[15]},
      {stage2_18[15],stage2_17[15],stage2_16[18],stage2_15[66],stage2_14[67]}
   );
   gpc1163_5 gpc6207 (
      {stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage1_16[16]},
      {stage1_17[16]},
      {stage2_18[16],stage2_17[16],stage2_16[19],stage2_15[67],stage2_14[68]}
   );
   gpc1163_5 gpc6208 (
      {stage1_14[90], stage1_14[91], stage1_14[92]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[17]},
      {stage1_17[17]},
      {stage2_18[17],stage2_17[17],stage2_16[20],stage2_15[68],stage2_14[69]}
   );
   gpc1163_5 gpc6209 (
      {stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage1_16[18]},
      {stage1_17[18]},
      {stage2_18[18],stage2_17[18],stage2_16[21],stage2_15[69],stage2_14[70]}
   );
   gpc1163_5 gpc6210 (
      {stage1_14[96], stage1_14[97], stage1_14[98]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage1_16[19]},
      {stage1_17[19]},
      {stage2_18[19],stage2_17[19],stage2_16[22],stage2_15[70],stage2_14[71]}
   );
   gpc1163_5 gpc6211 (
      {stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage1_16[20]},
      {stage1_17[20]},
      {stage2_18[20],stage2_17[20],stage2_16[23],stage2_15[71],stage2_14[72]}
   );
   gpc1163_5 gpc6212 (
      {stage1_14[102], stage1_14[103], stage1_14[104]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage1_16[21]},
      {stage1_17[21]},
      {stage2_18[21],stage2_17[21],stage2_16[24],stage2_15[72],stage2_14[73]}
   );
   gpc1163_5 gpc6213 (
      {stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage1_16[22]},
      {stage1_17[22]},
      {stage2_18[22],stage2_17[22],stage2_16[25],stage2_15[73],stage2_14[74]}
   );
   gpc1163_5 gpc6214 (
      {stage1_14[108], stage1_14[109], stage1_14[110]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage1_16[23]},
      {stage1_17[23]},
      {stage2_18[23],stage2_17[23],stage2_16[26],stage2_15[74],stage2_14[75]}
   );
   gpc1163_5 gpc6215 (
      {stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage1_16[24]},
      {stage1_17[24]},
      {stage2_18[24],stage2_17[24],stage2_16[27],stage2_15[75],stage2_14[76]}
   );
   gpc1163_5 gpc6216 (
      {stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage1_16[25]},
      {stage1_17[25]},
      {stage2_18[25],stage2_17[25],stage2_16[28],stage2_15[76],stage2_14[77]}
   );
   gpc1163_5 gpc6217 (
      {stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[26]},
      {stage1_17[26]},
      {stage2_18[26],stage2_17[26],stage2_16[29],stage2_15[77],stage2_14[78]}
   );
   gpc1163_5 gpc6218 (
      {stage1_14[120], stage1_14[121], stage1_14[122]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage1_16[27]},
      {stage1_17[27]},
      {stage2_18[27],stage2_17[27],stage2_16[30],stage2_15[78],stage2_14[79]}
   );
   gpc1163_5 gpc6219 (
      {stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage1_16[28]},
      {stage1_17[28]},
      {stage2_18[28],stage2_17[28],stage2_16[31],stage2_15[79],stage2_14[80]}
   );
   gpc1163_5 gpc6220 (
      {stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage1_16[29]},
      {stage1_17[29]},
      {stage2_18[29],stage2_17[29],stage2_16[32],stage2_15[80],stage2_14[81]}
   );
   gpc1163_5 gpc6221 (
      {stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage1_16[30]},
      {stage1_17[30]},
      {stage2_18[30],stage2_17[30],stage2_16[33],stage2_15[81],stage2_14[82]}
   );
   gpc1163_5 gpc6222 (
      {stage1_14[132], stage1_14[133], stage1_14[134]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[31]},
      {stage1_17[31]},
      {stage2_18[31],stage2_17[31],stage2_16[34],stage2_15[82],stage2_14[83]}
   );
   gpc606_5 gpc6223 (
      {stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140]},
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage2_18[32],stage2_17[32],stage2_16[35],stage2_15[83],stage2_14[84]}
   );
   gpc606_5 gpc6224 (
      {stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage2_18[33],stage2_17[33],stage2_16[36],stage2_15[84],stage2_14[85]}
   );
   gpc606_5 gpc6225 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152]},
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage2_18[34],stage2_17[34],stage2_16[37],stage2_15[85],stage2_14[86]}
   );
   gpc606_5 gpc6226 (
      {stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage2_18[35],stage2_17[35],stage2_16[38],stage2_15[86],stage2_14[87]}
   );
   gpc606_5 gpc6227 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163], stage1_14[164]},
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage2_18[36],stage2_17[36],stage2_16[39],stage2_15[87],stage2_14[88]}
   );
   gpc606_5 gpc6228 (
      {stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170]},
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage2_18[37],stage2_17[37],stage2_16[40],stage2_15[88],stage2_14[89]}
   );
   gpc615_5 gpc6229 (
      {stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_15[192]},
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage2_18[38],stage2_17[38],stage2_16[41],stage2_15[89],stage2_14[90]}
   );
   gpc615_5 gpc6230 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180]},
      {stage1_15[193]},
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage2_18[39],stage2_17[39],stage2_16[42],stage2_15[90],stage2_14[91]}
   );
   gpc615_5 gpc6231 (
      {stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage1_15[194]},
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage2_18[40],stage2_17[40],stage2_16[43],stage2_15[91],stage2_14[92]}
   );
   gpc615_5 gpc6232 (
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190]},
      {stage1_15[195]},
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage2_18[41],stage2_17[41],stage2_16[44],stage2_15[92],stage2_14[93]}
   );
   gpc615_5 gpc6233 (
      {stage1_14[191], stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195]},
      {stage1_15[196]},
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage2_18[42],stage2_17[42],stage2_16[45],stage2_15[93],stage2_14[94]}
   );
   gpc615_5 gpc6234 (
      {stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200]},
      {stage1_15[197]},
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage2_18[43],stage2_17[43],stage2_16[46],stage2_15[94],stage2_14[95]}
   );
   gpc615_5 gpc6235 (
      {stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_15[198]},
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage2_18[44],stage2_17[44],stage2_16[47],stage2_15[95],stage2_14[96]}
   );
   gpc615_5 gpc6236 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[199]},
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage2_18[45],stage2_17[45],stage2_16[48],stage2_15[96],stage2_14[97]}
   );
   gpc615_5 gpc6237 (
      {stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage1_15[200]},
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage2_18[46],stage2_17[46],stage2_16[49],stage2_15[97],stage2_14[98]}
   );
   gpc615_5 gpc6238 (
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220]},
      {stage1_15[201]},
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage2_18[47],stage2_17[47],stage2_16[50],stage2_15[98],stage2_14[99]}
   );
   gpc615_5 gpc6239 (
      {stage1_14[221], stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225]},
      {stage1_15[202]},
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage2_18[48],stage2_17[48],stage2_16[51],stage2_15[99],stage2_14[100]}
   );
   gpc615_5 gpc6240 (
      {stage1_14[226], stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230]},
      {stage1_15[203]},
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage2_18[49],stage2_17[49],stage2_16[52],stage2_15[100],stage2_14[101]}
   );
   gpc615_5 gpc6241 (
      {stage1_14[231], stage1_14[232], stage1_14[233], stage1_14[234], stage1_14[235]},
      {stage1_15[204]},
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage2_18[50],stage2_17[50],stage2_16[53],stage2_15[101],stage2_14[102]}
   );
   gpc615_5 gpc6242 (
      {stage1_14[236], stage1_14[237], stage1_14[238], stage1_14[239], stage1_14[240]},
      {stage1_15[205]},
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage2_18[51],stage2_17[51],stage2_16[54],stage2_15[102],stage2_14[103]}
   );
   gpc615_5 gpc6243 (
      {stage1_14[241], stage1_14[242], stage1_14[243], stage1_14[244], stage1_14[245]},
      {stage1_15[206]},
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage2_18[52],stage2_17[52],stage2_16[55],stage2_15[103],stage2_14[104]}
   );
   gpc1406_5 gpc6244 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211], stage1_15[212]},
      {stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[53],stage2_17[53],stage2_16[56],stage2_15[104]}
   );
   gpc1406_5 gpc6245 (
      {stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216], stage1_15[217], stage1_15[218]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39]},
      {stage1_18[1]},
      {stage2_19[1],stage2_18[54],stage2_17[54],stage2_16[57],stage2_15[105]}
   );
   gpc606_5 gpc6246 (
      {stage1_15[219], stage1_15[220], stage1_15[221], stage1_15[222], stage1_15[223], stage1_15[224]},
      {stage1_17[40], stage1_17[41], stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45]},
      {stage2_19[2],stage2_18[55],stage2_17[55],stage2_16[58],stage2_15[106]}
   );
   gpc606_5 gpc6247 (
      {stage1_15[225], stage1_15[226], stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230]},
      {stage1_17[46], stage1_17[47], stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51]},
      {stage2_19[3],stage2_18[56],stage2_17[56],stage2_16[59],stage2_15[107]}
   );
   gpc606_5 gpc6248 (
      {stage1_15[231], stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_17[52], stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage2_19[4],stage2_18[57],stage2_17[57],stage2_16[60],stage2_15[108]}
   );
   gpc606_5 gpc6249 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241], stage1_15[242]},
      {stage1_17[58], stage1_17[59], stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63]},
      {stage2_19[5],stage2_18[58],stage2_17[58],stage2_16[61],stage2_15[109]}
   );
   gpc606_5 gpc6250 (
      {stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246], stage1_15[247], stage1_15[248]},
      {stage1_17[64], stage1_17[65], stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69]},
      {stage2_19[6],stage2_18[59],stage2_17[59],stage2_16[62],stage2_15[110]}
   );
   gpc606_5 gpc6251 (
      {stage1_15[249], stage1_15[250], stage1_15[251], stage1_15[252], stage1_15[253], stage1_15[254]},
      {stage1_17[70], stage1_17[71], stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75]},
      {stage2_19[7],stage2_18[60],stage2_17[60],stage2_16[63],stage2_15[111]}
   );
   gpc606_5 gpc6252 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6], stage1_18[7]},
      {stage2_20[0],stage2_19[8],stage2_18[61],stage2_17[61],stage2_16[64]}
   );
   gpc606_5 gpc6253 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12], stage1_18[13]},
      {stage2_20[1],stage2_19[9],stage2_18[62],stage2_17[62],stage2_16[65]}
   );
   gpc606_5 gpc6254 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18], stage1_18[19]},
      {stage2_20[2],stage2_19[10],stage2_18[63],stage2_17[63],stage2_16[66]}
   );
   gpc606_5 gpc6255 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180], stage1_16[181]},
      {stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25]},
      {stage2_20[3],stage2_19[11],stage2_18[64],stage2_17[64],stage2_16[67]}
   );
   gpc606_5 gpc6256 (
      {stage1_17[76], stage1_17[77], stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[4],stage2_19[12],stage2_18[65],stage2_17[65]}
   );
   gpc606_5 gpc6257 (
      {stage1_17[82], stage1_17[83], stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[5],stage2_19[13],stage2_18[66],stage2_17[66]}
   );
   gpc606_5 gpc6258 (
      {stage1_17[88], stage1_17[89], stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[6],stage2_19[14],stage2_18[67],stage2_17[67]}
   );
   gpc606_5 gpc6259 (
      {stage1_17[94], stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[7],stage2_19[15],stage2_18[68],stage2_17[68]}
   );
   gpc606_5 gpc6260 (
      {stage1_17[100], stage1_17[101], stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[8],stage2_19[16],stage2_18[69],stage2_17[69]}
   );
   gpc606_5 gpc6261 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[9],stage2_19[17],stage2_18[70],stage2_17[70]}
   );
   gpc606_5 gpc6262 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[10],stage2_19[18],stage2_18[71],stage2_17[71]}
   );
   gpc606_5 gpc6263 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[11],stage2_19[19],stage2_18[72],stage2_17[72]}
   );
   gpc606_5 gpc6264 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[12],stage2_19[20],stage2_18[73],stage2_17[73]}
   );
   gpc606_5 gpc6265 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[13],stage2_19[21],stage2_18[74],stage2_17[74]}
   );
   gpc606_5 gpc6266 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[14],stage2_19[22],stage2_18[75],stage2_17[75]}
   );
   gpc606_5 gpc6267 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[15],stage2_19[23],stage2_18[76],stage2_17[76]}
   );
   gpc606_5 gpc6268 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[16],stage2_19[24],stage2_18[77],stage2_17[77]}
   );
   gpc606_5 gpc6269 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[17],stage2_19[25],stage2_18[78],stage2_17[78]}
   );
   gpc606_5 gpc6270 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[18],stage2_19[26],stage2_18[79],stage2_17[79]}
   );
   gpc606_5 gpc6271 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[19],stage2_19[27],stage2_18[80],stage2_17[80]}
   );
   gpc606_5 gpc6272 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[20],stage2_19[28],stage2_18[81],stage2_17[81]}
   );
   gpc606_5 gpc6273 (
      {stage1_17[178], stage1_17[179], stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[21],stage2_19[29],stage2_18[82],stage2_17[82]}
   );
   gpc606_5 gpc6274 (
      {stage1_17[184], stage1_17[185], stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[22],stage2_19[30],stage2_18[83],stage2_17[83]}
   );
   gpc606_5 gpc6275 (
      {stage1_17[190], stage1_17[191], stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[23],stage2_19[31],stage2_18[84],stage2_17[84]}
   );
   gpc606_5 gpc6276 (
      {stage1_17[196], stage1_17[197], stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[24],stage2_19[32],stage2_18[85],stage2_17[85]}
   );
   gpc606_5 gpc6277 (
      {stage1_17[202], stage1_17[203], stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[25],stage2_19[33],stage2_18[86],stage2_17[86]}
   );
   gpc606_5 gpc6278 (
      {stage1_17[208], stage1_17[209], stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[26],stage2_19[34],stage2_18[87],stage2_17[87]}
   );
   gpc606_5 gpc6279 (
      {stage1_17[214], stage1_17[215], stage1_17[216], stage1_17[217], 1'b0, 1'b0},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[27],stage2_19[35],stage2_18[88],stage2_17[88]}
   );
   gpc606_5 gpc6280 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[28],stage2_19[36],stage2_18[89],stage2_17[89]}
   );
   gpc606_5 gpc6281 (
      {stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[25],stage2_20[29],stage2_19[37],stage2_18[90]}
   );
   gpc606_5 gpc6282 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36], stage1_18[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[26],stage2_20[30],stage2_19[38],stage2_18[91]}
   );
   gpc606_5 gpc6283 (
      {stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42], stage1_18[43]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[27],stage2_20[31],stage2_19[39],stage2_18[92]}
   );
   gpc606_5 gpc6284 (
      {stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48], stage1_18[49]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[28],stage2_20[32],stage2_19[40],stage2_18[93]}
   );
   gpc606_5 gpc6285 (
      {stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54], stage1_18[55]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[29],stage2_20[33],stage2_19[41],stage2_18[94]}
   );
   gpc606_5 gpc6286 (
      {stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[30],stage2_20[34],stage2_19[42],stage2_18[95]}
   );
   gpc606_5 gpc6287 (
      {stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[31],stage2_20[35],stage2_19[43],stage2_18[96]}
   );
   gpc606_5 gpc6288 (
      {stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[32],stage2_20[36],stage2_19[44],stage2_18[97]}
   );
   gpc615_5 gpc6289 (
      {stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77], stage1_18[78]},
      {stage1_19[150]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[33],stage2_20[37],stage2_19[45],stage2_18[98]}
   );
   gpc615_5 gpc6290 (
      {stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_19[151]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[34],stage2_20[38],stage2_19[46],stage2_18[99]}
   );
   gpc615_5 gpc6291 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[152]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[35],stage2_20[39],stage2_19[47],stage2_18[100]}
   );
   gpc615_5 gpc6292 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[153]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[36],stage2_20[40],stage2_19[48],stage2_18[101]}
   );
   gpc615_5 gpc6293 (
      {stage1_18[94], stage1_18[95], stage1_18[96], stage1_18[97], stage1_18[98]},
      {stage1_19[154]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[37],stage2_20[41],stage2_19[49],stage2_18[102]}
   );
   gpc615_5 gpc6294 (
      {stage1_18[99], stage1_18[100], stage1_18[101], stage1_18[102], stage1_18[103]},
      {stage1_19[155]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[38],stage2_20[42],stage2_19[50],stage2_18[103]}
   );
   gpc615_5 gpc6295 (
      {stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107], stage1_18[108]},
      {stage1_19[156]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[39],stage2_20[43],stage2_19[51],stage2_18[104]}
   );
   gpc615_5 gpc6296 (
      {stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_19[157]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[40],stage2_20[44],stage2_19[52],stage2_18[105]}
   );
   gpc615_5 gpc6297 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118]},
      {stage1_19[158]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[41],stage2_20[45],stage2_19[53],stage2_18[106]}
   );
   gpc615_5 gpc6298 (
      {stage1_18[119], stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123]},
      {stage1_19[159]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[42],stage2_20[46],stage2_19[54],stage2_18[107]}
   );
   gpc615_5 gpc6299 (
      {stage1_18[124], stage1_18[125], stage1_18[126], stage1_18[127], stage1_18[128]},
      {stage1_19[160]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[43],stage2_20[47],stage2_19[55],stage2_18[108]}
   );
   gpc615_5 gpc6300 (
      {stage1_18[129], stage1_18[130], stage1_18[131], stage1_18[132], stage1_18[133]},
      {stage1_19[161]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[44],stage2_20[48],stage2_19[56],stage2_18[109]}
   );
   gpc615_5 gpc6301 (
      {stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137], stage1_18[138]},
      {stage1_19[162]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[45],stage2_20[49],stage2_19[57],stage2_18[110]}
   );
   gpc615_5 gpc6302 (
      {stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_19[163]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[46],stage2_20[50],stage2_19[58],stage2_18[111]}
   );
   gpc615_5 gpc6303 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148]},
      {stage1_19[164]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[47],stage2_20[51],stage2_19[59],stage2_18[112]}
   );
   gpc615_5 gpc6304 (
      {stage1_18[149], stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153]},
      {stage1_19[165]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[48],stage2_20[52],stage2_19[60],stage2_18[113]}
   );
   gpc615_5 gpc6305 (
      {stage1_18[154], stage1_18[155], stage1_18[156], stage1_18[157], stage1_18[158]},
      {stage1_19[166]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[49],stage2_20[53],stage2_19[61],stage2_18[114]}
   );
   gpc615_5 gpc6306 (
      {stage1_18[159], stage1_18[160], stage1_18[161], stage1_18[162], stage1_18[163]},
      {stage1_19[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[50],stage2_20[54],stage2_19[62],stage2_18[115]}
   );
   gpc615_5 gpc6307 (
      {stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167], stage1_18[168]},
      {stage1_19[168]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[51],stage2_20[55],stage2_19[63],stage2_18[116]}
   );
   gpc615_5 gpc6308 (
      {stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_19[169]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[52],stage2_20[56],stage2_19[64],stage2_18[117]}
   );
   gpc615_5 gpc6309 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[170]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[53],stage2_20[57],stage2_19[65],stage2_18[118]}
   );
   gpc615_5 gpc6310 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[171]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[54],stage2_20[58],stage2_19[66],stage2_18[119]}
   );
   gpc615_5 gpc6311 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[172]},
      {stage1_20[180], stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185]},
      {stage2_22[30],stage2_21[55],stage2_20[59],stage2_19[67],stage2_18[120]}
   );
   gpc615_5 gpc6312 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[173]},
      {stage1_20[186], stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage2_22[31],stage2_21[56],stage2_20[60],stage2_19[68],stage2_18[121]}
   );
   gpc615_5 gpc6313 (
      {stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197], stage1_18[198]},
      {stage1_19[174]},
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197]},
      {stage2_22[32],stage2_21[57],stage2_20[61],stage2_19[69],stage2_18[122]}
   );
   gpc615_5 gpc6314 (
      {stage1_18[199], stage1_18[200], stage1_18[201], stage1_18[202], stage1_18[203]},
      {stage1_19[175]},
      {stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203]},
      {stage2_22[33],stage2_21[58],stage2_20[62],stage2_19[70],stage2_18[123]}
   );
   gpc615_5 gpc6315 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[204]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[34],stage2_21[59],stage2_20[63],stage2_19[71]}
   );
   gpc615_5 gpc6316 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[205]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[35],stage2_21[60],stage2_20[64],stage2_19[72]}
   );
   gpc615_5 gpc6317 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[206]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[36],stage2_21[61],stage2_20[65],stage2_19[73]}
   );
   gpc615_5 gpc6318 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[207]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[37],stage2_21[62],stage2_20[66],stage2_19[74]}
   );
   gpc615_5 gpc6319 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[208]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[38],stage2_21[63],stage2_20[67],stage2_19[75]}
   );
   gpc606_5 gpc6320 (
      {stage1_20[209], stage1_20[210], stage1_20[211], stage1_20[212], stage1_20[213], stage1_20[214]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[39],stage2_21[64],stage2_20[68]}
   );
   gpc606_5 gpc6321 (
      {stage1_20[215], stage1_20[216], stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[40],stage2_21[65],stage2_20[69]}
   );
   gpc606_5 gpc6322 (
      {stage1_20[221], stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[41],stage2_21[66],stage2_20[70]}
   );
   gpc606_5 gpc6323 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[3],stage2_23[8],stage2_22[42],stage2_21[67]}
   );
   gpc606_5 gpc6324 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[4],stage2_23[9],stage2_22[43],stage2_21[68]}
   );
   gpc606_5 gpc6325 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[5],stage2_23[10],stage2_22[44],stage2_21[69]}
   );
   gpc606_5 gpc6326 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[6],stage2_23[11],stage2_22[45],stage2_21[70]}
   );
   gpc606_5 gpc6327 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[7],stage2_23[12],stage2_22[46],stage2_21[71]}
   );
   gpc606_5 gpc6328 (
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[8],stage2_23[13],stage2_22[47],stage2_21[72]}
   );
   gpc606_5 gpc6329 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[9],stage2_23[14],stage2_22[48],stage2_21[73]}
   );
   gpc606_5 gpc6330 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[10],stage2_23[15],stage2_22[49],stage2_21[74]}
   );
   gpc606_5 gpc6331 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[11],stage2_23[16],stage2_22[50],stage2_21[75]}
   );
   gpc606_5 gpc6332 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[12],stage2_23[17],stage2_22[51],stage2_21[76]}
   );
   gpc606_5 gpc6333 (
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[13],stage2_23[18],stage2_22[52],stage2_21[77]}
   );
   gpc606_5 gpc6334 (
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[14],stage2_23[19],stage2_22[53],stage2_21[78]}
   );
   gpc606_5 gpc6335 (
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[15],stage2_23[20],stage2_22[54],stage2_21[79]}
   );
   gpc606_5 gpc6336 (
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[16],stage2_23[21],stage2_22[55],stage2_21[80]}
   );
   gpc606_5 gpc6337 (
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[17],stage2_23[22],stage2_22[56],stage2_21[81]}
   );
   gpc606_5 gpc6338 (
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[18],stage2_23[23],stage2_22[57],stage2_21[82]}
   );
   gpc606_5 gpc6339 (
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[19],stage2_23[24],stage2_22[58],stage2_21[83]}
   );
   gpc606_5 gpc6340 (
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[20],stage2_23[25],stage2_22[59],stage2_21[84]}
   );
   gpc606_5 gpc6341 (
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[21],stage2_23[26],stage2_22[60],stage2_21[85]}
   );
   gpc606_5 gpc6342 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[22],stage2_23[27],stage2_22[61],stage2_21[86]}
   );
   gpc606_5 gpc6343 (
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[23],stage2_23[28],stage2_22[62],stage2_21[87]}
   );
   gpc606_5 gpc6344 (
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[24],stage2_23[29],stage2_22[63],stage2_21[88]}
   );
   gpc606_5 gpc6345 (
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[25],stage2_23[30],stage2_22[64],stage2_21[89]}
   );
   gpc606_5 gpc6346 (
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[26],stage2_23[31],stage2_22[65],stage2_21[90]}
   );
   gpc606_5 gpc6347 (
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[27],stage2_23[32],stage2_22[66],stage2_21[91]}
   );
   gpc606_5 gpc6348 (
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[28],stage2_23[33],stage2_22[67],stage2_21[92]}
   );
   gpc606_5 gpc6349 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[26],stage2_24[29],stage2_23[34],stage2_22[68]}
   );
   gpc615_5 gpc6350 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[156]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[27],stage2_24[30],stage2_23[35],stage2_22[69]}
   );
   gpc615_5 gpc6351 (
      {stage1_22[29], stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33]},
      {stage1_23[157]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[28],stage2_24[31],stage2_23[36],stage2_22[70]}
   );
   gpc615_5 gpc6352 (
      {stage1_22[34], stage1_22[35], stage1_22[36], stage1_22[37], stage1_22[38]},
      {stage1_23[158]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[29],stage2_24[32],stage2_23[37],stage2_22[71]}
   );
   gpc615_5 gpc6353 (
      {stage1_22[39], stage1_22[40], stage1_22[41], stage1_22[42], stage1_22[43]},
      {stage1_23[159]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[30],stage2_24[33],stage2_23[38],stage2_22[72]}
   );
   gpc615_5 gpc6354 (
      {stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47], stage1_22[48]},
      {stage1_23[160]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[31],stage2_24[34],stage2_23[39],stage2_22[73]}
   );
   gpc615_5 gpc6355 (
      {stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_23[161]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[32],stage2_24[35],stage2_23[40],stage2_22[74]}
   );
   gpc615_5 gpc6356 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58]},
      {stage1_23[162]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[33],stage2_24[36],stage2_23[41],stage2_22[75]}
   );
   gpc615_5 gpc6357 (
      {stage1_22[59], stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63]},
      {stage1_23[163]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[34],stage2_24[37],stage2_23[42],stage2_22[76]}
   );
   gpc615_5 gpc6358 (
      {stage1_22[64], stage1_22[65], stage1_22[66], stage1_22[67], stage1_22[68]},
      {stage1_23[164]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[35],stage2_24[38],stage2_23[43],stage2_22[77]}
   );
   gpc615_5 gpc6359 (
      {stage1_22[69], stage1_22[70], stage1_22[71], stage1_22[72], stage1_22[73]},
      {stage1_23[165]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[36],stage2_24[39],stage2_23[44],stage2_22[78]}
   );
   gpc615_5 gpc6360 (
      {stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77], stage1_22[78]},
      {stage1_23[166]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[37],stage2_24[40],stage2_23[45],stage2_22[79]}
   );
   gpc615_5 gpc6361 (
      {stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage1_23[167]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[38],stage2_24[41],stage2_23[46],stage2_22[80]}
   );
   gpc615_5 gpc6362 (
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88]},
      {stage1_23[168]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[39],stage2_24[42],stage2_23[47],stage2_22[81]}
   );
   gpc615_5 gpc6363 (
      {stage1_22[89], stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93]},
      {stage1_23[169]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[40],stage2_24[43],stage2_23[48],stage2_22[82]}
   );
   gpc615_5 gpc6364 (
      {stage1_22[94], stage1_22[95], stage1_22[96], stage1_22[97], stage1_22[98]},
      {stage1_23[170]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[41],stage2_24[44],stage2_23[49],stage2_22[83]}
   );
   gpc615_5 gpc6365 (
      {stage1_22[99], stage1_22[100], stage1_22[101], stage1_22[102], stage1_22[103]},
      {stage1_23[171]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[42],stage2_24[45],stage2_23[50],stage2_22[84]}
   );
   gpc615_5 gpc6366 (
      {stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108]},
      {stage1_23[172]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[43],stage2_24[46],stage2_23[51],stage2_22[85]}
   );
   gpc615_5 gpc6367 (
      {stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage1_23[173]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[44],stage2_24[47],stage2_23[52],stage2_22[86]}
   );
   gpc615_5 gpc6368 (
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118]},
      {stage1_23[174]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[45],stage2_24[48],stage2_23[53],stage2_22[87]}
   );
   gpc615_5 gpc6369 (
      {stage1_22[119], stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123]},
      {stage1_23[175]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[46],stage2_24[49],stage2_23[54],stage2_22[88]}
   );
   gpc615_5 gpc6370 (
      {stage1_22[124], stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128]},
      {stage1_23[176]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[47],stage2_24[50],stage2_23[55],stage2_22[89]}
   );
   gpc615_5 gpc6371 (
      {stage1_22[129], stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133]},
      {stage1_23[177]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[48],stage2_24[51],stage2_23[56],stage2_22[90]}
   );
   gpc615_5 gpc6372 (
      {stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138]},
      {stage1_23[178]},
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage2_26[23],stage2_25[49],stage2_24[52],stage2_23[57],stage2_22[91]}
   );
   gpc615_5 gpc6373 (
      {stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage1_23[179]},
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage2_26[24],stage2_25[50],stage2_24[53],stage2_23[58],stage2_22[92]}
   );
   gpc615_5 gpc6374 (
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148]},
      {stage1_23[180]},
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage2_26[25],stage2_25[51],stage2_24[54],stage2_23[59],stage2_22[93]}
   );
   gpc615_5 gpc6375 (
      {stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153]},
      {stage1_23[181]},
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage2_26[26],stage2_25[52],stage2_24[55],stage2_23[60],stage2_22[94]}
   );
   gpc615_5 gpc6376 (
      {stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157], stage1_22[158]},
      {stage1_23[182]},
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage2_26[27],stage2_25[53],stage2_24[56],stage2_23[61],stage2_22[95]}
   );
   gpc615_5 gpc6377 (
      {stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162], stage1_22[163]},
      {stage1_23[183]},
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage2_26[28],stage2_25[54],stage2_24[57],stage2_23[62],stage2_22[96]}
   );
   gpc615_5 gpc6378 (
      {stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167], stage1_22[168]},
      {stage1_23[184]},
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage2_26[29],stage2_25[55],stage2_24[58],stage2_23[63],stage2_22[97]}
   );
   gpc615_5 gpc6379 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173]},
      {stage1_23[185]},
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage2_26[30],stage2_25[56],stage2_24[59],stage2_23[64],stage2_22[98]}
   );
   gpc615_5 gpc6380 (
      {stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178]},
      {stage1_23[186]},
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage2_26[31],stage2_25[57],stage2_24[60],stage2_23[65],stage2_22[99]}
   );
   gpc615_5 gpc6381 (
      {stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182], stage1_22[183]},
      {stage1_23[187]},
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage2_26[32],stage2_25[58],stage2_24[61],stage2_23[66],stage2_22[100]}
   );
   gpc615_5 gpc6382 (
      {stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187], stage1_22[188]},
      {stage1_23[188]},
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage2_26[33],stage2_25[59],stage2_24[62],stage2_23[67],stage2_22[101]}
   );
   gpc615_5 gpc6383 (
      {stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192], stage1_22[193]},
      {stage1_23[189]},
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage2_26[34],stage2_25[60],stage2_24[63],stage2_23[68],stage2_22[102]}
   );
   gpc615_5 gpc6384 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[210]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[35],stage2_25[61],stage2_24[64],stage2_23[69]}
   );
   gpc615_5 gpc6385 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[211]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[36],stage2_25[62],stage2_24[65],stage2_23[70]}
   );
   gpc615_5 gpc6386 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[212]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[37],stage2_25[63],stage2_24[66],stage2_23[71]}
   );
   gpc615_5 gpc6387 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[213]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[38],stage2_25[64],stage2_24[67],stage2_23[72]}
   );
   gpc615_5 gpc6388 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[214]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[39],stage2_25[65],stage2_24[68],stage2_23[73]}
   );
   gpc615_5 gpc6389 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[215]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[40],stage2_25[66],stage2_24[69],stage2_23[74]}
   );
   gpc615_5 gpc6390 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[216]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[41],stage2_25[67],stage2_24[70],stage2_23[75]}
   );
   gpc615_5 gpc6391 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[217]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[42],stage2_25[68],stage2_24[71],stage2_23[76]}
   );
   gpc615_5 gpc6392 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[218]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[43],stage2_25[69],stage2_24[72],stage2_23[77]}
   );
   gpc615_5 gpc6393 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[219]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[44],stage2_25[70],stage2_24[73],stage2_23[78]}
   );
   gpc615_5 gpc6394 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[220]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[45],stage2_25[71],stage2_24[74],stage2_23[79]}
   );
   gpc615_5 gpc6395 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[221]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[46],stage2_25[72],stage2_24[75],stage2_23[80]}
   );
   gpc615_5 gpc6396 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[222]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[47],stage2_25[73],stage2_24[76],stage2_23[81]}
   );
   gpc615_5 gpc6397 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[223]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[48],stage2_25[74],stage2_24[77],stage2_23[82]}
   );
   gpc615_5 gpc6398 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[224]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[49],stage2_25[75],stage2_24[78],stage2_23[83]}
   );
   gpc615_5 gpc6399 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[225]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[50],stage2_25[76],stage2_24[79],stage2_23[84]}
   );
   gpc615_5 gpc6400 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[226]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[51],stage2_25[77],stage2_24[80],stage2_23[85]}
   );
   gpc615_5 gpc6401 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[227]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[52],stage2_25[78],stage2_24[81],stage2_23[86]}
   );
   gpc615_5 gpc6402 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[228]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[53],stage2_25[79],stage2_24[82],stage2_23[87]}
   );
   gpc615_5 gpc6403 (
      {stage1_23[285], stage1_23[286], stage1_23[287], stage1_23[288], stage1_23[289]},
      {stage1_24[229]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[54],stage2_25[80],stage2_24[83],stage2_23[88]}
   );
   gpc606_5 gpc6404 (
      {stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233], stage1_24[234], 1'b0},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[20],stage2_26[55],stage2_25[81],stage2_24[84]}
   );
   gpc606_5 gpc6405 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[1],stage2_27[21],stage2_26[56],stage2_25[82]}
   );
   gpc606_5 gpc6406 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[2],stage2_27[22],stage2_26[57],stage2_25[83]}
   );
   gpc606_5 gpc6407 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[3],stage2_27[23],stage2_26[58],stage2_25[84]}
   );
   gpc606_5 gpc6408 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[4],stage2_27[24],stage2_26[59],stage2_25[85]}
   );
   gpc606_5 gpc6409 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[5],stage2_27[25],stage2_26[60],stage2_25[86]}
   );
   gpc606_5 gpc6410 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[6],stage2_27[26],stage2_26[61],stage2_25[87]}
   );
   gpc606_5 gpc6411 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[7],stage2_27[27],stage2_26[62],stage2_25[88]}
   );
   gpc606_5 gpc6412 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[8],stage2_27[28],stage2_26[63],stage2_25[89]}
   );
   gpc606_5 gpc6413 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[9],stage2_27[29],stage2_26[64],stage2_25[90]}
   );
   gpc606_5 gpc6414 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[10],stage2_27[30],stage2_26[65],stage2_25[91]}
   );
   gpc615_5 gpc6415 (
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10]},
      {stage1_27[60]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[10],stage2_28[11],stage2_27[31],stage2_26[66]}
   );
   gpc615_5 gpc6416 (
      {stage1_26[11], stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15]},
      {stage1_27[61]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[11],stage2_28[12],stage2_27[32],stage2_26[67]}
   );
   gpc615_5 gpc6417 (
      {stage1_26[16], stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20]},
      {stage1_27[62]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[12],stage2_28[13],stage2_27[33],stage2_26[68]}
   );
   gpc615_5 gpc6418 (
      {stage1_26[21], stage1_26[22], stage1_26[23], stage1_26[24], stage1_26[25]},
      {stage1_27[63]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[13],stage2_28[14],stage2_27[34],stage2_26[69]}
   );
   gpc615_5 gpc6419 (
      {stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29], stage1_26[30]},
      {stage1_27[64]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[14],stage2_28[15],stage2_27[35],stage2_26[70]}
   );
   gpc615_5 gpc6420 (
      {stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[65]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[15],stage2_28[16],stage2_27[36],stage2_26[71]}
   );
   gpc615_5 gpc6421 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40]},
      {stage1_27[66]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[16],stage2_28[17],stage2_27[37],stage2_26[72]}
   );
   gpc615_5 gpc6422 (
      {stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45]},
      {stage1_27[67]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[17],stage2_28[18],stage2_27[38],stage2_26[73]}
   );
   gpc615_5 gpc6423 (
      {stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49], stage1_26[50]},
      {stage1_27[68]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[18],stage2_28[19],stage2_27[39],stage2_26[74]}
   );
   gpc615_5 gpc6424 (
      {stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54], stage1_26[55]},
      {stage1_27[69]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[19],stage2_28[20],stage2_27[40],stage2_26[75]}
   );
   gpc615_5 gpc6425 (
      {stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59], stage1_26[60]},
      {stage1_27[70]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[20],stage2_28[21],stage2_27[41],stage2_26[76]}
   );
   gpc615_5 gpc6426 (
      {stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage1_27[71]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[21],stage2_28[22],stage2_27[42],stage2_26[77]}
   );
   gpc615_5 gpc6427 (
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70]},
      {stage1_27[72]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[22],stage2_28[23],stage2_27[43],stage2_26[78]}
   );
   gpc615_5 gpc6428 (
      {stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75]},
      {stage1_27[73]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[23],stage2_28[24],stage2_27[44],stage2_26[79]}
   );
   gpc615_5 gpc6429 (
      {stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79], stage1_26[80]},
      {stage1_27[74]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[24],stage2_28[25],stage2_27[45],stage2_26[80]}
   );
   gpc615_5 gpc6430 (
      {stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84], stage1_26[85]},
      {stage1_27[75]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[25],stage2_28[26],stage2_27[46],stage2_26[81]}
   );
   gpc615_5 gpc6431 (
      {stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89], stage1_26[90]},
      {stage1_27[76]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[26],stage2_28[27],stage2_27[47],stage2_26[82]}
   );
   gpc615_5 gpc6432 (
      {stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage1_27[77]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[27],stage2_28[28],stage2_27[48],stage2_26[83]}
   );
   gpc615_5 gpc6433 (
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100]},
      {stage1_27[78]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[28],stage2_28[29],stage2_27[49],stage2_26[84]}
   );
   gpc615_5 gpc6434 (
      {stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105]},
      {stage1_27[79]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[29],stage2_28[30],stage2_27[50],stage2_26[85]}
   );
   gpc615_5 gpc6435 (
      {stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109], stage1_26[110]},
      {stage1_27[80]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[30],stage2_28[31],stage2_27[51],stage2_26[86]}
   );
   gpc615_5 gpc6436 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[81]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[31],stage2_28[32],stage2_27[52],stage2_26[87]}
   );
   gpc615_5 gpc6437 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[82]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[32],stage2_28[33],stage2_27[53],stage2_26[88]}
   );
   gpc615_5 gpc6438 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[83]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[33],stage2_28[34],stage2_27[54],stage2_26[89]}
   );
   gpc615_5 gpc6439 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[84]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[34],stage2_28[35],stage2_27[55],stage2_26[90]}
   );
   gpc615_5 gpc6440 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[85]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[35],stage2_28[36],stage2_27[56],stage2_26[91]}
   );
   gpc615_5 gpc6441 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[86]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[36],stage2_28[37],stage2_27[57],stage2_26[92]}
   );
   gpc615_5 gpc6442 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[87]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[37],stage2_28[38],stage2_27[58],stage2_26[93]}
   );
   gpc615_5 gpc6443 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[88]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[38],stage2_28[39],stage2_27[59],stage2_26[94]}
   );
   gpc623_5 gpc6444 (
      {stage1_26[151], stage1_26[152], stage1_26[153]},
      {stage1_27[89], stage1_27[90]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[39],stage2_28[40],stage2_27[60],stage2_26[95]}
   );
   gpc615_5 gpc6445 (
      {stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage1_28[180]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[30],stage2_29[40],stage2_28[41],stage2_27[61]}
   );
   gpc615_5 gpc6446 (
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100]},
      {stage1_28[181]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[31],stage2_29[41],stage2_28[42],stage2_27[62]}
   );
   gpc615_5 gpc6447 (
      {stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105]},
      {stage1_28[182]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[32],stage2_29[42],stage2_28[43],stage2_27[63]}
   );
   gpc615_5 gpc6448 (
      {stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109], stage1_27[110]},
      {stage1_28[183]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[33],stage2_29[43],stage2_28[44],stage2_27[64]}
   );
   gpc615_5 gpc6449 (
      {stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114], stage1_27[115]},
      {stage1_28[184]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[34],stage2_29[44],stage2_28[45],stage2_27[65]}
   );
   gpc615_5 gpc6450 (
      {stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119], stage1_27[120]},
      {stage1_28[185]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[35],stage2_29[45],stage2_28[46],stage2_27[66]}
   );
   gpc615_5 gpc6451 (
      {stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage1_28[186]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[36],stage2_29[46],stage2_28[47],stage2_27[67]}
   );
   gpc615_5 gpc6452 (
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130]},
      {stage1_28[187]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[37],stage2_29[47],stage2_28[48],stage2_27[68]}
   );
   gpc615_5 gpc6453 (
      {stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135]},
      {stage1_28[188]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[38],stage2_29[48],stage2_28[49],stage2_27[69]}
   );
   gpc615_5 gpc6454 (
      {stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139], stage1_27[140]},
      {stage1_28[189]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[39],stage2_29[49],stage2_28[50],stage2_27[70]}
   );
   gpc615_5 gpc6455 (
      {stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144], stage1_27[145]},
      {stage1_28[190]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[40],stage2_29[50],stage2_28[51],stage2_27[71]}
   );
   gpc615_5 gpc6456 (
      {stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149], stage1_27[150]},
      {stage1_28[191]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[41],stage2_29[51],stage2_28[52],stage2_27[72]}
   );
   gpc615_5 gpc6457 (
      {stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage1_28[192]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[42],stage2_29[52],stage2_28[53],stage2_27[73]}
   );
   gpc615_5 gpc6458 (
      {stage1_27[156], stage1_27[157], stage1_27[158], stage1_27[159], stage1_27[160]},
      {stage1_28[193]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[43],stage2_29[53],stage2_28[54],stage2_27[74]}
   );
   gpc615_5 gpc6459 (
      {stage1_27[161], stage1_27[162], stage1_27[163], stage1_27[164], stage1_27[165]},
      {stage1_28[194]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[44],stage2_29[54],stage2_28[55],stage2_27[75]}
   );
   gpc615_5 gpc6460 (
      {stage1_27[166], stage1_27[167], stage1_27[168], stage1_27[169], stage1_27[170]},
      {stage1_28[195]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[45],stage2_29[55],stage2_28[56],stage2_27[76]}
   );
   gpc615_5 gpc6461 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[196]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[46],stage2_29[56],stage2_28[57],stage2_27[77]}
   );
   gpc615_5 gpc6462 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[197]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[47],stage2_29[57],stage2_28[58],stage2_27[78]}
   );
   gpc615_5 gpc6463 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[198]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[48],stage2_29[58],stage2_28[59],stage2_27[79]}
   );
   gpc615_5 gpc6464 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[199]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[49],stage2_29[59],stage2_28[60],stage2_27[80]}
   );
   gpc615_5 gpc6465 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[200]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[50],stage2_29[60],stage2_28[61],stage2_27[81]}
   );
   gpc615_5 gpc6466 (
      {stage1_27[196], stage1_27[197], stage1_27[198], stage1_27[199], stage1_27[200]},
      {stage1_28[201]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[51],stage2_29[61],stage2_28[62],stage2_27[82]}
   );
   gpc615_5 gpc6467 (
      {stage1_27[201], stage1_27[202], stage1_27[203], stage1_27[204], stage1_27[205]},
      {stage1_28[202]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[52],stage2_29[62],stage2_28[63],stage2_27[83]}
   );
   gpc615_5 gpc6468 (
      {stage1_27[206], stage1_27[207], stage1_27[208], stage1_27[209], stage1_27[210]},
      {stage1_28[203]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[53],stage2_29[63],stage2_28[64],stage2_27[84]}
   );
   gpc606_5 gpc6469 (
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[24],stage2_30[54],stage2_29[64],stage2_28[65]}
   );
   gpc606_5 gpc6470 (
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[25],stage2_30[55],stage2_29[65],stage2_28[66]}
   );
   gpc606_5 gpc6471 (
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[26],stage2_30[56],stage2_29[66],stage2_28[67]}
   );
   gpc606_5 gpc6472 (
      {stage1_28[222], stage1_28[223], stage1_28[224], stage1_28[225], stage1_28[226], stage1_28[227]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[27],stage2_30[57],stage2_29[67],stage2_28[68]}
   );
   gpc606_5 gpc6473 (
      {stage1_28[228], stage1_28[229], stage1_28[230], stage1_28[231], stage1_28[232], stage1_28[233]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[28],stage2_30[58],stage2_29[68],stage2_28[69]}
   );
   gpc606_5 gpc6474 (
      {stage1_28[234], stage1_28[235], stage1_28[236], stage1_28[237], stage1_28[238], stage1_28[239]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[29],stage2_30[59],stage2_29[69],stage2_28[70]}
   );
   gpc606_5 gpc6475 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[6],stage2_31[30],stage2_30[60],stage2_29[70]}
   );
   gpc606_5 gpc6476 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[7],stage2_31[31],stage2_30[61],stage2_29[71]}
   );
   gpc606_5 gpc6477 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[8],stage2_31[32],stage2_30[62],stage2_29[72]}
   );
   gpc606_5 gpc6478 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[9],stage2_31[33],stage2_30[63],stage2_29[73]}
   );
   gpc606_5 gpc6479 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[10],stage2_31[34],stage2_30[64],stage2_29[74]}
   );
   gpc606_5 gpc6480 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[11],stage2_31[35],stage2_30[65],stage2_29[75]}
   );
   gpc606_5 gpc6481 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[12],stage2_31[36],stage2_30[66],stage2_29[76]}
   );
   gpc2135_5 gpc6482 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40]},
      {stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_32[0]},
      {stage1_33[0], stage1_33[1]},
      {stage2_34[0],stage2_33[7],stage2_32[13],stage2_31[37],stage2_30[67]}
   );
   gpc207_4 gpc6483 (
      {stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[1], stage1_32[2]},
      {stage2_33[8],stage2_32[14],stage2_31[38],stage2_30[68]}
   );
   gpc207_4 gpc6484 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_32[3], stage1_32[4]},
      {stage2_33[9],stage2_32[15],stage2_31[39],stage2_30[69]}
   );
   gpc207_4 gpc6485 (
      {stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_32[5], stage1_32[6]},
      {stage2_33[10],stage2_32[16],stage2_31[40],stage2_30[70]}
   );
   gpc207_4 gpc6486 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66], stage1_30[67], stage1_30[68]},
      {stage1_32[7], stage1_32[8]},
      {stage2_33[11],stage2_32[17],stage2_31[41],stage2_30[71]}
   );
   gpc207_4 gpc6487 (
      {stage1_30[69], stage1_30[70], stage1_30[71], stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75]},
      {stage1_32[9], stage1_32[10]},
      {stage2_33[12],stage2_32[18],stage2_31[42],stage2_30[72]}
   );
   gpc606_5 gpc6488 (
      {stage1_30[76], stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16]},
      {stage2_34[1],stage2_33[13],stage2_32[19],stage2_31[43],stage2_30[73]}
   );
   gpc606_5 gpc6489 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87]},
      {stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22]},
      {stage2_34[2],stage2_33[14],stage2_32[20],stage2_31[44],stage2_30[74]}
   );
   gpc606_5 gpc6490 (
      {stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93]},
      {stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28]},
      {stage2_34[3],stage2_33[15],stage2_32[21],stage2_31[45],stage2_30[75]}
   );
   gpc606_5 gpc6491 (
      {stage1_30[94], stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34]},
      {stage2_34[4],stage2_33[16],stage2_32[22],stage2_31[46],stage2_30[76]}
   );
   gpc606_5 gpc6492 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105]},
      {stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40]},
      {stage2_34[5],stage2_33[17],stage2_32[23],stage2_31[47],stage2_30[77]}
   );
   gpc606_5 gpc6493 (
      {stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111]},
      {stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46]},
      {stage2_34[6],stage2_33[18],stage2_32[24],stage2_31[48],stage2_30[78]}
   );
   gpc606_5 gpc6494 (
      {stage1_30[112], stage1_30[113], stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117]},
      {stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52]},
      {stage2_34[7],stage2_33[19],stage2_32[25],stage2_31[49],stage2_30[79]}
   );
   gpc606_5 gpc6495 (
      {stage1_30[118], stage1_30[119], stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123]},
      {stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58]},
      {stage2_34[8],stage2_33[20],stage2_32[26],stage2_31[50],stage2_30[80]}
   );
   gpc606_5 gpc6496 (
      {stage1_30[124], stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64]},
      {stage2_34[9],stage2_33[21],stage2_32[27],stage2_31[51],stage2_30[81]}
   );
   gpc606_5 gpc6497 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135]},
      {stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70]},
      {stage2_34[10],stage2_33[22],stage2_32[28],stage2_31[52],stage2_30[82]}
   );
   gpc606_5 gpc6498 (
      {stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141]},
      {stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76]},
      {stage2_34[11],stage2_33[23],stage2_32[29],stage2_31[53],stage2_30[83]}
   );
   gpc606_5 gpc6499 (
      {stage1_30[142], stage1_30[143], stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147]},
      {stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82]},
      {stage2_34[12],stage2_33[24],stage2_32[30],stage2_31[54],stage2_30[84]}
   );
   gpc606_5 gpc6500 (
      {stage1_30[148], stage1_30[149], stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153]},
      {stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88]},
      {stage2_34[13],stage2_33[25],stage2_32[31],stage2_31[55],stage2_30[85]}
   );
   gpc606_5 gpc6501 (
      {stage1_30[154], stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94]},
      {stage2_34[14],stage2_33[26],stage2_32[32],stage2_31[56],stage2_30[86]}
   );
   gpc606_5 gpc6502 (
      {stage1_30[160], stage1_30[161], stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165]},
      {stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100]},
      {stage2_34[15],stage2_33[27],stage2_32[33],stage2_31[57],stage2_30[87]}
   );
   gpc606_5 gpc6503 (
      {stage1_30[166], stage1_30[167], stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171]},
      {stage1_32[101], stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106]},
      {stage2_34[16],stage2_33[28],stage2_32[34],stage2_31[58],stage2_30[88]}
   );
   gpc606_5 gpc6504 (
      {stage1_30[172], stage1_30[173], stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177]},
      {stage1_32[107], stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112]},
      {stage2_34[17],stage2_33[29],stage2_32[35],stage2_31[59],stage2_30[89]}
   );
   gpc606_5 gpc6505 (
      {stage1_30[178], stage1_30[179], stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183]},
      {stage1_32[113], stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118]},
      {stage2_34[18],stage2_33[30],stage2_32[36],stage2_31[60],stage2_30[90]}
   );
   gpc606_5 gpc6506 (
      {stage1_30[184], stage1_30[185], stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189]},
      {stage1_32[119], stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124]},
      {stage2_34[19],stage2_33[31],stage2_32[37],stage2_31[61],stage2_30[91]}
   );
   gpc606_5 gpc6507 (
      {stage1_30[190], stage1_30[191], stage1_30[192], stage1_30[193], stage1_30[194], stage1_30[195]},
      {stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130]},
      {stage2_34[20],stage2_33[32],stage2_32[38],stage2_31[62],stage2_30[92]}
   );
   gpc606_5 gpc6508 (
      {stage1_30[196], stage1_30[197], stage1_30[198], stage1_30[199], stage1_30[200], stage1_30[201]},
      {stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136]},
      {stage2_34[21],stage2_33[33],stage2_32[39],stage2_31[63],stage2_30[93]}
   );
   gpc606_5 gpc6509 (
      {stage1_30[202], stage1_30[203], stage1_30[204], stage1_30[205], stage1_30[206], stage1_30[207]},
      {stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140], stage1_32[141], stage1_32[142]},
      {stage2_34[22],stage2_33[34],stage2_32[40],stage2_31[64],stage2_30[94]}
   );
   gpc606_5 gpc6510 (
      {stage1_30[208], stage1_30[209], stage1_30[210], stage1_30[211], stage1_30[212], stage1_30[213]},
      {stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146], stage1_32[147], stage1_32[148]},
      {stage2_34[23],stage2_33[35],stage2_32[41],stage2_31[65],stage2_30[95]}
   );
   gpc606_5 gpc6511 (
      {stage1_30[214], stage1_30[215], stage1_30[216], stage1_30[217], stage1_30[218], stage1_30[219]},
      {stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152], stage1_32[153], stage1_32[154]},
      {stage2_34[24],stage2_33[36],stage2_32[42],stage2_31[66],stage2_30[96]}
   );
   gpc606_5 gpc6512 (
      {stage1_30[220], stage1_30[221], stage1_30[222], stage1_30[223], stage1_30[224], stage1_30[225]},
      {stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158], stage1_32[159], stage1_32[160]},
      {stage2_34[25],stage2_33[37],stage2_32[43],stage2_31[67],stage2_30[97]}
   );
   gpc606_5 gpc6513 (
      {stage1_30[226], stage1_30[227], stage1_30[228], stage1_30[229], stage1_30[230], stage1_30[231]},
      {stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164], stage1_32[165], stage1_32[166]},
      {stage2_34[26],stage2_33[38],stage2_32[44],stage2_31[68],stage2_30[98]}
   );
   gpc615_5 gpc6514 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49]},
      {stage1_32[167]},
      {stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6], stage1_33[7]},
      {stage2_35[0],stage2_34[27],stage2_33[39],stage2_32[45],stage2_31[69]}
   );
   gpc615_5 gpc6515 (
      {stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54]},
      {stage1_32[168]},
      {stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12], stage1_33[13]},
      {stage2_35[1],stage2_34[28],stage2_33[40],stage2_32[46],stage2_31[70]}
   );
   gpc615_5 gpc6516 (
      {stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage1_32[169]},
      {stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18], stage1_33[19]},
      {stage2_35[2],stage2_34[29],stage2_33[41],stage2_32[47],stage2_31[71]}
   );
   gpc615_5 gpc6517 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64]},
      {stage1_32[170]},
      {stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24], stage1_33[25]},
      {stage2_35[3],stage2_34[30],stage2_33[42],stage2_32[48],stage2_31[72]}
   );
   gpc615_5 gpc6518 (
      {stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69]},
      {stage1_32[171]},
      {stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30], stage1_33[31]},
      {stage2_35[4],stage2_34[31],stage2_33[43],stage2_32[49],stage2_31[73]}
   );
   gpc615_5 gpc6519 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[172]},
      {stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36], stage1_33[37]},
      {stage2_35[5],stage2_34[32],stage2_33[44],stage2_32[50],stage2_31[74]}
   );
   gpc615_5 gpc6520 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79]},
      {stage1_32[173]},
      {stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42], stage1_33[43]},
      {stage2_35[6],stage2_34[33],stage2_33[45],stage2_32[51],stage2_31[75]}
   );
   gpc615_5 gpc6521 (
      {stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84]},
      {stage1_32[174]},
      {stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48], stage1_33[49]},
      {stage2_35[7],stage2_34[34],stage2_33[46],stage2_32[52],stage2_31[76]}
   );
   gpc615_5 gpc6522 (
      {stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_32[175]},
      {stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54], stage1_33[55]},
      {stage2_35[8],stage2_34[35],stage2_33[47],stage2_32[53],stage2_31[77]}
   );
   gpc615_5 gpc6523 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94]},
      {stage1_32[176]},
      {stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60], stage1_33[61]},
      {stage2_35[9],stage2_34[36],stage2_33[48],stage2_32[54],stage2_31[78]}
   );
   gpc615_5 gpc6524 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99]},
      {stage1_32[177]},
      {stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66], stage1_33[67]},
      {stage2_35[10],stage2_34[37],stage2_33[49],stage2_32[55],stage2_31[79]}
   );
   gpc615_5 gpc6525 (
      {stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_32[178]},
      {stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72], stage1_33[73]},
      {stage2_35[11],stage2_34[38],stage2_33[50],stage2_32[56],stage2_31[80]}
   );
   gpc615_5 gpc6526 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[179]},
      {stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78], stage1_33[79]},
      {stage2_35[12],stage2_34[39],stage2_33[51],stage2_32[57],stage2_31[81]}
   );
   gpc615_5 gpc6527 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[180]},
      {stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84], stage1_33[85]},
      {stage2_35[13],stage2_34[40],stage2_33[52],stage2_32[58],stage2_31[82]}
   );
   gpc615_5 gpc6528 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[181]},
      {stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90], stage1_33[91]},
      {stage2_35[14],stage2_34[41],stage2_33[53],stage2_32[59],stage2_31[83]}
   );
   gpc615_5 gpc6529 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[182]},
      {stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96], stage1_33[97]},
      {stage2_35[15],stage2_34[42],stage2_33[54],stage2_32[60],stage2_31[84]}
   );
   gpc615_5 gpc6530 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[183]},
      {stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102], stage1_33[103]},
      {stage2_35[16],stage2_34[43],stage2_33[55],stage2_32[61],stage2_31[85]}
   );
   gpc615_5 gpc6531 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[184]},
      {stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108], stage1_33[109]},
      {stage2_35[17],stage2_34[44],stage2_33[56],stage2_32[62],stage2_31[86]}
   );
   gpc615_5 gpc6532 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[185]},
      {stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114], stage1_33[115]},
      {stage2_35[18],stage2_34[45],stage2_33[57],stage2_32[63],stage2_31[87]}
   );
   gpc615_5 gpc6533 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[186]},
      {stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120], stage1_33[121]},
      {stage2_35[19],stage2_34[46],stage2_33[58],stage2_32[64],stage2_31[88]}
   );
   gpc615_5 gpc6534 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[187]},
      {stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126], stage1_33[127]},
      {stage2_35[20],stage2_34[47],stage2_33[59],stage2_32[65],stage2_31[89]}
   );
   gpc615_5 gpc6535 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[188]},
      {stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132], stage1_33[133]},
      {stage2_35[21],stage2_34[48],stage2_33[60],stage2_32[66],stage2_31[90]}
   );
   gpc615_5 gpc6536 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[189]},
      {stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138], stage1_33[139]},
      {stage2_35[22],stage2_34[49],stage2_33[61],stage2_32[67],stage2_31[91]}
   );
   gpc615_5 gpc6537 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[190]},
      {stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144], stage1_33[145]},
      {stage2_35[23],stage2_34[50],stage2_33[62],stage2_32[68],stage2_31[92]}
   );
   gpc615_5 gpc6538 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[191]},
      {stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150], stage1_33[151]},
      {stage2_35[24],stage2_34[51],stage2_33[63],stage2_32[69],stage2_31[93]}
   );
   gpc615_5 gpc6539 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[192]},
      {stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156], stage1_33[157]},
      {stage2_35[25],stage2_34[52],stage2_33[64],stage2_32[70],stage2_31[94]}
   );
   gpc615_5 gpc6540 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[193]},
      {stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162], stage1_33[163]},
      {stage2_35[26],stage2_34[53],stage2_33[65],stage2_32[71],stage2_31[95]}
   );
   gpc606_5 gpc6541 (
      {stage1_32[194], stage1_32[195], stage1_32[196], stage1_32[197], stage1_32[198], stage1_32[199]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[27],stage2_34[54],stage2_33[66],stage2_32[72]}
   );
   gpc606_5 gpc6542 (
      {stage1_32[200], stage1_32[201], stage1_32[202], stage1_32[203], stage1_32[204], stage1_32[205]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[28],stage2_34[55],stage2_33[67],stage2_32[73]}
   );
   gpc606_5 gpc6543 (
      {stage1_32[206], stage1_32[207], stage1_32[208], stage1_32[209], stage1_32[210], stage1_32[211]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[29],stage2_34[56],stage2_33[68],stage2_32[74]}
   );
   gpc606_5 gpc6544 (
      {stage1_32[212], stage1_32[213], stage1_32[214], stage1_32[215], stage1_32[216], stage1_32[217]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[30],stage2_34[57],stage2_33[69],stage2_32[75]}
   );
   gpc606_5 gpc6545 (
      {stage1_32[218], stage1_32[219], stage1_32[220], stage1_32[221], stage1_32[222], stage1_32[223]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[31],stage2_34[58],stage2_33[70],stage2_32[76]}
   );
   gpc606_5 gpc6546 (
      {stage1_32[224], stage1_32[225], stage1_32[226], stage1_32[227], stage1_32[228], stage1_32[229]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[32],stage2_34[59],stage2_33[71],stage2_32[77]}
   );
   gpc606_5 gpc6547 (
      {stage1_32[230], stage1_32[231], stage1_32[232], stage1_32[233], stage1_32[234], stage1_32[235]},
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage2_36[6],stage2_35[33],stage2_34[60],stage2_33[72],stage2_32[78]}
   );
   gpc606_5 gpc6548 (
      {stage1_32[236], stage1_32[237], stage1_32[238], stage1_32[239], stage1_32[240], stage1_32[241]},
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage2_36[7],stage2_35[34],stage2_34[61],stage2_33[73],stage2_32[79]}
   );
   gpc606_5 gpc6549 (
      {stage1_32[242], stage1_32[243], stage1_32[244], stage1_32[245], stage1_32[246], stage1_32[247]},
      {stage1_34[48], stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53]},
      {stage2_36[8],stage2_35[35],stage2_34[62],stage2_33[74],stage2_32[80]}
   );
   gpc606_5 gpc6550 (
      {stage1_32[248], stage1_32[249], stage1_32[250], stage1_32[251], stage1_32[252], stage1_32[253]},
      {stage1_34[54], stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59]},
      {stage2_36[9],stage2_35[36],stage2_34[63],stage2_33[75],stage2_32[81]}
   );
   gpc606_5 gpc6551 (
      {stage1_32[254], stage1_32[255], stage1_32[256], stage1_32[257], stage1_32[258], stage1_32[259]},
      {stage1_34[60], stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage2_36[10],stage2_35[37],stage2_34[64],stage2_33[76],stage2_32[82]}
   );
   gpc606_5 gpc6552 (
      {stage1_32[260], stage1_32[261], stage1_32[262], stage1_32[263], stage1_32[264], stage1_32[265]},
      {stage1_34[66], stage1_34[67], stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71]},
      {stage2_36[11],stage2_35[38],stage2_34[65],stage2_33[77],stage2_32[83]}
   );
   gpc606_5 gpc6553 (
      {stage1_32[266], stage1_32[267], stage1_32[268], stage1_32[269], stage1_32[270], stage1_32[271]},
      {stage1_34[72], stage1_34[73], stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77]},
      {stage2_36[12],stage2_35[39],stage2_34[66],stage2_33[78],stage2_32[84]}
   );
   gpc606_5 gpc6554 (
      {stage1_32[272], stage1_32[273], stage1_32[274], stage1_32[275], stage1_32[276], stage1_32[277]},
      {stage1_34[78], stage1_34[79], stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83]},
      {stage2_36[13],stage2_35[40],stage2_34[67],stage2_33[79],stage2_32[85]}
   );
   gpc606_5 gpc6555 (
      {stage1_32[278], stage1_32[279], stage1_32[280], stage1_32[281], stage1_32[282], stage1_32[283]},
      {stage1_34[84], stage1_34[85], stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89]},
      {stage2_36[14],stage2_35[41],stage2_34[68],stage2_33[80],stage2_32[86]}
   );
   gpc606_5 gpc6556 (
      {stage1_32[284], stage1_32[285], stage1_32[286], stage1_32[287], stage1_32[288], stage1_32[289]},
      {stage1_34[90], stage1_34[91], stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95]},
      {stage2_36[15],stage2_35[42],stage2_34[69],stage2_33[81],stage2_32[87]}
   );
   gpc606_5 gpc6557 (
      {stage1_32[290], stage1_32[291], stage1_32[292], stage1_32[293], stage1_32[294], stage1_32[295]},
      {stage1_34[96], stage1_34[97], stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101]},
      {stage2_36[16],stage2_35[43],stage2_34[70],stage2_33[82],stage2_32[88]}
   );
   gpc606_5 gpc6558 (
      {stage1_32[296], stage1_32[297], stage1_32[298], stage1_32[299], stage1_32[300], stage1_32[301]},
      {stage1_34[102], stage1_34[103], stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107]},
      {stage2_36[17],stage2_35[44],stage2_34[71],stage2_33[83],stage2_32[89]}
   );
   gpc606_5 gpc6559 (
      {stage1_32[302], stage1_32[303], stage1_32[304], stage1_32[305], stage1_32[306], stage1_32[307]},
      {stage1_34[108], stage1_34[109], stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113]},
      {stage2_36[18],stage2_35[45],stage2_34[72],stage2_33[84],stage2_32[90]}
   );
   gpc606_5 gpc6560 (
      {stage1_32[308], stage1_32[309], stage1_32[310], stage1_32[311], stage1_32[312], stage1_32[313]},
      {stage1_34[114], stage1_34[115], stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119]},
      {stage2_36[19],stage2_35[46],stage2_34[73],stage2_33[85],stage2_32[91]}
   );
   gpc606_5 gpc6561 (
      {stage1_32[314], stage1_32[315], stage1_32[316], stage1_32[317], stage1_32[318], stage1_32[319]},
      {stage1_34[120], stage1_34[121], stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125]},
      {stage2_36[20],stage2_35[47],stage2_34[74],stage2_33[86],stage2_32[92]}
   );
   gpc606_5 gpc6562 (
      {stage1_32[320], stage1_32[321], stage1_32[322], stage1_32[323], stage1_32[324], stage1_32[325]},
      {stage1_34[126], stage1_34[127], stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131]},
      {stage2_36[21],stage2_35[48],stage2_34[75],stage2_33[87],stage2_32[93]}
   );
   gpc606_5 gpc6563 (
      {stage1_32[326], stage1_32[327], stage1_32[328], stage1_32[329], stage1_32[330], stage1_32[331]},
      {stage1_34[132], stage1_34[133], stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137]},
      {stage2_36[22],stage2_35[49],stage2_34[76],stage2_33[88],stage2_32[94]}
   );
   gpc606_5 gpc6564 (
      {stage1_32[332], stage1_32[333], stage1_32[334], stage1_32[335], stage1_32[336], stage1_32[337]},
      {stage1_34[138], stage1_34[139], stage1_34[140], stage1_34[141], stage1_34[142], stage1_34[143]},
      {stage2_36[23],stage2_35[50],stage2_34[77],stage2_33[89],stage2_32[95]}
   );
   gpc606_5 gpc6565 (
      {stage1_32[338], stage1_32[339], stage1_32[340], stage1_32[341], stage1_32[342], stage1_32[343]},
      {stage1_34[144], stage1_34[145], stage1_34[146], stage1_34[147], stage1_34[148], stage1_34[149]},
      {stage2_36[24],stage2_35[51],stage2_34[78],stage2_33[90],stage2_32[96]}
   );
   gpc606_5 gpc6566 (
      {stage1_32[344], stage1_32[345], stage1_32[346], stage1_32[347], stage1_32[348], stage1_32[349]},
      {stage1_34[150], stage1_34[151], stage1_34[152], stage1_34[153], stage1_34[154], stage1_34[155]},
      {stage2_36[25],stage2_35[52],stage2_34[79],stage2_33[91],stage2_32[97]}
   );
   gpc606_5 gpc6567 (
      {stage1_32[350], stage1_32[351], stage1_32[352], stage1_32[353], stage1_32[354], stage1_32[355]},
      {stage1_34[156], stage1_34[157], stage1_34[158], stage1_34[159], stage1_34[160], stage1_34[161]},
      {stage2_36[26],stage2_35[53],stage2_34[80],stage2_33[92],stage2_32[98]}
   );
   gpc606_5 gpc6568 (
      {stage1_32[356], stage1_32[357], stage1_32[358], stage1_32[359], stage1_32[360], stage1_32[361]},
      {stage1_34[162], stage1_34[163], stage1_34[164], stage1_34[165], stage1_34[166], stage1_34[167]},
      {stage2_36[27],stage2_35[54],stage2_34[81],stage2_33[93],stage2_32[99]}
   );
   gpc606_5 gpc6569 (
      {stage1_32[362], stage1_32[363], stage1_32[364], stage1_32[365], stage1_32[366], stage1_32[367]},
      {stage1_34[168], stage1_34[169], stage1_34[170], stage1_34[171], stage1_34[172], stage1_34[173]},
      {stage2_36[28],stage2_35[55],stage2_34[82],stage2_33[94],stage2_32[100]}
   );
   gpc606_5 gpc6570 (
      {stage1_32[368], stage1_32[369], stage1_32[370], stage1_32[371], stage1_32[372], stage1_32[373]},
      {stage1_34[174], stage1_34[175], stage1_34[176], stage1_34[177], stage1_34[178], stage1_34[179]},
      {stage2_36[29],stage2_35[56],stage2_34[83],stage2_33[95],stage2_32[101]}
   );
   gpc606_5 gpc6571 (
      {stage1_32[374], stage1_32[375], stage1_32[376], stage1_32[377], stage1_32[378], stage1_32[379]},
      {stage1_34[180], stage1_34[181], stage1_34[182], stage1_34[183], stage1_34[184], stage1_34[185]},
      {stage2_36[30],stage2_35[57],stage2_34[84],stage2_33[96],stage2_32[102]}
   );
   gpc606_5 gpc6572 (
      {stage1_32[380], stage1_32[381], stage1_32[382], stage1_32[383], stage1_32[384], stage1_32[385]},
      {stage1_34[186], stage1_34[187], stage1_34[188], stage1_34[189], stage1_34[190], stage1_34[191]},
      {stage2_36[31],stage2_35[58],stage2_34[85],stage2_33[97],stage2_32[103]}
   );
   gpc606_5 gpc6573 (
      {stage1_32[386], stage1_32[387], stage1_32[388], stage1_32[389], stage1_32[390], stage1_32[391]},
      {stage1_34[192], stage1_34[193], stage1_34[194], stage1_34[195], stage1_34[196], stage1_34[197]},
      {stage2_36[32],stage2_35[59],stage2_34[86],stage2_33[98],stage2_32[104]}
   );
   gpc606_5 gpc6574 (
      {stage1_32[392], stage1_32[393], stage1_32[394], stage1_32[395], stage1_32[396], stage1_32[397]},
      {stage1_34[198], stage1_34[199], stage1_34[200], stage1_34[201], stage1_34[202], stage1_34[203]},
      {stage2_36[33],stage2_35[60],stage2_34[87],stage2_33[99],stage2_32[105]}
   );
   gpc606_5 gpc6575 (
      {stage1_32[398], stage1_32[399], stage1_32[400], stage1_32[401], stage1_32[402], stage1_32[403]},
      {stage1_34[204], stage1_34[205], stage1_34[206], stage1_34[207], stage1_34[208], stage1_34[209]},
      {stage2_36[34],stage2_35[61],stage2_34[88],stage2_33[100],stage2_32[106]}
   );
   gpc606_5 gpc6576 (
      {stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168], stage1_33[169]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[35],stage2_35[62],stage2_34[89],stage2_33[101]}
   );
   gpc606_5 gpc6577 (
      {stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174], stage1_33[175]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[36],stage2_35[63],stage2_34[90],stage2_33[102]}
   );
   gpc606_5 gpc6578 (
      {stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180], stage1_33[181]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[37],stage2_35[64],stage2_34[91],stage2_33[103]}
   );
   gpc606_5 gpc6579 (
      {stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186], stage1_33[187]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[38],stage2_35[65],stage2_34[92],stage2_33[104]}
   );
   gpc606_5 gpc6580 (
      {stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192], stage1_33[193]},
      {stage1_35[24], stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29]},
      {stage2_37[4],stage2_36[39],stage2_35[66],stage2_34[93],stage2_33[105]}
   );
   gpc606_5 gpc6581 (
      {stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198], stage1_33[199]},
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage2_37[5],stage2_36[40],stage2_35[67],stage2_34[94],stage2_33[106]}
   );
   gpc615_5 gpc6582 (
      {stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage1_34[210]},
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage2_37[6],stage2_36[41],stage2_35[68],stage2_34[95],stage2_33[107]}
   );
   gpc615_5 gpc6583 (
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209]},
      {stage1_34[211]},
      {stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage2_37[7],stage2_36[42],stage2_35[69],stage2_34[96],stage2_33[108]}
   );
   gpc606_5 gpc6584 (
      {stage1_34[212], stage1_34[213], stage1_34[214], stage1_34[215], stage1_34[216], stage1_34[217]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[8],stage2_36[43],stage2_35[70],stage2_34[97]}
   );
   gpc606_5 gpc6585 (
      {stage1_34[218], stage1_34[219], stage1_34[220], stage1_34[221], stage1_34[222], stage1_34[223]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[9],stage2_36[44],stage2_35[71],stage2_34[98]}
   );
   gpc606_5 gpc6586 (
      {stage1_34[224], stage1_34[225], stage1_34[226], stage1_34[227], stage1_34[228], stage1_34[229]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[10],stage2_36[45],stage2_35[72],stage2_34[99]}
   );
   gpc606_5 gpc6587 (
      {stage1_34[230], stage1_34[231], stage1_34[232], stage1_34[233], stage1_34[234], stage1_34[235]},
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23]},
      {stage2_38[3],stage2_37[11],stage2_36[46],stage2_35[73],stage2_34[100]}
   );
   gpc606_5 gpc6588 (
      {stage1_34[236], stage1_34[237], stage1_34[238], stage1_34[239], stage1_34[240], stage1_34[241]},
      {stage1_36[24], stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29]},
      {stage2_38[4],stage2_37[12],stage2_36[47],stage2_35[74],stage2_34[101]}
   );
   gpc615_5 gpc6589 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[30]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[5],stage2_37[13],stage2_36[48],stage2_35[75]}
   );
   gpc615_5 gpc6590 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[31]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[6],stage2_37[14],stage2_36[49],stage2_35[76]}
   );
   gpc615_5 gpc6591 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[32]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[7],stage2_37[15],stage2_36[50],stage2_35[77]}
   );
   gpc615_5 gpc6592 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[33]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[8],stage2_37[16],stage2_36[51],stage2_35[78]}
   );
   gpc615_5 gpc6593 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[34]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[9],stage2_37[17],stage2_36[52],stage2_35[79]}
   );
   gpc615_5 gpc6594 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[35]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[10],stage2_37[18],stage2_36[53],stage2_35[80]}
   );
   gpc615_5 gpc6595 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[36]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[11],stage2_37[19],stage2_36[54],stage2_35[81]}
   );
   gpc615_5 gpc6596 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[37]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[12],stage2_37[20],stage2_36[55],stage2_35[82]}
   );
   gpc615_5 gpc6597 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[38]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[13],stage2_37[21],stage2_36[56],stage2_35[83]}
   );
   gpc615_5 gpc6598 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[39]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[14],stage2_37[22],stage2_36[57],stage2_35[84]}
   );
   gpc615_5 gpc6599 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[40]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[15],stage2_37[23],stage2_36[58],stage2_35[85]}
   );
   gpc615_5 gpc6600 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[41]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[16],stage2_37[24],stage2_36[59],stage2_35[86]}
   );
   gpc615_5 gpc6601 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[42]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[17],stage2_37[25],stage2_36[60],stage2_35[87]}
   );
   gpc615_5 gpc6602 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[43]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[18],stage2_37[26],stage2_36[61],stage2_35[88]}
   );
   gpc615_5 gpc6603 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[44]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[19],stage2_37[27],stage2_36[62],stage2_35[89]}
   );
   gpc615_5 gpc6604 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[45]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[20],stage2_37[28],stage2_36[63],stage2_35[90]}
   );
   gpc615_5 gpc6605 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[46]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[21],stage2_37[29],stage2_36[64],stage2_35[91]}
   );
   gpc615_5 gpc6606 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[47]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[22],stage2_37[30],stage2_36[65],stage2_35[92]}
   );
   gpc615_5 gpc6607 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[48]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[23],stage2_37[31],stage2_36[66],stage2_35[93]}
   );
   gpc615_5 gpc6608 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[49]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[24],stage2_37[32],stage2_36[67],stage2_35[94]}
   );
   gpc615_5 gpc6609 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[50]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[25],stage2_37[33],stage2_36[68],stage2_35[95]}
   );
   gpc615_5 gpc6610 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[51]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[26],stage2_37[34],stage2_36[69],stage2_35[96]}
   );
   gpc615_5 gpc6611 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[52]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[27],stage2_37[35],stage2_36[70],stage2_35[97]}
   );
   gpc615_5 gpc6612 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[53]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[28],stage2_37[36],stage2_36[71],stage2_35[98]}
   );
   gpc615_5 gpc6613 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[54]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[29],stage2_37[37],stage2_36[72],stage2_35[99]}
   );
   gpc1163_5 gpc6614 (
      {stage1_36[55], stage1_36[56], stage1_36[57]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage1_38[0]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[25],stage2_38[30],stage2_37[38],stage2_36[73]}
   );
   gpc606_5 gpc6615 (
      {stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61], stage1_36[62], stage1_36[63]},
      {stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6]},
      {stage2_40[1],stage2_39[26],stage2_38[31],stage2_37[39],stage2_36[74]}
   );
   gpc606_5 gpc6616 (
      {stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67], stage1_36[68], stage1_36[69]},
      {stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12]},
      {stage2_40[2],stage2_39[27],stage2_38[32],stage2_37[40],stage2_36[75]}
   );
   gpc606_5 gpc6617 (
      {stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73], stage1_36[74], stage1_36[75]},
      {stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18]},
      {stage2_40[3],stage2_39[28],stage2_38[33],stage2_37[41],stage2_36[76]}
   );
   gpc606_5 gpc6618 (
      {stage1_36[76], stage1_36[77], stage1_36[78], stage1_36[79], stage1_36[80], stage1_36[81]},
      {stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24]},
      {stage2_40[4],stage2_39[29],stage2_38[34],stage2_37[42],stage2_36[77]}
   );
   gpc606_5 gpc6619 (
      {stage1_36[82], stage1_36[83], stage1_36[84], stage1_36[85], stage1_36[86], stage1_36[87]},
      {stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30]},
      {stage2_40[5],stage2_39[30],stage2_38[35],stage2_37[43],stage2_36[78]}
   );
   gpc606_5 gpc6620 (
      {stage1_36[88], stage1_36[89], stage1_36[90], stage1_36[91], stage1_36[92], stage1_36[93]},
      {stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36]},
      {stage2_40[6],stage2_39[31],stage2_38[36],stage2_37[44],stage2_36[79]}
   );
   gpc606_5 gpc6621 (
      {stage1_36[94], stage1_36[95], stage1_36[96], stage1_36[97], stage1_36[98], stage1_36[99]},
      {stage1_38[37], stage1_38[38], stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42]},
      {stage2_40[7],stage2_39[32],stage2_38[37],stage2_37[45],stage2_36[80]}
   );
   gpc606_5 gpc6622 (
      {stage1_36[100], stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105]},
      {stage1_38[43], stage1_38[44], stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48]},
      {stage2_40[8],stage2_39[33],stage2_38[38],stage2_37[46],stage2_36[81]}
   );
   gpc606_5 gpc6623 (
      {stage1_36[106], stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111]},
      {stage1_38[49], stage1_38[50], stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54]},
      {stage2_40[9],stage2_39[34],stage2_38[39],stage2_37[47],stage2_36[82]}
   );
   gpc606_5 gpc6624 (
      {stage1_36[112], stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117]},
      {stage1_38[55], stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage2_40[10],stage2_39[35],stage2_38[40],stage2_37[48],stage2_36[83]}
   );
   gpc606_5 gpc6625 (
      {stage1_36[118], stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123]},
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65], stage1_38[66]},
      {stage2_40[11],stage2_39[36],stage2_38[41],stage2_37[49],stage2_36[84]}
   );
   gpc606_5 gpc6626 (
      {stage1_36[124], stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129]},
      {stage1_38[67], stage1_38[68], stage1_38[69], stage1_38[70], stage1_38[71], stage1_38[72]},
      {stage2_40[12],stage2_39[37],stage2_38[42],stage2_37[50],stage2_36[85]}
   );
   gpc606_5 gpc6627 (
      {stage1_36[130], stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135]},
      {stage1_38[73], stage1_38[74], stage1_38[75], stage1_38[76], stage1_38[77], stage1_38[78]},
      {stage2_40[13],stage2_39[38],stage2_38[43],stage2_37[51],stage2_36[86]}
   );
   gpc606_5 gpc6628 (
      {stage1_36[136], stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141]},
      {stage1_38[79], stage1_38[80], stage1_38[81], stage1_38[82], stage1_38[83], stage1_38[84]},
      {stage2_40[14],stage2_39[39],stage2_38[44],stage2_37[52],stage2_36[87]}
   );
   gpc606_5 gpc6629 (
      {stage1_36[142], stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147]},
      {stage1_38[85], stage1_38[86], stage1_38[87], stage1_38[88], stage1_38[89], stage1_38[90]},
      {stage2_40[15],stage2_39[40],stage2_38[45],stage2_37[53],stage2_36[88]}
   );
   gpc606_5 gpc6630 (
      {stage1_36[148], stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153]},
      {stage1_38[91], stage1_38[92], stage1_38[93], stage1_38[94], stage1_38[95], stage1_38[96]},
      {stage2_40[16],stage2_39[41],stage2_38[46],stage2_37[54],stage2_36[89]}
   );
   gpc606_5 gpc6631 (
      {stage1_36[154], stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159]},
      {stage1_38[97], stage1_38[98], stage1_38[99], stage1_38[100], stage1_38[101], stage1_38[102]},
      {stage2_40[17],stage2_39[42],stage2_38[47],stage2_37[55],stage2_36[90]}
   );
   gpc606_5 gpc6632 (
      {stage1_36[160], stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165]},
      {stage1_38[103], stage1_38[104], stage1_38[105], stage1_38[106], stage1_38[107], stage1_38[108]},
      {stage2_40[18],stage2_39[43],stage2_38[48],stage2_37[56],stage2_36[91]}
   );
   gpc606_5 gpc6633 (
      {stage1_36[166], stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171]},
      {stage1_38[109], stage1_38[110], stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114]},
      {stage2_40[19],stage2_39[44],stage2_38[49],stage2_37[57],stage2_36[92]}
   );
   gpc606_5 gpc6634 (
      {stage1_36[172], stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177]},
      {stage1_38[115], stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage2_40[20],stage2_39[45],stage2_38[50],stage2_37[58],stage2_36[93]}
   );
   gpc606_5 gpc6635 (
      {stage1_36[178], stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183]},
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125], stage1_38[126]},
      {stage2_40[21],stage2_39[46],stage2_38[51],stage2_37[59],stage2_36[94]}
   );
   gpc606_5 gpc6636 (
      {stage1_36[184], stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189]},
      {stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130], stage1_38[131], stage1_38[132]},
      {stage2_40[22],stage2_39[47],stage2_38[52],stage2_37[60],stage2_36[95]}
   );
   gpc606_5 gpc6637 (
      {stage1_36[190], stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195]},
      {stage1_38[133], stage1_38[134], stage1_38[135], stage1_38[136], stage1_38[137], stage1_38[138]},
      {stage2_40[23],stage2_39[48],stage2_38[53],stage2_37[61],stage2_36[96]}
   );
   gpc606_5 gpc6638 (
      {stage1_36[196], stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201]},
      {stage1_38[139], stage1_38[140], stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144]},
      {stage2_40[24],stage2_39[49],stage2_38[54],stage2_37[62],stage2_36[97]}
   );
   gpc606_5 gpc6639 (
      {stage1_36[202], stage1_36[203], stage1_36[204], stage1_36[205], stage1_36[206], stage1_36[207]},
      {stage1_38[145], stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage2_40[25],stage2_39[50],stage2_38[55],stage2_37[63],stage2_36[98]}
   );
   gpc606_5 gpc6640 (
      {stage1_36[208], stage1_36[209], stage1_36[210], stage1_36[211], stage1_36[212], stage1_36[213]},
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155], stage1_38[156]},
      {stage2_40[26],stage2_39[51],stage2_38[56],stage2_37[64],stage2_36[99]}
   );
   gpc606_5 gpc6641 (
      {stage1_36[214], stage1_36[215], stage1_36[216], stage1_36[217], stage1_36[218], stage1_36[219]},
      {stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160], stage1_38[161], stage1_38[162]},
      {stage2_40[27],stage2_39[52],stage2_38[57],stage2_37[65],stage2_36[100]}
   );
   gpc606_5 gpc6642 (
      {stage1_36[220], stage1_36[221], stage1_36[222], stage1_36[223], stage1_36[224], stage1_36[225]},
      {stage1_38[163], stage1_38[164], stage1_38[165], stage1_38[166], stage1_38[167], stage1_38[168]},
      {stage2_40[28],stage2_39[53],stage2_38[58],stage2_37[66],stage2_36[101]}
   );
   gpc606_5 gpc6643 (
      {stage1_36[226], stage1_36[227], stage1_36[228], stage1_36[229], stage1_36[230], stage1_36[231]},
      {stage1_38[169], stage1_38[170], stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174]},
      {stage2_40[29],stage2_39[54],stage2_38[59],stage2_37[67],stage2_36[102]}
   );
   gpc606_5 gpc6644 (
      {stage1_36[232], stage1_36[233], stage1_36[234], stage1_36[235], stage1_36[236], stage1_36[237]},
      {stage1_38[175], stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage2_40[30],stage2_39[55],stage2_38[60],stage2_37[68],stage2_36[103]}
   );
   gpc606_5 gpc6645 (
      {stage1_36[238], stage1_36[239], stage1_36[240], stage1_36[241], stage1_36[242], stage1_36[243]},
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185], stage1_38[186]},
      {stage2_40[31],stage2_39[56],stage2_38[61],stage2_37[69],stage2_36[104]}
   );
   gpc606_5 gpc6646 (
      {stage1_36[244], stage1_36[245], stage1_36[246], stage1_36[247], stage1_36[248], stage1_36[249]},
      {stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190], stage1_38[191], stage1_38[192]},
      {stage2_40[32],stage2_39[57],stage2_38[62],stage2_37[70],stage2_36[105]}
   );
   gpc606_5 gpc6647 (
      {stage1_36[250], stage1_36[251], stage1_36[252], stage1_36[253], stage1_36[254], stage1_36[255]},
      {stage1_38[193], stage1_38[194], stage1_38[195], stage1_38[196], stage1_38[197], stage1_38[198]},
      {stage2_40[33],stage2_39[58],stage2_38[63],stage2_37[71],stage2_36[106]}
   );
   gpc606_5 gpc6648 (
      {stage1_36[256], stage1_36[257], stage1_36[258], stage1_36[259], stage1_36[260], stage1_36[261]},
      {stage1_38[199], stage1_38[200], stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204]},
      {stage2_40[34],stage2_39[59],stage2_38[64],stage2_37[72],stage2_36[107]}
   );
   gpc606_5 gpc6649 (
      {stage1_36[262], stage1_36[263], stage1_36[264], stage1_36[265], stage1_36[266], stage1_36[267]},
      {stage1_38[205], stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage2_40[35],stage2_39[60],stage2_38[65],stage2_37[73],stage2_36[108]}
   );
   gpc606_5 gpc6650 (
      {stage1_36[268], stage1_36[269], stage1_36[270], stage1_36[271], stage1_36[272], stage1_36[273]},
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215], stage1_38[216]},
      {stage2_40[36],stage2_39[61],stage2_38[66],stage2_37[74],stage2_36[109]}
   );
   gpc606_5 gpc6651 (
      {stage1_36[274], stage1_36[275], stage1_36[276], stage1_36[277], stage1_36[278], stage1_36[279]},
      {stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220], stage1_38[221], stage1_38[222]},
      {stage2_40[37],stage2_39[62],stage2_38[67],stage2_37[75],stage2_36[110]}
   );
   gpc606_5 gpc6652 (
      {stage1_36[280], stage1_36[281], stage1_36[282], stage1_36[283], stage1_36[284], stage1_36[285]},
      {stage1_38[223], stage1_38[224], stage1_38[225], stage1_38[226], stage1_38[227], stage1_38[228]},
      {stage2_40[38],stage2_39[63],stage2_38[68],stage2_37[76],stage2_36[111]}
   );
   gpc606_5 gpc6653 (
      {stage1_36[286], stage1_36[287], stage1_36[288], stage1_36[289], stage1_36[290], stage1_36[291]},
      {stage1_38[229], stage1_38[230], stage1_38[231], stage1_38[232], stage1_38[233], stage1_38[234]},
      {stage2_40[39],stage2_39[64],stage2_38[69],stage2_37[77],stage2_36[112]}
   );
   gpc606_5 gpc6654 (
      {stage1_36[292], stage1_36[293], stage1_36[294], stage1_36[295], stage1_36[296], stage1_36[297]},
      {stage1_38[235], stage1_38[236], stage1_38[237], stage1_38[238], stage1_38[239], stage1_38[240]},
      {stage2_40[40],stage2_39[65],stage2_38[70],stage2_37[78],stage2_36[113]}
   );
   gpc606_5 gpc6655 (
      {stage1_36[298], stage1_36[299], stage1_36[300], stage1_36[301], stage1_36[302], stage1_36[303]},
      {stage1_38[241], stage1_38[242], stage1_38[243], stage1_38[244], stage1_38[245], stage1_38[246]},
      {stage2_40[41],stage2_39[66],stage2_38[71],stage2_37[79],stage2_36[114]}
   );
   gpc606_5 gpc6656 (
      {stage1_36[304], stage1_36[305], stage1_36[306], stage1_36[307], stage1_36[308], stage1_36[309]},
      {stage1_38[247], stage1_38[248], stage1_38[249], stage1_38[250], stage1_38[251], stage1_38[252]},
      {stage2_40[42],stage2_39[67],stage2_38[72],stage2_37[80],stage2_36[115]}
   );
   gpc606_5 gpc6657 (
      {stage1_36[310], stage1_36[311], stage1_36[312], stage1_36[313], stage1_36[314], stage1_36[315]},
      {stage1_38[253], stage1_38[254], stage1_38[255], stage1_38[256], stage1_38[257], stage1_38[258]},
      {stage2_40[43],stage2_39[68],stage2_38[73],stage2_37[81],stage2_36[116]}
   );
   gpc615_5 gpc6658 (
      {stage1_36[316], stage1_36[317], stage1_36[318], stage1_36[319], stage1_36[320]},
      {stage1_37[156]},
      {stage1_38[259], stage1_38[260], stage1_38[261], stage1_38[262], stage1_38[263], stage1_38[264]},
      {stage2_40[44],stage2_39[69],stage2_38[74],stage2_37[82],stage2_36[117]}
   );
   gpc615_5 gpc6659 (
      {stage1_36[321], stage1_36[322], stage1_36[323], stage1_36[324], stage1_36[325]},
      {stage1_37[157]},
      {stage1_38[265], stage1_38[266], stage1_38[267], stage1_38[268], stage1_38[269], stage1_38[270]},
      {stage2_40[45],stage2_39[70],stage2_38[75],stage2_37[83],stage2_36[118]}
   );
   gpc615_5 gpc6660 (
      {stage1_36[326], stage1_36[327], stage1_36[328], stage1_36[329], stage1_36[330]},
      {stage1_37[158]},
      {stage1_38[271], stage1_38[272], stage1_38[273], stage1_38[274], stage1_38[275], stage1_38[276]},
      {stage2_40[46],stage2_39[71],stage2_38[76],stage2_37[84],stage2_36[119]}
   );
   gpc606_5 gpc6661 (
      {stage1_37[159], stage1_37[160], stage1_37[161], stage1_37[162], stage1_37[163], stage1_37[164]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[47],stage2_39[72],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc6662 (
      {stage1_37[165], stage1_37[166], stage1_37[167], stage1_37[168], stage1_37[169], stage1_37[170]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[48],stage2_39[73],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc6663 (
      {stage1_37[171], stage1_37[172], stage1_37[173], stage1_37[174], stage1_37[175], stage1_37[176]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[49],stage2_39[74],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc6664 (
      {stage1_37[177], stage1_37[178], stage1_37[179], stage1_37[180], stage1_37[181], stage1_37[182]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[50],stage2_39[75],stage2_38[80],stage2_37[88]}
   );
   gpc606_5 gpc6665 (
      {stage1_37[183], stage1_37[184], stage1_37[185], stage1_37[186], stage1_37[187], stage1_37[188]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[51],stage2_39[76],stage2_38[81],stage2_37[89]}
   );
   gpc606_5 gpc6666 (
      {stage1_37[189], stage1_37[190], stage1_37[191], stage1_37[192], stage1_37[193], stage1_37[194]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[52],stage2_39[77],stage2_38[82],stage2_37[90]}
   );
   gpc606_5 gpc6667 (
      {stage1_37[195], stage1_37[196], stage1_37[197], stage1_37[198], stage1_37[199], stage1_37[200]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[53],stage2_39[78],stage2_38[83],stage2_37[91]}
   );
   gpc606_5 gpc6668 (
      {stage1_37[201], stage1_37[202], stage1_37[203], stage1_37[204], stage1_37[205], stage1_37[206]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[54],stage2_39[79],stage2_38[84],stage2_37[92]}
   );
   gpc606_5 gpc6669 (
      {stage1_37[207], stage1_37[208], stage1_37[209], stage1_37[210], stage1_37[211], stage1_37[212]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[55],stage2_39[80],stage2_38[85],stage2_37[93]}
   );
   gpc606_5 gpc6670 (
      {stage1_37[213], stage1_37[214], stage1_37[215], stage1_37[216], stage1_37[217], stage1_37[218]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[56],stage2_39[81],stage2_38[86],stage2_37[94]}
   );
   gpc606_5 gpc6671 (
      {stage1_37[219], stage1_37[220], stage1_37[221], stage1_37[222], stage1_37[223], stage1_37[224]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[57],stage2_39[82],stage2_38[87],stage2_37[95]}
   );
   gpc606_5 gpc6672 (
      {stage1_37[225], stage1_37[226], stage1_37[227], stage1_37[228], stage1_37[229], stage1_37[230]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[58],stage2_39[83],stage2_38[88],stage2_37[96]}
   );
   gpc606_5 gpc6673 (
      {stage1_37[231], stage1_37[232], stage1_37[233], stage1_37[234], stage1_37[235], stage1_37[236]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[59],stage2_39[84],stage2_38[89],stage2_37[97]}
   );
   gpc606_5 gpc6674 (
      {stage1_37[237], stage1_37[238], stage1_37[239], stage1_37[240], stage1_37[241], stage1_37[242]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[60],stage2_39[85],stage2_38[90],stage2_37[98]}
   );
   gpc606_5 gpc6675 (
      {stage1_37[243], stage1_37[244], stage1_37[245], stage1_37[246], stage1_37[247], stage1_37[248]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[61],stage2_39[86],stage2_38[91],stage2_37[99]}
   );
   gpc606_5 gpc6676 (
      {stage1_37[249], stage1_37[250], stage1_37[251], stage1_37[252], stage1_37[253], stage1_37[254]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[62],stage2_39[87],stage2_38[92],stage2_37[100]}
   );
   gpc606_5 gpc6677 (
      {stage1_37[255], stage1_37[256], stage1_37[257], stage1_37[258], stage1_37[259], stage1_37[260]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[63],stage2_39[88],stage2_38[93],stage2_37[101]}
   );
   gpc606_5 gpc6678 (
      {stage1_37[261], stage1_37[262], stage1_37[263], stage1_37[264], stage1_37[265], stage1_37[266]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[64],stage2_39[89],stage2_38[94],stage2_37[102]}
   );
   gpc606_5 gpc6679 (
      {stage1_37[267], stage1_37[268], stage1_37[269], stage1_37[270], stage1_37[271], stage1_37[272]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[65],stage2_39[90],stage2_38[95],stage2_37[103]}
   );
   gpc606_5 gpc6680 (
      {stage1_37[273], stage1_37[274], stage1_37[275], stage1_37[276], stage1_37[277], stage1_37[278]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[66],stage2_39[91],stage2_38[96],stage2_37[104]}
   );
   gpc606_5 gpc6681 (
      {stage1_37[279], stage1_37[280], stage1_37[281], stage1_37[282], stage1_37[283], stage1_37[284]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[67],stage2_39[92],stage2_38[97],stage2_37[105]}
   );
   gpc606_5 gpc6682 (
      {stage1_37[285], stage1_37[286], stage1_37[287], stage1_37[288], stage1_37[289], stage1_37[290]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[68],stage2_39[93],stage2_38[98],stage2_37[106]}
   );
   gpc606_5 gpc6683 (
      {stage1_37[291], stage1_37[292], stage1_37[293], stage1_37[294], stage1_37[295], stage1_37[296]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[69],stage2_39[94],stage2_38[99],stage2_37[107]}
   );
   gpc606_5 gpc6684 (
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[0],stage2_41[23],stage2_40[70],stage2_39[95]}
   );
   gpc606_5 gpc6685 (
      {stage1_39[145], stage1_39[146], stage1_39[147], stage1_39[148], stage1_39[149], stage1_39[150]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage2_43[1],stage2_42[1],stage2_41[24],stage2_40[71],stage2_39[96]}
   );
   gpc606_5 gpc6686 (
      {stage1_39[151], stage1_39[152], stage1_39[153], stage1_39[154], stage1_39[155], stage1_39[156]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage2_43[2],stage2_42[2],stage2_41[25],stage2_40[72],stage2_39[97]}
   );
   gpc606_5 gpc6687 (
      {stage1_39[157], stage1_39[158], stage1_39[159], stage1_39[160], stage1_39[161], stage1_39[162]},
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage2_43[3],stage2_42[3],stage2_41[26],stage2_40[73],stage2_39[98]}
   );
   gpc606_5 gpc6688 (
      {stage1_39[163], stage1_39[164], stage1_39[165], stage1_39[166], stage1_39[167], stage1_39[168]},
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage2_43[4],stage2_42[4],stage2_41[27],stage2_40[74],stage2_39[99]}
   );
   gpc615_5 gpc6689 (
      {stage1_39[169], stage1_39[170], stage1_39[171], stage1_39[172], stage1_39[173]},
      {stage1_40[0]},
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage2_43[5],stage2_42[5],stage2_41[28],stage2_40[75],stage2_39[100]}
   );
   gpc615_5 gpc6690 (
      {stage1_39[174], stage1_39[175], stage1_39[176], stage1_39[177], stage1_39[178]},
      {stage1_40[1]},
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage2_43[6],stage2_42[6],stage2_41[29],stage2_40[76],stage2_39[101]}
   );
   gpc615_5 gpc6691 (
      {stage1_39[179], stage1_39[180], stage1_39[181], stage1_39[182], stage1_39[183]},
      {stage1_40[2]},
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage2_43[7],stage2_42[7],stage2_41[30],stage2_40[77],stage2_39[102]}
   );
   gpc615_5 gpc6692 (
      {stage1_39[184], stage1_39[185], stage1_39[186], stage1_39[187], stage1_39[188]},
      {stage1_40[3]},
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52], stage1_41[53]},
      {stage2_43[8],stage2_42[8],stage2_41[31],stage2_40[78],stage2_39[103]}
   );
   gpc615_5 gpc6693 (
      {stage1_39[189], stage1_39[190], stage1_39[191], stage1_39[192], stage1_39[193]},
      {stage1_40[4]},
      {stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57], stage1_41[58], stage1_41[59]},
      {stage2_43[9],stage2_42[9],stage2_41[32],stage2_40[79],stage2_39[104]}
   );
   gpc606_5 gpc6694 (
      {stage1_40[5], stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[10],stage2_42[10],stage2_41[33],stage2_40[80]}
   );
   gpc606_5 gpc6695 (
      {stage1_40[11], stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[11],stage2_42[11],stage2_41[34],stage2_40[81]}
   );
   gpc606_5 gpc6696 (
      {stage1_40[17], stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[12],stage2_42[12],stage2_41[35],stage2_40[82]}
   );
   gpc606_5 gpc6697 (
      {stage1_40[23], stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[13],stage2_42[13],stage2_41[36],stage2_40[83]}
   );
   gpc606_5 gpc6698 (
      {stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[14],stage2_42[14],stage2_41[37],stage2_40[84]}
   );
   gpc606_5 gpc6699 (
      {stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[15],stage2_42[15],stage2_41[38],stage2_40[85]}
   );
   gpc606_5 gpc6700 (
      {stage1_40[41], stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[16],stage2_42[16],stage2_41[39],stage2_40[86]}
   );
   gpc606_5 gpc6701 (
      {stage1_40[47], stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[17],stage2_42[17],stage2_41[40],stage2_40[87]}
   );
   gpc606_5 gpc6702 (
      {stage1_40[53], stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[18],stage2_42[18],stage2_41[41],stage2_40[88]}
   );
   gpc606_5 gpc6703 (
      {stage1_40[59], stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[19],stage2_42[19],stage2_41[42],stage2_40[89]}
   );
   gpc606_5 gpc6704 (
      {stage1_40[65], stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[20],stage2_42[20],stage2_41[43],stage2_40[90]}
   );
   gpc606_5 gpc6705 (
      {stage1_40[71], stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[21],stage2_42[21],stage2_41[44],stage2_40[91]}
   );
   gpc606_5 gpc6706 (
      {stage1_40[77], stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[22],stage2_42[22],stage2_41[45],stage2_40[92]}
   );
   gpc606_5 gpc6707 (
      {stage1_40[83], stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[23],stage2_42[23],stage2_41[46],stage2_40[93]}
   );
   gpc606_5 gpc6708 (
      {stage1_40[89], stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[24],stage2_42[24],stage2_41[47],stage2_40[94]}
   );
   gpc606_5 gpc6709 (
      {stage1_40[95], stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[25],stage2_42[25],stage2_41[48],stage2_40[95]}
   );
   gpc606_5 gpc6710 (
      {stage1_40[101], stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[26],stage2_42[26],stage2_41[49],stage2_40[96]}
   );
   gpc606_5 gpc6711 (
      {stage1_40[107], stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[27],stage2_42[27],stage2_41[50],stage2_40[97]}
   );
   gpc606_5 gpc6712 (
      {stage1_40[113], stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[28],stage2_42[28],stage2_41[51],stage2_40[98]}
   );
   gpc606_5 gpc6713 (
      {stage1_40[119], stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[29],stage2_42[29],stage2_41[52],stage2_40[99]}
   );
   gpc606_5 gpc6714 (
      {stage1_40[125], stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[30],stage2_42[30],stage2_41[53],stage2_40[100]}
   );
   gpc606_5 gpc6715 (
      {stage1_40[131], stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[31],stage2_42[31],stage2_41[54],stage2_40[101]}
   );
   gpc606_5 gpc6716 (
      {stage1_40[137], stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[32],stage2_42[32],stage2_41[55],stage2_40[102]}
   );
   gpc606_5 gpc6717 (
      {stage1_40[143], stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148]},
      {stage1_42[138], stage1_42[139], stage1_42[140], stage1_42[141], stage1_42[142], stage1_42[143]},
      {stage2_44[23],stage2_43[33],stage2_42[33],stage2_41[56],stage2_40[103]}
   );
   gpc606_5 gpc6718 (
      {stage1_40[149], stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154]},
      {stage1_42[144], stage1_42[145], stage1_42[146], stage1_42[147], stage1_42[148], stage1_42[149]},
      {stage2_44[24],stage2_43[34],stage2_42[34],stage2_41[57],stage2_40[104]}
   );
   gpc606_5 gpc6719 (
      {stage1_40[155], stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160]},
      {stage1_42[150], stage1_42[151], stage1_42[152], stage1_42[153], stage1_42[154], stage1_42[155]},
      {stage2_44[25],stage2_43[35],stage2_42[35],stage2_41[58],stage2_40[105]}
   );
   gpc606_5 gpc6720 (
      {stage1_40[161], stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166]},
      {stage1_42[156], stage1_42[157], stage1_42[158], stage1_42[159], stage1_42[160], stage1_42[161]},
      {stage2_44[26],stage2_43[36],stage2_42[36],stage2_41[59],stage2_40[106]}
   );
   gpc606_5 gpc6721 (
      {stage1_40[167], stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172]},
      {stage1_42[162], stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage2_44[27],stage2_43[37],stage2_42[37],stage2_41[60],stage2_40[107]}
   );
   gpc606_5 gpc6722 (
      {stage1_40[173], stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178]},
      {stage1_42[168], stage1_42[169], stage1_42[170], stage1_42[171], stage1_42[172], stage1_42[173]},
      {stage2_44[28],stage2_43[38],stage2_42[38],stage2_41[61],stage2_40[108]}
   );
   gpc606_5 gpc6723 (
      {stage1_40[179], stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184]},
      {stage1_42[174], stage1_42[175], stage1_42[176], stage1_42[177], stage1_42[178], stage1_42[179]},
      {stage2_44[29],stage2_43[39],stage2_42[39],stage2_41[62],stage2_40[109]}
   );
   gpc606_5 gpc6724 (
      {stage1_40[185], stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190]},
      {stage1_42[180], stage1_42[181], stage1_42[182], stage1_42[183], stage1_42[184], stage1_42[185]},
      {stage2_44[30],stage2_43[40],stage2_42[40],stage2_41[63],stage2_40[110]}
   );
   gpc606_5 gpc6725 (
      {stage1_40[191], stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196]},
      {stage1_42[186], stage1_42[187], stage1_42[188], stage1_42[189], stage1_42[190], stage1_42[191]},
      {stage2_44[31],stage2_43[41],stage2_42[41],stage2_41[64],stage2_40[111]}
   );
   gpc606_5 gpc6726 (
      {stage1_40[197], stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202]},
      {stage1_42[192], stage1_42[193], stage1_42[194], stage1_42[195], stage1_42[196], stage1_42[197]},
      {stage2_44[32],stage2_43[42],stage2_42[42],stage2_41[65],stage2_40[112]}
   );
   gpc606_5 gpc6727 (
      {stage1_41[60], stage1_41[61], stage1_41[62], stage1_41[63], stage1_41[64], stage1_41[65]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[33],stage2_43[43],stage2_42[43],stage2_41[66]}
   );
   gpc606_5 gpc6728 (
      {stage1_41[66], stage1_41[67], stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[34],stage2_43[44],stage2_42[44],stage2_41[67]}
   );
   gpc606_5 gpc6729 (
      {stage1_41[72], stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[35],stage2_43[45],stage2_42[45],stage2_41[68]}
   );
   gpc606_5 gpc6730 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82], stage1_41[83]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[36],stage2_43[46],stage2_42[46],stage2_41[69]}
   );
   gpc606_5 gpc6731 (
      {stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87], stage1_41[88], stage1_41[89]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[37],stage2_43[47],stage2_42[47],stage2_41[70]}
   );
   gpc606_5 gpc6732 (
      {stage1_41[90], stage1_41[91], stage1_41[92], stage1_41[93], stage1_41[94], stage1_41[95]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[38],stage2_43[48],stage2_42[48],stage2_41[71]}
   );
   gpc606_5 gpc6733 (
      {stage1_41[96], stage1_41[97], stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[39],stage2_43[49],stage2_42[49],stage2_41[72]}
   );
   gpc606_5 gpc6734 (
      {stage1_41[102], stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[40],stage2_43[50],stage2_42[50],stage2_41[73]}
   );
   gpc606_5 gpc6735 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112], stage1_41[113]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[41],stage2_43[51],stage2_42[51],stage2_41[74]}
   );
   gpc606_5 gpc6736 (
      {stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117], stage1_41[118], stage1_41[119]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[42],stage2_43[52],stage2_42[52],stage2_41[75]}
   );
   gpc606_5 gpc6737 (
      {stage1_41[120], stage1_41[121], stage1_41[122], stage1_41[123], stage1_41[124], stage1_41[125]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[43],stage2_43[53],stage2_42[53],stage2_41[76]}
   );
   gpc606_5 gpc6738 (
      {stage1_41[126], stage1_41[127], stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[44],stage2_43[54],stage2_42[54],stage2_41[77]}
   );
   gpc606_5 gpc6739 (
      {stage1_41[132], stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[45],stage2_43[55],stage2_42[55],stage2_41[78]}
   );
   gpc606_5 gpc6740 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142], stage1_41[143]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[46],stage2_43[56],stage2_42[56],stage2_41[79]}
   );
   gpc606_5 gpc6741 (
      {stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147], stage1_41[148], stage1_41[149]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[47],stage2_43[57],stage2_42[57],stage2_41[80]}
   );
   gpc606_5 gpc6742 (
      {stage1_41[150], stage1_41[151], stage1_41[152], stage1_41[153], stage1_41[154], stage1_41[155]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[48],stage2_43[58],stage2_42[58],stage2_41[81]}
   );
   gpc606_5 gpc6743 (
      {stage1_41[156], stage1_41[157], stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[49],stage2_43[59],stage2_42[59],stage2_41[82]}
   );
   gpc606_5 gpc6744 (
      {stage1_41[162], stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[50],stage2_43[60],stage2_42[60],stage2_41[83]}
   );
   gpc606_5 gpc6745 (
      {stage1_41[168], stage1_41[169], stage1_41[170], stage1_41[171], stage1_41[172], stage1_41[173]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[51],stage2_43[61],stage2_42[61],stage2_41[84]}
   );
   gpc606_5 gpc6746 (
      {stage1_41[174], stage1_41[175], stage1_41[176], stage1_41[177], stage1_41[178], stage1_41[179]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[52],stage2_43[62],stage2_42[62],stage2_41[85]}
   );
   gpc606_5 gpc6747 (
      {stage1_41[180], stage1_41[181], stage1_41[182], stage1_41[183], stage1_41[184], stage1_41[185]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[53],stage2_43[63],stage2_42[63],stage2_41[86]}
   );
   gpc606_5 gpc6748 (
      {stage1_41[186], stage1_41[187], stage1_41[188], stage1_41[189], stage1_41[190], stage1_41[191]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[54],stage2_43[64],stage2_42[64],stage2_41[87]}
   );
   gpc606_5 gpc6749 (
      {stage1_41[192], stage1_41[193], stage1_41[194], stage1_41[195], stage1_41[196], stage1_41[197]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[55],stage2_43[65],stage2_42[65],stage2_41[88]}
   );
   gpc606_5 gpc6750 (
      {stage1_41[198], stage1_41[199], stage1_41[200], stage1_41[201], stage1_41[202], stage1_41[203]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[56],stage2_43[66],stage2_42[66],stage2_41[89]}
   );
   gpc606_5 gpc6751 (
      {stage1_41[204], stage1_41[205], stage1_41[206], stage1_41[207], stage1_41[208], stage1_41[209]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[57],stage2_43[67],stage2_42[67],stage2_41[90]}
   );
   gpc606_5 gpc6752 (
      {stage1_41[210], stage1_41[211], stage1_41[212], stage1_41[213], stage1_41[214], stage1_41[215]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[58],stage2_43[68],stage2_42[68],stage2_41[91]}
   );
   gpc606_5 gpc6753 (
      {stage1_41[216], stage1_41[217], stage1_41[218], stage1_41[219], stage1_41[220], stage1_41[221]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[59],stage2_43[69],stage2_42[69],stage2_41[92]}
   );
   gpc606_5 gpc6754 (
      {stage1_41[222], stage1_41[223], stage1_41[224], stage1_41[225], stage1_41[226], stage1_41[227]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[60],stage2_43[70],stage2_42[70],stage2_41[93]}
   );
   gpc606_5 gpc6755 (
      {stage1_41[228], stage1_41[229], stage1_41[230], stage1_41[231], stage1_41[232], stage1_41[233]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[61],stage2_43[71],stage2_42[71],stage2_41[94]}
   );
   gpc606_5 gpc6756 (
      {stage1_41[234], stage1_41[235], stage1_41[236], stage1_41[237], stage1_41[238], stage1_41[239]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[62],stage2_43[72],stage2_42[72],stage2_41[95]}
   );
   gpc606_5 gpc6757 (
      {stage1_41[240], stage1_41[241], stage1_41[242], stage1_41[243], stage1_41[244], stage1_41[245]},
      {stage1_43[180], stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage2_45[30],stage2_44[63],stage2_43[73],stage2_42[73],stage2_41[96]}
   );
   gpc606_5 gpc6758 (
      {stage1_41[246], stage1_41[247], stage1_41[248], stage1_41[249], stage1_41[250], stage1_41[251]},
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190], stage1_43[191]},
      {stage2_45[31],stage2_44[64],stage2_43[74],stage2_42[74],stage2_41[97]}
   );
   gpc615_5 gpc6759 (
      {stage1_42[198], stage1_42[199], stage1_42[200], stage1_42[201], stage1_42[202]},
      {stage1_43[192]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[32],stage2_44[65],stage2_43[75],stage2_42[75]}
   );
   gpc615_5 gpc6760 (
      {stage1_42[203], stage1_42[204], stage1_42[205], stage1_42[206], stage1_42[207]},
      {stage1_43[193]},
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage2_46[1],stage2_45[33],stage2_44[66],stage2_43[76],stage2_42[76]}
   );
   gpc615_5 gpc6761 (
      {stage1_42[208], stage1_42[209], stage1_42[210], stage1_42[211], stage1_42[212]},
      {stage1_43[194]},
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage2_46[2],stage2_45[34],stage2_44[67],stage2_43[77],stage2_42[77]}
   );
   gpc615_5 gpc6762 (
      {stage1_42[213], stage1_42[214], stage1_42[215], stage1_42[216], stage1_42[217]},
      {stage1_43[195]},
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage2_46[3],stage2_45[35],stage2_44[68],stage2_43[78],stage2_42[78]}
   );
   gpc615_5 gpc6763 (
      {stage1_42[218], stage1_42[219], stage1_42[220], stage1_42[221], stage1_42[222]},
      {stage1_43[196]},
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage2_46[4],stage2_45[36],stage2_44[69],stage2_43[79],stage2_42[79]}
   );
   gpc615_5 gpc6764 (
      {stage1_42[223], stage1_42[224], stage1_42[225], stage1_42[226], stage1_42[227]},
      {stage1_43[197]},
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage2_46[5],stage2_45[37],stage2_44[70],stage2_43[80],stage2_42[80]}
   );
   gpc1415_5 gpc6765 (
      {stage1_43[198], stage1_43[199], stage1_43[200], stage1_43[201], stage1_43[202]},
      {stage1_44[36]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3]},
      {stage1_46[0]},
      {stage2_47[0],stage2_46[6],stage2_45[38],stage2_44[71],stage2_43[81]}
   );
   gpc1415_5 gpc6766 (
      {stage1_43[203], stage1_43[204], stage1_43[205], stage1_43[206], stage1_43[207]},
      {stage1_44[37]},
      {stage1_45[4], stage1_45[5], stage1_45[6], stage1_45[7]},
      {stage1_46[1]},
      {stage2_47[1],stage2_46[7],stage2_45[39],stage2_44[72],stage2_43[82]}
   );
   gpc1415_5 gpc6767 (
      {stage1_43[208], stage1_43[209], stage1_43[210], stage1_43[211], stage1_43[212]},
      {stage1_44[38]},
      {stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage1_46[2]},
      {stage2_47[2],stage2_46[8],stage2_45[40],stage2_44[73],stage2_43[83]}
   );
   gpc1415_5 gpc6768 (
      {stage1_43[213], stage1_43[214], stage1_43[215], stage1_43[216], stage1_43[217]},
      {stage1_44[39]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15]},
      {stage1_46[3]},
      {stage2_47[3],stage2_46[9],stage2_45[41],stage2_44[74],stage2_43[84]}
   );
   gpc606_5 gpc6769 (
      {stage1_44[40], stage1_44[41], stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45]},
      {stage1_46[4], stage1_46[5], stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9]},
      {stage2_48[0],stage2_47[4],stage2_46[10],stage2_45[42],stage2_44[75]}
   );
   gpc606_5 gpc6770 (
      {stage1_44[46], stage1_44[47], stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51]},
      {stage1_46[10], stage1_46[11], stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15]},
      {stage2_48[1],stage2_47[5],stage2_46[11],stage2_45[43],stage2_44[76]}
   );
   gpc606_5 gpc6771 (
      {stage1_44[52], stage1_44[53], stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57]},
      {stage1_46[16], stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage2_48[2],stage2_47[6],stage2_46[12],stage2_45[44],stage2_44[77]}
   );
   gpc606_5 gpc6772 (
      {stage1_44[58], stage1_44[59], stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63]},
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27]},
      {stage2_48[3],stage2_47[7],stage2_46[13],stage2_45[45],stage2_44[78]}
   );
   gpc606_5 gpc6773 (
      {stage1_44[64], stage1_44[65], stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69]},
      {stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33]},
      {stage2_48[4],stage2_47[8],stage2_46[14],stage2_45[46],stage2_44[79]}
   );
   gpc606_5 gpc6774 (
      {stage1_44[70], stage1_44[71], stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75]},
      {stage1_46[34], stage1_46[35], stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39]},
      {stage2_48[5],stage2_47[9],stage2_46[15],stage2_45[47],stage2_44[80]}
   );
   gpc606_5 gpc6775 (
      {stage1_44[76], stage1_44[77], stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81]},
      {stage1_46[40], stage1_46[41], stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45]},
      {stage2_48[6],stage2_47[10],stage2_46[16],stage2_45[48],stage2_44[81]}
   );
   gpc606_5 gpc6776 (
      {stage1_44[82], stage1_44[83], stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87]},
      {stage1_46[46], stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage2_48[7],stage2_47[11],stage2_46[17],stage2_45[49],stage2_44[82]}
   );
   gpc606_5 gpc6777 (
      {stage1_44[88], stage1_44[89], stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93]},
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57]},
      {stage2_48[8],stage2_47[12],stage2_46[18],stage2_45[50],stage2_44[83]}
   );
   gpc606_5 gpc6778 (
      {stage1_44[94], stage1_44[95], stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99]},
      {stage1_46[58], stage1_46[59], stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63]},
      {stage2_48[9],stage2_47[13],stage2_46[19],stage2_45[51],stage2_44[84]}
   );
   gpc606_5 gpc6779 (
      {stage1_44[100], stage1_44[101], stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105]},
      {stage1_46[64], stage1_46[65], stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69]},
      {stage2_48[10],stage2_47[14],stage2_46[20],stage2_45[52],stage2_44[85]}
   );
   gpc606_5 gpc6780 (
      {stage1_44[106], stage1_44[107], stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111]},
      {stage1_46[70], stage1_46[71], stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75]},
      {stage2_48[11],stage2_47[15],stage2_46[21],stage2_45[53],stage2_44[86]}
   );
   gpc606_5 gpc6781 (
      {stage1_44[112], stage1_44[113], stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117]},
      {stage1_46[76], stage1_46[77], stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81]},
      {stage2_48[12],stage2_47[16],stage2_46[22],stage2_45[54],stage2_44[87]}
   );
   gpc606_5 gpc6782 (
      {stage1_44[118], stage1_44[119], stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123]},
      {stage1_46[82], stage1_46[83], stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87]},
      {stage2_48[13],stage2_47[17],stage2_46[23],stage2_45[55],stage2_44[88]}
   );
   gpc615_5 gpc6783 (
      {stage1_44[124], stage1_44[125], stage1_44[126], stage1_44[127], stage1_44[128]},
      {stage1_45[16]},
      {stage1_46[88], stage1_46[89], stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93]},
      {stage2_48[14],stage2_47[18],stage2_46[24],stage2_45[56],stage2_44[89]}
   );
   gpc615_5 gpc6784 (
      {stage1_44[129], stage1_44[130], stage1_44[131], stage1_44[132], stage1_44[133]},
      {stage1_45[17]},
      {stage1_46[94], stage1_46[95], stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99]},
      {stage2_48[15],stage2_47[19],stage2_46[25],stage2_45[57],stage2_44[90]}
   );
   gpc615_5 gpc6785 (
      {stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137], stage1_44[138]},
      {stage1_45[18]},
      {stage1_46[100], stage1_46[101], stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105]},
      {stage2_48[16],stage2_47[20],stage2_46[26],stage2_45[58],stage2_44[91]}
   );
   gpc615_5 gpc6786 (
      {stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_45[19]},
      {stage1_46[106], stage1_46[107], stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111]},
      {stage2_48[17],stage2_47[21],stage2_46[27],stage2_45[59],stage2_44[92]}
   );
   gpc615_5 gpc6787 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148]},
      {stage1_45[20]},
      {stage1_46[112], stage1_46[113], stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117]},
      {stage2_48[18],stage2_47[22],stage2_46[28],stage2_45[60],stage2_44[93]}
   );
   gpc615_5 gpc6788 (
      {stage1_44[149], stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153]},
      {stage1_45[21]},
      {stage1_46[118], stage1_46[119], stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123]},
      {stage2_48[19],stage2_47[23],stage2_46[29],stage2_45[61],stage2_44[94]}
   );
   gpc615_5 gpc6789 (
      {stage1_44[154], stage1_44[155], stage1_44[156], stage1_44[157], stage1_44[158]},
      {stage1_45[22]},
      {stage1_46[124], stage1_46[125], stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129]},
      {stage2_48[20],stage2_47[24],stage2_46[30],stage2_45[62],stage2_44[95]}
   );
   gpc615_5 gpc6790 (
      {stage1_44[159], stage1_44[160], stage1_44[161], stage1_44[162], stage1_44[163]},
      {stage1_45[23]},
      {stage1_46[130], stage1_46[131], stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135]},
      {stage2_48[21],stage2_47[25],stage2_46[31],stage2_45[63],stage2_44[96]}
   );
   gpc615_5 gpc6791 (
      {stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167], stage1_44[168]},
      {stage1_45[24]},
      {stage1_46[136], stage1_46[137], stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141]},
      {stage2_48[22],stage2_47[26],stage2_46[32],stage2_45[64],stage2_44[97]}
   );
   gpc615_5 gpc6792 (
      {stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_45[25]},
      {stage1_46[142], stage1_46[143], stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147]},
      {stage2_48[23],stage2_47[27],stage2_46[33],stage2_45[65],stage2_44[98]}
   );
   gpc615_5 gpc6793 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178]},
      {stage1_45[26]},
      {stage1_46[148], stage1_46[149], stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153]},
      {stage2_48[24],stage2_47[28],stage2_46[34],stage2_45[66],stage2_44[99]}
   );
   gpc615_5 gpc6794 (
      {stage1_44[179], stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183]},
      {stage1_45[27]},
      {stage1_46[154], stage1_46[155], stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159]},
      {stage2_48[25],stage2_47[29],stage2_46[35],stage2_45[67],stage2_44[100]}
   );
   gpc615_5 gpc6795 (
      {stage1_44[184], stage1_44[185], stage1_44[186], stage1_44[187], stage1_44[188]},
      {stage1_45[28]},
      {stage1_46[160], stage1_46[161], stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165]},
      {stage2_48[26],stage2_47[30],stage2_46[36],stage2_45[68],stage2_44[101]}
   );
   gpc615_5 gpc6796 (
      {stage1_44[189], stage1_44[190], stage1_44[191], stage1_44[192], stage1_44[193]},
      {stage1_45[29]},
      {stage1_46[166], stage1_46[167], stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171]},
      {stage2_48[27],stage2_47[31],stage2_46[37],stage2_45[69],stage2_44[102]}
   );
   gpc615_5 gpc6797 (
      {stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197], stage1_44[198]},
      {stage1_45[30]},
      {stage1_46[172], stage1_46[173], stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177]},
      {stage2_48[28],stage2_47[32],stage2_46[38],stage2_45[70],stage2_44[103]}
   );
   gpc615_5 gpc6798 (
      {stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_45[31]},
      {stage1_46[178], stage1_46[179], stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183]},
      {stage2_48[29],stage2_47[33],stage2_46[39],stage2_45[71],stage2_44[104]}
   );
   gpc615_5 gpc6799 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208]},
      {stage1_45[32]},
      {stage1_46[184], stage1_46[185], stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189]},
      {stage2_48[30],stage2_47[34],stage2_46[40],stage2_45[72],stage2_44[105]}
   );
   gpc615_5 gpc6800 (
      {stage1_44[209], stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213]},
      {stage1_45[33]},
      {stage1_46[190], stage1_46[191], stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195]},
      {stage2_48[31],stage2_47[35],stage2_46[41],stage2_45[73],stage2_44[106]}
   );
   gpc615_5 gpc6801 (
      {stage1_44[214], stage1_44[215], stage1_44[216], stage1_44[217], stage1_44[218]},
      {stage1_45[34]},
      {stage1_46[196], stage1_46[197], stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201]},
      {stage2_48[32],stage2_47[36],stage2_46[42],stage2_45[74],stage2_44[107]}
   );
   gpc615_5 gpc6802 (
      {stage1_44[219], stage1_44[220], stage1_44[221], stage1_44[222], stage1_44[223]},
      {stage1_45[35]},
      {stage1_46[202], stage1_46[203], stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207]},
      {stage2_48[33],stage2_47[37],stage2_46[43],stage2_45[75],stage2_44[108]}
   );
   gpc615_5 gpc6803 (
      {stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227], stage1_44[228]},
      {stage1_45[36]},
      {stage1_46[208], stage1_46[209], stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213]},
      {stage2_48[34],stage2_47[38],stage2_46[44],stage2_45[76],stage2_44[109]}
   );
   gpc615_5 gpc6804 (
      {stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_45[37]},
      {stage1_46[214], stage1_46[215], stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219]},
      {stage2_48[35],stage2_47[39],stage2_46[45],stage2_45[77],stage2_44[110]}
   );
   gpc615_5 gpc6805 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238]},
      {stage1_45[38]},
      {stage1_46[220], stage1_46[221], stage1_46[222], stage1_46[223], stage1_46[224], stage1_46[225]},
      {stage2_48[36],stage2_47[40],stage2_46[46],stage2_45[78],stage2_44[111]}
   );
   gpc615_5 gpc6806 (
      {stage1_44[239], stage1_44[240], stage1_44[241], stage1_44[242], stage1_44[243]},
      {stage1_45[39]},
      {stage1_46[226], stage1_46[227], stage1_46[228], stage1_46[229], stage1_46[230], stage1_46[231]},
      {stage2_48[37],stage2_47[41],stage2_46[47],stage2_45[79],stage2_44[112]}
   );
   gpc606_5 gpc6807 (
      {stage1_45[40], stage1_45[41], stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[38],stage2_47[42],stage2_46[48],stage2_45[80]}
   );
   gpc606_5 gpc6808 (
      {stage1_45[46], stage1_45[47], stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[39],stage2_47[43],stage2_46[49],stage2_45[81]}
   );
   gpc606_5 gpc6809 (
      {stage1_45[52], stage1_45[53], stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[40],stage2_47[44],stage2_46[50],stage2_45[82]}
   );
   gpc606_5 gpc6810 (
      {stage1_45[58], stage1_45[59], stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[41],stage2_47[45],stage2_46[51],stage2_45[83]}
   );
   gpc606_5 gpc6811 (
      {stage1_45[64], stage1_45[65], stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[42],stage2_47[46],stage2_46[52],stage2_45[84]}
   );
   gpc606_5 gpc6812 (
      {stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[43],stage2_47[47],stage2_46[53],stage2_45[85]}
   );
   gpc606_5 gpc6813 (
      {stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[44],stage2_47[48],stage2_46[54],stage2_45[86]}
   );
   gpc606_5 gpc6814 (
      {stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[45],stage2_47[49],stage2_46[55],stage2_45[87]}
   );
   gpc606_5 gpc6815 (
      {stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[46],stage2_47[50],stage2_46[56],stage2_45[88]}
   );
   gpc606_5 gpc6816 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98], stage1_45[99]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[47],stage2_47[51],stage2_46[57],stage2_45[89]}
   );
   gpc606_5 gpc6817 (
      {stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103], stage1_45[104], stage1_45[105]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[48],stage2_47[52],stage2_46[58],stage2_45[90]}
   );
   gpc606_5 gpc6818 (
      {stage1_45[106], stage1_45[107], stage1_45[108], stage1_45[109], stage1_45[110], stage1_45[111]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[49],stage2_47[53],stage2_46[59],stage2_45[91]}
   );
   gpc606_5 gpc6819 (
      {stage1_45[112], stage1_45[113], stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[50],stage2_47[54],stage2_46[60],stage2_45[92]}
   );
   gpc606_5 gpc6820 (
      {stage1_45[118], stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[51],stage2_47[55],stage2_46[61],stage2_45[93]}
   );
   gpc606_5 gpc6821 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128], stage1_45[129]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[52],stage2_47[56],stage2_46[62],stage2_45[94]}
   );
   gpc606_5 gpc6822 (
      {stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133], stage1_45[134], stage1_45[135]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[53],stage2_47[57],stage2_46[63],stage2_45[95]}
   );
   gpc606_5 gpc6823 (
      {stage1_45[136], stage1_45[137], stage1_45[138], stage1_45[139], stage1_45[140], stage1_45[141]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[54],stage2_47[58],stage2_46[64],stage2_45[96]}
   );
   gpc615_5 gpc6824 (
      {stage1_45[142], stage1_45[143], stage1_45[144], stage1_45[145], stage1_45[146]},
      {stage1_46[232]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[55],stage2_47[59],stage2_46[65],stage2_45[97]}
   );
   gpc615_5 gpc6825 (
      {stage1_45[147], stage1_45[148], stage1_45[149], stage1_45[150], stage1_45[151]},
      {stage1_46[233]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[56],stage2_47[60],stage2_46[66],stage2_45[98]}
   );
   gpc615_5 gpc6826 (
      {stage1_45[152], stage1_45[153], stage1_45[154], stage1_45[155], stage1_45[156]},
      {stage1_46[234]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[57],stage2_47[61],stage2_46[67],stage2_45[99]}
   );
   gpc615_5 gpc6827 (
      {stage1_46[235], stage1_46[236], stage1_46[237], stage1_46[238], stage1_46[239]},
      {stage1_47[120]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[20],stage2_48[58],stage2_47[62],stage2_46[68]}
   );
   gpc615_5 gpc6828 (
      {stage1_46[240], stage1_46[241], stage1_46[242], stage1_46[243], stage1_46[244]},
      {stage1_47[121]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[21],stage2_48[59],stage2_47[63],stage2_46[69]}
   );
   gpc615_5 gpc6829 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[122]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[22],stage2_48[60],stage2_47[64],stage2_46[70]}
   );
   gpc615_5 gpc6830 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[123]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[23],stage2_48[61],stage2_47[65],stage2_46[71]}
   );
   gpc615_5 gpc6831 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[124]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[24],stage2_48[62],stage2_47[66],stage2_46[72]}
   );
   gpc615_5 gpc6832 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[125]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[25],stage2_48[63],stage2_47[67],stage2_46[73]}
   );
   gpc615_5 gpc6833 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[126]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[26],stage2_48[64],stage2_47[68],stage2_46[74]}
   );
   gpc615_5 gpc6834 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[127]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[27],stage2_48[65],stage2_47[69],stage2_46[75]}
   );
   gpc615_5 gpc6835 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[128]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[28],stage2_48[66],stage2_47[70],stage2_46[76]}
   );
   gpc615_5 gpc6836 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[129]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[29],stage2_48[67],stage2_47[71],stage2_46[77]}
   );
   gpc615_5 gpc6837 (
      {stage1_47[130], stage1_47[131], stage1_47[132], stage1_47[133], stage1_47[134]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[30],stage2_48[68],stage2_47[72]}
   );
   gpc615_5 gpc6838 (
      {stage1_47[135], stage1_47[136], stage1_47[137], stage1_47[138], stage1_47[139]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[31],stage2_48[69],stage2_47[73]}
   );
   gpc615_5 gpc6839 (
      {stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143], stage1_47[144]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[32],stage2_48[70],stage2_47[74]}
   );
   gpc615_5 gpc6840 (
      {stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[33],stage2_48[71],stage2_47[75]}
   );
   gpc615_5 gpc6841 (
      {stage1_47[150], stage1_47[151], stage1_47[152], stage1_47[153], stage1_47[154]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[34],stage2_48[72],stage2_47[76]}
   );
   gpc615_5 gpc6842 (
      {stage1_47[155], stage1_47[156], stage1_47[157], stage1_47[158], stage1_47[159]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[35],stage2_48[73],stage2_47[77]}
   );
   gpc615_5 gpc6843 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[36],stage2_48[74],stage2_47[78]}
   );
   gpc615_5 gpc6844 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[37],stage2_48[75],stage2_47[79]}
   );
   gpc615_5 gpc6845 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[38],stage2_48[76],stage2_47[80]}
   );
   gpc615_5 gpc6846 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[39],stage2_48[77],stage2_47[81]}
   );
   gpc615_5 gpc6847 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[40],stage2_48[78],stage2_47[82]}
   );
   gpc615_5 gpc6848 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[41],stage2_48[79],stage2_47[83]}
   );
   gpc615_5 gpc6849 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[42],stage2_48[80],stage2_47[84]}
   );
   gpc615_5 gpc6850 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[43],stage2_48[81],stage2_47[85]}
   );
   gpc615_5 gpc6851 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[74]},
      {stage1_49[84], stage1_49[85], stage1_49[86], stage1_49[87], stage1_49[88], stage1_49[89]},
      {stage2_51[14],stage2_50[24],stage2_49[44],stage2_48[82],stage2_47[86]}
   );
   gpc615_5 gpc6852 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[75]},
      {stage1_49[90], stage1_49[91], stage1_49[92], stage1_49[93], stage1_49[94], stage1_49[95]},
      {stage2_51[15],stage2_50[25],stage2_49[45],stage2_48[83],stage2_47[87]}
   );
   gpc615_5 gpc6853 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[76]},
      {stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99], stage1_49[100], stage1_49[101]},
      {stage2_51[16],stage2_50[26],stage2_49[46],stage2_48[84],stage2_47[88]}
   );
   gpc615_5 gpc6854 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[77]},
      {stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105], stage1_49[106], stage1_49[107]},
      {stage2_51[17],stage2_50[27],stage2_49[47],stage2_48[85],stage2_47[89]}
   );
   gpc615_5 gpc6855 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[78]},
      {stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111], stage1_49[112], stage1_49[113]},
      {stage2_51[18],stage2_50[28],stage2_49[48],stage2_48[86],stage2_47[90]}
   );
   gpc615_5 gpc6856 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[79]},
      {stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117], stage1_49[118], stage1_49[119]},
      {stage2_51[19],stage2_50[29],stage2_49[49],stage2_48[87],stage2_47[91]}
   );
   gpc615_5 gpc6857 (
      {stage1_47[230], stage1_47[231], stage1_47[232], stage1_47[233], stage1_47[234]},
      {stage1_48[80]},
      {stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123], stage1_49[124], stage1_49[125]},
      {stage2_51[20],stage2_50[30],stage2_49[50],stage2_48[88],stage2_47[92]}
   );
   gpc615_5 gpc6858 (
      {stage1_47[235], stage1_47[236], stage1_47[237], stage1_47[238], stage1_47[239]},
      {stage1_48[81]},
      {stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129], stage1_49[130], stage1_49[131]},
      {stage2_51[21],stage2_50[31],stage2_49[51],stage2_48[89],stage2_47[93]}
   );
   gpc615_5 gpc6859 (
      {stage1_47[240], stage1_47[241], stage1_47[242], stage1_47[243], stage1_47[244]},
      {stage1_48[82]},
      {stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135], stage1_49[136], stage1_49[137]},
      {stage2_51[22],stage2_50[32],stage2_49[52],stage2_48[90],stage2_47[94]}
   );
   gpc615_5 gpc6860 (
      {stage1_47[245], stage1_47[246], stage1_47[247], stage1_47[248], stage1_47[249]},
      {stage1_48[83]},
      {stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141], stage1_49[142], stage1_49[143]},
      {stage2_51[23],stage2_50[33],stage2_49[53],stage2_48[91],stage2_47[95]}
   );
   gpc615_5 gpc6861 (
      {stage1_47[250], stage1_47[251], stage1_47[252], stage1_47[253], stage1_47[254]},
      {stage1_48[84]},
      {stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147], stage1_49[148], stage1_49[149]},
      {stage2_51[24],stage2_50[34],stage2_49[54],stage2_48[92],stage2_47[96]}
   );
   gpc615_5 gpc6862 (
      {stage1_47[255], stage1_47[256], stage1_47[257], stage1_47[258], stage1_47[259]},
      {stage1_48[85]},
      {stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153], stage1_49[154], stage1_49[155]},
      {stage2_51[25],stage2_50[35],stage2_49[55],stage2_48[93],stage2_47[97]}
   );
   gpc615_5 gpc6863 (
      {stage1_47[260], stage1_47[261], stage1_47[262], stage1_47[263], stage1_47[264]},
      {stage1_48[86]},
      {stage1_49[156], stage1_49[157], stage1_49[158], stage1_49[159], stage1_49[160], stage1_49[161]},
      {stage2_51[26],stage2_50[36],stage2_49[56],stage2_48[94],stage2_47[98]}
   );
   gpc615_5 gpc6864 (
      {stage1_47[265], stage1_47[266], stage1_47[267], stage1_47[268], stage1_47[269]},
      {stage1_48[87]},
      {stage1_49[162], stage1_49[163], stage1_49[164], stage1_49[165], stage1_49[166], stage1_49[167]},
      {stage2_51[27],stage2_50[37],stage2_49[57],stage2_48[95],stage2_47[99]}
   );
   gpc606_5 gpc6865 (
      {stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91], stage1_48[92], stage1_48[93]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[28],stage2_50[38],stage2_49[58],stage2_48[96]}
   );
   gpc606_5 gpc6866 (
      {stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97], stage1_48[98], stage1_48[99]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[29],stage2_50[39],stage2_49[59],stage2_48[97]}
   );
   gpc606_5 gpc6867 (
      {stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103], stage1_48[104], stage1_48[105]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[30],stage2_50[40],stage2_49[60],stage2_48[98]}
   );
   gpc606_5 gpc6868 (
      {stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109], stage1_48[110], stage1_48[111]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[31],stage2_50[41],stage2_49[61],stage2_48[99]}
   );
   gpc606_5 gpc6869 (
      {stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115], stage1_48[116], stage1_48[117]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[32],stage2_50[42],stage2_49[62],stage2_48[100]}
   );
   gpc606_5 gpc6870 (
      {stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121], stage1_48[122], stage1_48[123]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[33],stage2_50[43],stage2_49[63],stage2_48[101]}
   );
   gpc606_5 gpc6871 (
      {stage1_48[124], stage1_48[125], stage1_48[126], stage1_48[127], stage1_48[128], stage1_48[129]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[34],stage2_50[44],stage2_49[64],stage2_48[102]}
   );
   gpc606_5 gpc6872 (
      {stage1_48[130], stage1_48[131], stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[35],stage2_50[45],stage2_49[65],stage2_48[103]}
   );
   gpc606_5 gpc6873 (
      {stage1_48[136], stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[36],stage2_50[46],stage2_49[66],stage2_48[104]}
   );
   gpc606_5 gpc6874 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146], stage1_48[147]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[37],stage2_50[47],stage2_49[67],stage2_48[105]}
   );
   gpc606_5 gpc6875 (
      {stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151], stage1_48[152], stage1_48[153]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[38],stage2_50[48],stage2_49[68],stage2_48[106]}
   );
   gpc606_5 gpc6876 (
      {stage1_48[154], stage1_48[155], stage1_48[156], stage1_48[157], stage1_48[158], stage1_48[159]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[39],stage2_50[49],stage2_49[69],stage2_48[107]}
   );
   gpc606_5 gpc6877 (
      {stage1_48[160], stage1_48[161], stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[40],stage2_50[50],stage2_49[70],stage2_48[108]}
   );
   gpc606_5 gpc6878 (
      {stage1_49[168], stage1_49[169], stage1_49[170], stage1_49[171], stage1_49[172], stage1_49[173]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[13],stage2_51[41],stage2_50[51],stage2_49[71]}
   );
   gpc606_5 gpc6879 (
      {stage1_49[174], stage1_49[175], stage1_49[176], stage1_49[177], stage1_49[178], stage1_49[179]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[14],stage2_51[42],stage2_50[52],stage2_49[72]}
   );
   gpc606_5 gpc6880 (
      {stage1_49[180], stage1_49[181], stage1_49[182], stage1_49[183], stage1_49[184], stage1_49[185]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[15],stage2_51[43],stage2_50[53],stage2_49[73]}
   );
   gpc606_5 gpc6881 (
      {stage1_49[186], stage1_49[187], stage1_49[188], stage1_49[189], stage1_49[190], stage1_49[191]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[16],stage2_51[44],stage2_50[54],stage2_49[74]}
   );
   gpc606_5 gpc6882 (
      {stage1_49[192], stage1_49[193], stage1_49[194], stage1_49[195], stage1_49[196], stage1_49[197]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[17],stage2_51[45],stage2_50[55],stage2_49[75]}
   );
   gpc615_5 gpc6883 (
      {stage1_49[198], stage1_49[199], stage1_49[200], stage1_49[201], stage1_49[202]},
      {stage1_50[78]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[18],stage2_51[46],stage2_50[56],stage2_49[76]}
   );
   gpc1163_5 gpc6884 (
      {stage1_50[79], stage1_50[80], stage1_50[81]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage1_52[0]},
      {stage1_53[0]},
      {stage2_54[0],stage2_53[6],stage2_52[19],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc6885 (
      {stage1_50[82], stage1_50[83], stage1_50[84]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage1_52[1]},
      {stage1_53[1]},
      {stage2_54[1],stage2_53[7],stage2_52[20],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc6886 (
      {stage1_50[85], stage1_50[86], stage1_50[87]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage1_52[2]},
      {stage1_53[2]},
      {stage2_54[2],stage2_53[8],stage2_52[21],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc6887 (
      {stage1_50[88], stage1_50[89], stage1_50[90]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage1_52[3]},
      {stage1_53[3]},
      {stage2_54[3],stage2_53[9],stage2_52[22],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc6888 (
      {stage1_50[91], stage1_50[92], stage1_50[93]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage1_52[4]},
      {stage1_53[4]},
      {stage2_54[4],stage2_53[10],stage2_52[23],stage2_51[51],stage2_50[61]}
   );
   gpc615_5 gpc6889 (
      {stage1_50[94], stage1_50[95], stage1_50[96], stage1_50[97], stage1_50[98]},
      {stage1_51[66]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[11],stage2_52[24],stage2_51[52],stage2_50[62]}
   );
   gpc615_5 gpc6890 (
      {stage1_50[99], stage1_50[100], stage1_50[101], stage1_50[102], stage1_50[103]},
      {stage1_51[67]},
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage2_54[6],stage2_53[12],stage2_52[25],stage2_51[53],stage2_50[63]}
   );
   gpc615_5 gpc6891 (
      {stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107], stage1_50[108]},
      {stage1_51[68]},
      {stage1_52[17], stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22]},
      {stage2_54[7],stage2_53[13],stage2_52[26],stage2_51[54],stage2_50[64]}
   );
   gpc615_5 gpc6892 (
      {stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112], stage1_50[113]},
      {stage1_51[69]},
      {stage1_52[23], stage1_52[24], stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28]},
      {stage2_54[8],stage2_53[14],stage2_52[27],stage2_51[55],stage2_50[65]}
   );
   gpc615_5 gpc6893 (
      {stage1_50[114], stage1_50[115], stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[70]},
      {stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34]},
      {stage2_54[9],stage2_53[15],stage2_52[28],stage2_51[56],stage2_50[66]}
   );
   gpc615_5 gpc6894 (
      {stage1_50[119], stage1_50[120], stage1_50[121], stage1_50[122], stage1_50[123]},
      {stage1_51[71]},
      {stage1_52[35], stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40]},
      {stage2_54[10],stage2_53[16],stage2_52[29],stage2_51[57],stage2_50[67]}
   );
   gpc615_5 gpc6895 (
      {stage1_50[124], stage1_50[125], stage1_50[126], stage1_50[127], stage1_50[128]},
      {stage1_51[72]},
      {stage1_52[41], stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46]},
      {stage2_54[11],stage2_53[17],stage2_52[30],stage2_51[58],stage2_50[68]}
   );
   gpc615_5 gpc6896 (
      {stage1_50[129], stage1_50[130], stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[73]},
      {stage1_52[47], stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52]},
      {stage2_54[12],stage2_53[18],stage2_52[31],stage2_51[59],stage2_50[69]}
   );
   gpc606_5 gpc6897 (
      {stage1_51[74], stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79]},
      {stage1_53[5], stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10]},
      {stage2_55[0],stage2_54[13],stage2_53[19],stage2_52[32],stage2_51[60]}
   );
   gpc606_5 gpc6898 (
      {stage1_51[80], stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85]},
      {stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16]},
      {stage2_55[1],stage2_54[14],stage2_53[20],stage2_52[33],stage2_51[61]}
   );
   gpc606_5 gpc6899 (
      {stage1_51[86], stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91]},
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22]},
      {stage2_55[2],stage2_54[15],stage2_53[21],stage2_52[34],stage2_51[62]}
   );
   gpc606_5 gpc6900 (
      {stage1_51[92], stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97]},
      {stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28]},
      {stage2_55[3],stage2_54[16],stage2_53[22],stage2_52[35],stage2_51[63]}
   );
   gpc606_5 gpc6901 (
      {stage1_51[98], stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103]},
      {stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage2_55[4],stage2_54[17],stage2_53[23],stage2_52[36],stage2_51[64]}
   );
   gpc606_5 gpc6902 (
      {stage1_51[104], stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109]},
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40]},
      {stage2_55[5],stage2_54[18],stage2_53[24],stage2_52[37],stage2_51[65]}
   );
   gpc606_5 gpc6903 (
      {stage1_51[110], stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115]},
      {stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46]},
      {stage2_55[6],stage2_54[19],stage2_53[25],stage2_52[38],stage2_51[66]}
   );
   gpc606_5 gpc6904 (
      {stage1_51[116], stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121]},
      {stage1_53[47], stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52]},
      {stage2_55[7],stage2_54[20],stage2_53[26],stage2_52[39],stage2_51[67]}
   );
   gpc606_5 gpc6905 (
      {stage1_51[122], stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127]},
      {stage1_53[53], stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58]},
      {stage2_55[8],stage2_54[21],stage2_53[27],stage2_52[40],stage2_51[68]}
   );
   gpc606_5 gpc6906 (
      {stage1_51[128], stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133]},
      {stage1_53[59], stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64]},
      {stage2_55[9],stage2_54[22],stage2_53[28],stage2_52[41],stage2_51[69]}
   );
   gpc606_5 gpc6907 (
      {stage1_51[134], stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139]},
      {stage1_53[65], stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70]},
      {stage2_55[10],stage2_54[23],stage2_53[29],stage2_52[42],stage2_51[70]}
   );
   gpc606_5 gpc6908 (
      {stage1_51[140], stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145]},
      {stage1_53[71], stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76]},
      {stage2_55[11],stage2_54[24],stage2_53[30],stage2_52[43],stage2_51[71]}
   );
   gpc606_5 gpc6909 (
      {stage1_51[146], stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151]},
      {stage1_53[77], stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82]},
      {stage2_55[12],stage2_54[25],stage2_53[31],stage2_52[44],stage2_51[72]}
   );
   gpc606_5 gpc6910 (
      {stage1_51[152], stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157]},
      {stage1_53[83], stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88]},
      {stage2_55[13],stage2_54[26],stage2_53[32],stage2_52[45],stage2_51[73]}
   );
   gpc606_5 gpc6911 (
      {stage1_51[158], stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163]},
      {stage1_53[89], stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94]},
      {stage2_55[14],stage2_54[27],stage2_53[33],stage2_52[46],stage2_51[74]}
   );
   gpc606_5 gpc6912 (
      {stage1_51[164], stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169]},
      {stage1_53[95], stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100]},
      {stage2_55[15],stage2_54[28],stage2_53[34],stage2_52[47],stage2_51[75]}
   );
   gpc606_5 gpc6913 (
      {stage1_51[170], stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175]},
      {stage1_53[101], stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106]},
      {stage2_55[16],stage2_54[29],stage2_53[35],stage2_52[48],stage2_51[76]}
   );
   gpc606_5 gpc6914 (
      {stage1_51[176], stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181]},
      {stage1_53[107], stage1_53[108], stage1_53[109], stage1_53[110], stage1_53[111], stage1_53[112]},
      {stage2_55[17],stage2_54[30],stage2_53[36],stage2_52[49],stage2_51[77]}
   );
   gpc606_5 gpc6915 (
      {stage1_51[182], stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187]},
      {stage1_53[113], stage1_53[114], stage1_53[115], stage1_53[116], stage1_53[117], stage1_53[118]},
      {stage2_55[18],stage2_54[31],stage2_53[37],stage2_52[50],stage2_51[78]}
   );
   gpc606_5 gpc6916 (
      {stage1_51[188], stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193]},
      {stage1_53[119], stage1_53[120], stage1_53[121], stage1_53[122], stage1_53[123], stage1_53[124]},
      {stage2_55[19],stage2_54[32],stage2_53[38],stage2_52[51],stage2_51[79]}
   );
   gpc606_5 gpc6917 (
      {stage1_51[194], stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199]},
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129], stage1_53[130]},
      {stage2_55[20],stage2_54[33],stage2_53[39],stage2_52[52],stage2_51[80]}
   );
   gpc606_5 gpc6918 (
      {stage1_51[200], stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_53[131], stage1_53[132], stage1_53[133], stage1_53[134], stage1_53[135], stage1_53[136]},
      {stage2_55[21],stage2_54[34],stage2_53[40],stage2_52[53],stage2_51[81]}
   );
   gpc606_5 gpc6919 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210], stage1_51[211]},
      {stage1_53[137], stage1_53[138], stage1_53[139], stage1_53[140], stage1_53[141], stage1_53[142]},
      {stage2_55[22],stage2_54[35],stage2_53[41],stage2_52[54],stage2_51[82]}
   );
   gpc606_5 gpc6920 (
      {stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215], stage1_51[216], stage1_51[217]},
      {stage1_53[143], stage1_53[144], stage1_53[145], stage1_53[146], stage1_53[147], stage1_53[148]},
      {stage2_55[23],stage2_54[36],stage2_53[42],stage2_52[55],stage2_51[83]}
   );
   gpc606_5 gpc6921 (
      {stage1_51[218], stage1_51[219], stage1_51[220], stage1_51[221], stage1_51[222], stage1_51[223]},
      {stage1_53[149], stage1_53[150], stage1_53[151], stage1_53[152], stage1_53[153], stage1_53[154]},
      {stage2_55[24],stage2_54[37],stage2_53[43],stage2_52[56],stage2_51[84]}
   );
   gpc606_5 gpc6922 (
      {stage1_52[53], stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[25],stage2_54[38],stage2_53[44],stage2_52[57]}
   );
   gpc606_5 gpc6923 (
      {stage1_52[59], stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[26],stage2_54[39],stage2_53[45],stage2_52[58]}
   );
   gpc606_5 gpc6924 (
      {stage1_52[65], stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[27],stage2_54[40],stage2_53[46],stage2_52[59]}
   );
   gpc606_5 gpc6925 (
      {stage1_52[71], stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[28],stage2_54[41],stage2_53[47],stage2_52[60]}
   );
   gpc606_5 gpc6926 (
      {stage1_52[77], stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[29],stage2_54[42],stage2_53[48],stage2_52[61]}
   );
   gpc606_5 gpc6927 (
      {stage1_52[83], stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[30],stage2_54[43],stage2_53[49],stage2_52[62]}
   );
   gpc606_5 gpc6928 (
      {stage1_52[89], stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[31],stage2_54[44],stage2_53[50],stage2_52[63]}
   );
   gpc606_5 gpc6929 (
      {stage1_52[95], stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[32],stage2_54[45],stage2_53[51],stage2_52[64]}
   );
   gpc606_5 gpc6930 (
      {stage1_52[101], stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[33],stage2_54[46],stage2_53[52],stage2_52[65]}
   );
   gpc606_5 gpc6931 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111], stage1_52[112]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[34],stage2_54[47],stage2_53[53],stage2_52[66]}
   );
   gpc606_5 gpc6932 (
      {stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116], stage1_52[117], stage1_52[118]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[35],stage2_54[48],stage2_53[54],stage2_52[67]}
   );
   gpc606_5 gpc6933 (
      {stage1_52[119], stage1_52[120], stage1_52[121], stage1_52[122], stage1_52[123], stage1_52[124]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[36],stage2_54[49],stage2_53[55],stage2_52[68]}
   );
   gpc606_5 gpc6934 (
      {stage1_52[125], stage1_52[126], stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[37],stage2_54[50],stage2_53[56],stage2_52[69]}
   );
   gpc606_5 gpc6935 (
      {stage1_52[131], stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[38],stage2_54[51],stage2_53[57],stage2_52[70]}
   );
   gpc606_5 gpc6936 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141], stage1_52[142]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[39],stage2_54[52],stage2_53[58],stage2_52[71]}
   );
   gpc606_5 gpc6937 (
      {stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146], stage1_52[147], stage1_52[148]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[40],stage2_54[53],stage2_53[59],stage2_52[72]}
   );
   gpc606_5 gpc6938 (
      {stage1_52[149], stage1_52[150], stage1_52[151], stage1_52[152], stage1_52[153], stage1_52[154]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[41],stage2_54[54],stage2_53[60],stage2_52[73]}
   );
   gpc606_5 gpc6939 (
      {stage1_52[155], stage1_52[156], stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[42],stage2_54[55],stage2_53[61],stage2_52[74]}
   );
   gpc606_5 gpc6940 (
      {stage1_52[161], stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[43],stage2_54[56],stage2_53[62],stage2_52[75]}
   );
   gpc606_5 gpc6941 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171], stage1_52[172]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[44],stage2_54[57],stage2_53[63],stage2_52[76]}
   );
   gpc606_5 gpc6942 (
      {stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176], stage1_52[177], stage1_52[178]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[45],stage2_54[58],stage2_53[64],stage2_52[77]}
   );
   gpc606_5 gpc6943 (
      {stage1_52[179], stage1_52[180], stage1_52[181], stage1_52[182], stage1_52[183], stage1_52[184]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[46],stage2_54[59],stage2_53[65],stage2_52[78]}
   );
   gpc606_5 gpc6944 (
      {stage1_52[185], stage1_52[186], stage1_52[187], stage1_52[188], stage1_52[189], stage1_52[190]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[47],stage2_54[60],stage2_53[66],stage2_52[79]}
   );
   gpc606_5 gpc6945 (
      {stage1_52[191], stage1_52[192], stage1_52[193], stage1_52[194], stage1_52[195], stage1_52[196]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[48],stage2_54[61],stage2_53[67],stage2_52[80]}
   );
   gpc606_5 gpc6946 (
      {stage1_52[197], stage1_52[198], stage1_52[199], stage1_52[200], stage1_52[201], stage1_52[202]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[49],stage2_54[62],stage2_53[68],stage2_52[81]}
   );
   gpc606_5 gpc6947 (
      {stage1_52[203], stage1_52[204], stage1_52[205], stage1_52[206], stage1_52[207], stage1_52[208]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[50],stage2_54[63],stage2_53[69],stage2_52[82]}
   );
   gpc606_5 gpc6948 (
      {stage1_52[209], stage1_52[210], stage1_52[211], stage1_52[212], stage1_52[213], stage1_52[214]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[51],stage2_54[64],stage2_53[70],stage2_52[83]}
   );
   gpc606_5 gpc6949 (
      {stage1_52[215], stage1_52[216], stage1_52[217], stage1_52[218], stage1_52[219], stage1_52[220]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[52],stage2_54[65],stage2_53[71],stage2_52[84]}
   );
   gpc606_5 gpc6950 (
      {stage1_52[221], stage1_52[222], stage1_52[223], stage1_52[224], stage1_52[225], stage1_52[226]},
      {stage1_54[168], stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173]},
      {stage2_56[28],stage2_55[53],stage2_54[66],stage2_53[72],stage2_52[85]}
   );
   gpc606_5 gpc6951 (
      {stage1_52[227], stage1_52[228], stage1_52[229], stage1_52[230], stage1_52[231], stage1_52[232]},
      {stage1_54[174], stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179]},
      {stage2_56[29],stage2_55[54],stage2_54[67],stage2_53[73],stage2_52[86]}
   );
   gpc606_5 gpc6952 (
      {stage1_52[233], stage1_52[234], stage1_52[235], stage1_52[236], stage1_52[237], stage1_52[238]},
      {stage1_54[180], stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185]},
      {stage2_56[30],stage2_55[55],stage2_54[68],stage2_53[74],stage2_52[87]}
   );
   gpc606_5 gpc6953 (
      {stage1_52[239], stage1_52[240], stage1_52[241], stage1_52[242], stage1_52[243], stage1_52[244]},
      {stage1_54[186], stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191]},
      {stage2_56[31],stage2_55[56],stage2_54[69],stage2_53[75],stage2_52[88]}
   );
   gpc606_5 gpc6954 (
      {stage1_52[245], stage1_52[246], stage1_52[247], stage1_52[248], stage1_52[249], stage1_52[250]},
      {stage1_54[192], stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage2_56[32],stage2_55[57],stage2_54[70],stage2_53[76],stage2_52[89]}
   );
   gpc606_5 gpc6955 (
      {stage1_52[251], stage1_52[252], stage1_52[253], stage1_52[254], stage1_52[255], stage1_52[256]},
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202], stage1_54[203]},
      {stage2_56[33],stage2_55[58],stage2_54[71],stage2_53[77],stage2_52[90]}
   );
   gpc606_5 gpc6956 (
      {stage1_52[257], stage1_52[258], stage1_52[259], stage1_52[260], stage1_52[261], stage1_52[262]},
      {stage1_54[204], stage1_54[205], stage1_54[206], stage1_54[207], stage1_54[208], stage1_54[209]},
      {stage2_56[34],stage2_55[59],stage2_54[72],stage2_53[78],stage2_52[91]}
   );
   gpc606_5 gpc6957 (
      {stage1_52[263], stage1_52[264], stage1_52[265], stage1_52[266], stage1_52[267], stage1_52[268]},
      {stage1_54[210], stage1_54[211], stage1_54[212], stage1_54[213], stage1_54[214], stage1_54[215]},
      {stage2_56[35],stage2_55[60],stage2_54[73],stage2_53[79],stage2_52[92]}
   );
   gpc606_5 gpc6958 (
      {stage1_53[155], stage1_53[156], stage1_53[157], stage1_53[158], stage1_53[159], stage1_53[160]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[36],stage2_55[61],stage2_54[74],stage2_53[80]}
   );
   gpc606_5 gpc6959 (
      {stage1_53[161], stage1_53[162], stage1_53[163], stage1_53[164], stage1_53[165], stage1_53[166]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[37],stage2_55[62],stage2_54[75],stage2_53[81]}
   );
   gpc606_5 gpc6960 (
      {stage1_53[167], stage1_53[168], stage1_53[169], stage1_53[170], stage1_53[171], stage1_53[172]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[38],stage2_55[63],stage2_54[76],stage2_53[82]}
   );
   gpc2135_5 gpc6961 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[0], stage1_56[1], stage1_56[2]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[0],stage2_57[3],stage2_56[39],stage2_55[64]}
   );
   gpc2135_5 gpc6962 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[1],stage2_57[4],stage2_56[40],stage2_55[65]}
   );
   gpc2135_5 gpc6963 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[6], stage1_56[7], stage1_56[8]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[2],stage2_57[5],stage2_56[41],stage2_55[66]}
   );
   gpc2135_5 gpc6964 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[3],stage2_57[6],stage2_56[42],stage2_55[67]}
   );
   gpc2135_5 gpc6965 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12], stage1_56[13], stage1_56[14]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[4],stage2_57[7],stage2_56[43],stage2_55[68]}
   );
   gpc2135_5 gpc6966 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[5],stage2_57[8],stage2_56[44],stage2_55[69]}
   );
   gpc2135_5 gpc6967 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[18], stage1_56[19], stage1_56[20]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[6],stage2_57[9],stage2_56[45],stage2_55[70]}
   );
   gpc2135_5 gpc6968 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[7],stage2_57[10],stage2_56[46],stage2_55[71]}
   );
   gpc2135_5 gpc6969 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[24], stage1_56[25], stage1_56[26]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[8],stage2_57[11],stage2_56[47],stage2_55[72]}
   );
   gpc2135_5 gpc6970 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[9],stage2_57[12],stage2_56[48],stage2_55[73]}
   );
   gpc2135_5 gpc6971 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[30], stage1_56[31], stage1_56[32]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[10],stage2_57[13],stage2_56[49],stage2_55[74]}
   );
   gpc2135_5 gpc6972 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[11],stage2_57[14],stage2_56[50],stage2_55[75]}
   );
   gpc2135_5 gpc6973 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[12],stage2_57[15],stage2_56[51],stage2_55[76]}
   );
   gpc2135_5 gpc6974 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[13],stage2_57[16],stage2_56[52],stage2_55[77]}
   );
   gpc2135_5 gpc6975 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[14],stage2_57[17],stage2_56[53],stage2_55[78]}
   );
   gpc2135_5 gpc6976 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[15],stage2_57[18],stage2_56[54],stage2_55[79]}
   );
   gpc2135_5 gpc6977 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[16],stage2_57[19],stage2_56[55],stage2_55[80]}
   );
   gpc2135_5 gpc6978 (
      {stage1_55[103], stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[17],stage2_57[20],stage2_56[56],stage2_55[81]}
   );
   gpc2135_5 gpc6979 (
      {stage1_55[108], stage1_55[109], stage1_55[110], stage1_55[111], stage1_55[112]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[18]},
      {stage1_58[36], stage1_58[37]},
      {stage2_59[18],stage2_58[18],stage2_57[21],stage2_56[57],stage2_55[82]}
   );
   gpc2135_5 gpc6980 (
      {stage1_55[113], stage1_55[114], stage1_55[115], stage1_55[116], stage1_55[117]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[19]},
      {stage1_58[38], stage1_58[39]},
      {stage2_59[19],stage2_58[19],stage2_57[22],stage2_56[58],stage2_55[83]}
   );
   gpc2135_5 gpc6981 (
      {stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121], stage1_55[122]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[20]},
      {stage1_58[40], stage1_58[41]},
      {stage2_59[20],stage2_58[20],stage2_57[23],stage2_56[59],stage2_55[84]}
   );
   gpc2135_5 gpc6982 (
      {stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[21]},
      {stage1_58[42], stage1_58[43]},
      {stage2_59[21],stage2_58[21],stage2_57[24],stage2_56[60],stage2_55[85]}
   );
   gpc2135_5 gpc6983 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[22]},
      {stage1_58[44], stage1_58[45]},
      {stage2_59[22],stage2_58[22],stage2_57[25],stage2_56[61],stage2_55[86]}
   );
   gpc2135_5 gpc6984 (
      {stage1_55[133], stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[23]},
      {stage1_58[46], stage1_58[47]},
      {stage2_59[23],stage2_58[23],stage2_57[26],stage2_56[62],stage2_55[87]}
   );
   gpc2135_5 gpc6985 (
      {stage1_55[138], stage1_55[139], stage1_55[140], stage1_55[141], stage1_55[142]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[24]},
      {stage1_58[48], stage1_58[49]},
      {stage2_59[24],stage2_58[24],stage2_57[27],stage2_56[63],stage2_55[88]}
   );
   gpc2135_5 gpc6986 (
      {stage1_55[143], stage1_55[144], stage1_55[145], stage1_55[146], stage1_55[147]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[25]},
      {stage1_58[50], stage1_58[51]},
      {stage2_59[25],stage2_58[25],stage2_57[28],stage2_56[64],stage2_55[89]}
   );
   gpc2135_5 gpc6987 (
      {stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151], stage1_55[152]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[26]},
      {stage1_58[52], stage1_58[53]},
      {stage2_59[26],stage2_58[26],stage2_57[29],stage2_56[65],stage2_55[90]}
   );
   gpc2135_5 gpc6988 (
      {stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[27]},
      {stage1_58[54], stage1_58[55]},
      {stage2_59[27],stage2_58[27],stage2_57[30],stage2_56[66],stage2_55[91]}
   );
   gpc2135_5 gpc6989 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[28]},
      {stage1_58[56], stage1_58[57]},
      {stage2_59[28],stage2_58[28],stage2_57[31],stage2_56[67],stage2_55[92]}
   );
   gpc2135_5 gpc6990 (
      {stage1_55[163], stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[29]},
      {stage1_58[58], stage1_58[59]},
      {stage2_59[29],stage2_58[29],stage2_57[32],stage2_56[68],stage2_55[93]}
   );
   gpc606_5 gpc6991 (
      {stage1_55[168], stage1_55[169], stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[30],stage2_58[30],stage2_57[33],stage2_56[69],stage2_55[94]}
   );
   gpc615_5 gpc6992 (
      {stage1_55[174], stage1_55[175], stage1_55[176], stage1_55[177], stage1_55[178]},
      {stage1_56[90]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[31],stage2_58[31],stage2_57[34],stage2_56[70],stage2_55[95]}
   );
   gpc615_5 gpc6993 (
      {stage1_55[179], stage1_55[180], stage1_55[181], stage1_55[182], stage1_55[183]},
      {stage1_56[91]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[32],stage2_58[32],stage2_57[35],stage2_56[71],stage2_55[96]}
   );
   gpc615_5 gpc6994 (
      {stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187], stage1_55[188]},
      {stage1_56[92]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[33],stage2_58[33],stage2_57[36],stage2_56[72],stage2_55[97]}
   );
   gpc615_5 gpc6995 (
      {stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_56[93]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[34],stage2_58[34],stage2_57[37],stage2_56[73],stage2_55[98]}
   );
   gpc615_5 gpc6996 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198]},
      {stage1_56[94]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[35],stage2_58[35],stage2_57[38],stage2_56[74],stage2_55[99]}
   );
   gpc615_5 gpc6997 (
      {stage1_55[199], stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203]},
      {stage1_56[95]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[36],stage2_58[36],stage2_57[39],stage2_56[75],stage2_55[100]}
   );
   gpc615_5 gpc6998 (
      {stage1_55[204], stage1_55[205], stage1_55[206], stage1_55[207], stage1_55[208]},
      {stage1_56[96]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[37],stage2_58[37],stage2_57[40],stage2_56[76],stage2_55[101]}
   );
   gpc615_5 gpc6999 (
      {stage1_55[209], stage1_55[210], stage1_55[211], stage1_55[212], stage1_55[213]},
      {stage1_56[97]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[38],stage2_58[38],stage2_57[41],stage2_56[77],stage2_55[102]}
   );
   gpc615_5 gpc7000 (
      {stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217], stage1_55[218]},
      {stage1_56[98]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[39],stage2_58[39],stage2_57[42],stage2_56[78],stage2_55[103]}
   );
   gpc606_5 gpc7001 (
      {stage1_56[99], stage1_56[100], stage1_56[101], stage1_56[102], stage1_56[103], stage1_56[104]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[0],stage2_59[40],stage2_58[40],stage2_57[43],stage2_56[79]}
   );
   gpc606_5 gpc7002 (
      {stage1_56[105], stage1_56[106], stage1_56[107], stage1_56[108], stage1_56[109], stage1_56[110]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[1],stage2_59[41],stage2_58[41],stage2_57[44],stage2_56[80]}
   );
   gpc606_5 gpc7003 (
      {stage1_56[111], stage1_56[112], stage1_56[113], stage1_56[114], stage1_56[115], stage1_56[116]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[2],stage2_59[42],stage2_58[42],stage2_57[45],stage2_56[81]}
   );
   gpc606_5 gpc7004 (
      {stage1_56[117], stage1_56[118], stage1_56[119], stage1_56[120], stage1_56[121], stage1_56[122]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[3],stage2_59[43],stage2_58[43],stage2_57[46],stage2_56[82]}
   );
   gpc606_5 gpc7005 (
      {stage1_56[123], stage1_56[124], stage1_56[125], stage1_56[126], stage1_56[127], stage1_56[128]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[4],stage2_59[44],stage2_58[44],stage2_57[47],stage2_56[83]}
   );
   gpc606_5 gpc7006 (
      {stage1_56[129], stage1_56[130], stage1_56[131], stage1_56[132], stage1_56[133], stage1_56[134]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[5],stage2_59[45],stage2_58[45],stage2_57[48],stage2_56[84]}
   );
   gpc606_5 gpc7007 (
      {stage1_56[135], stage1_56[136], stage1_56[137], stage1_56[138], stage1_56[139], stage1_56[140]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[6],stage2_59[46],stage2_58[46],stage2_57[49],stage2_56[85]}
   );
   gpc606_5 gpc7008 (
      {stage1_56[141], stage1_56[142], stage1_56[143], stage1_56[144], stage1_56[145], stage1_56[146]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[7],stage2_59[47],stage2_58[47],stage2_57[50],stage2_56[86]}
   );
   gpc606_5 gpc7009 (
      {stage1_56[147], stage1_56[148], stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[8],stage2_59[48],stage2_58[48],stage2_57[51],stage2_56[87]}
   );
   gpc606_5 gpc7010 (
      {stage1_56[153], stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_58[114], stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage2_60[9],stage2_59[49],stage2_58[49],stage2_57[52],stage2_56[88]}
   );
   gpc606_5 gpc7011 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163], stage1_56[164]},
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124], stage1_58[125]},
      {stage2_60[10],stage2_59[50],stage2_58[50],stage2_57[53],stage2_56[89]}
   );
   gpc606_5 gpc7012 (
      {stage1_56[165], stage1_56[166], stage1_56[167], stage1_56[168], stage1_56[169], stage1_56[170]},
      {stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129], stage1_58[130], stage1_58[131]},
      {stage2_60[11],stage2_59[51],stage2_58[51],stage2_57[54],stage2_56[90]}
   );
   gpc606_5 gpc7013 (
      {stage1_56[171], stage1_56[172], stage1_56[173], stage1_56[174], stage1_56[175], stage1_56[176]},
      {stage1_58[132], stage1_58[133], stage1_58[134], stage1_58[135], stage1_58[136], stage1_58[137]},
      {stage2_60[12],stage2_59[52],stage2_58[52],stage2_57[55],stage2_56[91]}
   );
   gpc606_5 gpc7014 (
      {stage1_56[177], stage1_56[178], stage1_56[179], stage1_56[180], stage1_56[181], stage1_56[182]},
      {stage1_58[138], stage1_58[139], stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143]},
      {stage2_60[13],stage2_59[53],stage2_58[53],stage2_57[56],stage2_56[92]}
   );
   gpc606_5 gpc7015 (
      {stage1_56[183], stage1_56[184], stage1_56[185], stage1_56[186], stage1_56[187], stage1_56[188]},
      {stage1_58[144], stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage2_60[14],stage2_59[54],stage2_58[54],stage2_57[57],stage2_56[93]}
   );
   gpc606_5 gpc7016 (
      {stage1_56[189], stage1_56[190], stage1_56[191], stage1_56[192], stage1_56[193], stage1_56[194]},
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154], stage1_58[155]},
      {stage2_60[15],stage2_59[55],stage2_58[55],stage2_57[58],stage2_56[94]}
   );
   gpc606_5 gpc7017 (
      {stage1_56[195], stage1_56[196], stage1_56[197], stage1_56[198], stage1_56[199], stage1_56[200]},
      {stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159], stage1_58[160], stage1_58[161]},
      {stage2_60[16],stage2_59[56],stage2_58[56],stage2_57[59],stage2_56[95]}
   );
   gpc606_5 gpc7018 (
      {stage1_56[201], stage1_56[202], stage1_56[203], stage1_56[204], stage1_56[205], stage1_56[206]},
      {stage1_58[162], stage1_58[163], stage1_58[164], stage1_58[165], stage1_58[166], stage1_58[167]},
      {stage2_60[17],stage2_59[57],stage2_58[57],stage2_57[60],stage2_56[96]}
   );
   gpc606_5 gpc7019 (
      {stage1_56[207], stage1_56[208], stage1_56[209], stage1_56[210], stage1_56[211], stage1_56[212]},
      {stage1_58[168], stage1_58[169], stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173]},
      {stage2_60[18],stage2_59[58],stage2_58[58],stage2_57[61],stage2_56[97]}
   );
   gpc606_5 gpc7020 (
      {stage1_56[213], stage1_56[214], stage1_56[215], stage1_56[216], stage1_56[217], stage1_56[218]},
      {stage1_58[174], stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage2_60[19],stage2_59[59],stage2_58[59],stage2_57[62],stage2_56[98]}
   );
   gpc606_5 gpc7021 (
      {stage1_56[219], stage1_56[220], stage1_56[221], stage1_56[222], stage1_56[223], stage1_56[224]},
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184], stage1_58[185]},
      {stage2_60[20],stage2_59[60],stage2_58[60],stage2_57[63],stage2_56[99]}
   );
   gpc606_5 gpc7022 (
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[21],stage2_59[61],stage2_58[61],stage2_57[64]}
   );
   gpc606_5 gpc7023 (
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[22],stage2_59[62],stage2_58[62],stage2_57[65]}
   );
   gpc606_5 gpc7024 (
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[23],stage2_59[63],stage2_58[63],stage2_57[66]}
   );
   gpc606_5 gpc7025 (
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[24],stage2_59[64],stage2_58[64],stage2_57[67]}
   );
   gpc606_5 gpc7026 (
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage2_61[4],stage2_60[25],stage2_59[65],stage2_58[65],stage2_57[68]}
   );
   gpc606_5 gpc7027 (
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage2_61[5],stage2_60[26],stage2_59[66],stage2_58[66],stage2_57[69]}
   );
   gpc606_5 gpc7028 (
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage2_61[6],stage2_60[27],stage2_59[67],stage2_58[67],stage2_57[70]}
   );
   gpc606_5 gpc7029 (
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage1_59[42], stage1_59[43], stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47]},
      {stage2_61[7],stage2_60[28],stage2_59[68],stage2_58[68],stage2_57[71]}
   );
   gpc606_5 gpc7030 (
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage1_59[48], stage1_59[49], stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53]},
      {stage2_61[8],stage2_60[29],stage2_59[69],stage2_58[69],stage2_57[72]}
   );
   gpc606_5 gpc7031 (
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage1_59[54], stage1_59[55], stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59]},
      {stage2_61[9],stage2_60[30],stage2_59[70],stage2_58[70],stage2_57[73]}
   );
   gpc606_5 gpc7032 (
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage1_59[60], stage1_59[61], stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65]},
      {stage2_61[10],stage2_60[31],stage2_59[71],stage2_58[71],stage2_57[74]}
   );
   gpc606_5 gpc7033 (
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage1_59[66], stage1_59[67], stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71]},
      {stage2_61[11],stage2_60[32],stage2_59[72],stage2_58[72],stage2_57[75]}
   );
   gpc606_5 gpc7034 (
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage1_59[72], stage1_59[73], stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77]},
      {stage2_61[12],stage2_60[33],stage2_59[73],stage2_58[73],stage2_57[76]}
   );
   gpc606_5 gpc7035 (
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage1_59[78], stage1_59[79], stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83]},
      {stage2_61[13],stage2_60[34],stage2_59[74],stage2_58[74],stage2_57[77]}
   );
   gpc606_5 gpc7036 (
      {stage1_57[174], stage1_57[175], stage1_57[176], stage1_57[177], stage1_57[178], stage1_57[179]},
      {stage1_59[84], stage1_59[85], stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89]},
      {stage2_61[14],stage2_60[35],stage2_59[75],stage2_58[75],stage2_57[78]}
   );
   gpc117_4 gpc7037 (
      {stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189], stage1_58[190], stage1_58[191], stage1_58[192]},
      {stage1_59[90]},
      {stage1_60[0]},
      {stage2_61[15],stage2_60[36],stage2_59[76],stage2_58[76]}
   );
   gpc117_4 gpc7038 (
      {stage1_58[193], stage1_58[194], stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[91]},
      {stage1_60[1]},
      {stage2_61[16],stage2_60[37],stage2_59[77],stage2_58[77]}
   );
   gpc117_4 gpc7039 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204], stage1_58[205], stage1_58[206]},
      {stage1_59[92]},
      {stage1_60[2]},
      {stage2_61[17],stage2_60[38],stage2_59[78],stage2_58[78]}
   );
   gpc117_4 gpc7040 (
      {stage1_58[207], stage1_58[208], stage1_58[209], stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213]},
      {stage1_59[93]},
      {stage1_60[3]},
      {stage2_61[18],stage2_60[39],stage2_59[79],stage2_58[79]}
   );
   gpc606_5 gpc7041 (
      {stage1_58[214], stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_60[4], stage1_60[5], stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9]},
      {stage2_62[0],stage2_61[19],stage2_60[40],stage2_59[80],stage2_58[80]}
   );
   gpc606_5 gpc7042 (
      {stage1_58[220], stage1_58[221], stage1_58[222], stage1_58[223], stage1_58[224], stage1_58[225]},
      {stage1_60[10], stage1_60[11], stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15]},
      {stage2_62[1],stage2_61[20],stage2_60[41],stage2_59[81],stage2_58[81]}
   );
   gpc606_5 gpc7043 (
      {stage1_58[226], stage1_58[227], stage1_58[228], stage1_58[229], stage1_58[230], stage1_58[231]},
      {stage1_60[16], stage1_60[17], stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21]},
      {stage2_62[2],stage2_61[21],stage2_60[42],stage2_59[82],stage2_58[82]}
   );
   gpc606_5 gpc7044 (
      {stage1_58[232], stage1_58[233], stage1_58[234], stage1_58[235], stage1_58[236], stage1_58[237]},
      {stage1_60[22], stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage2_62[3],stage2_61[22],stage2_60[43],stage2_59[83],stage2_58[83]}
   );
   gpc606_5 gpc7045 (
      {stage1_58[238], stage1_58[239], stage1_58[240], stage1_58[241], stage1_58[242], 1'b0},
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33]},
      {stage2_62[4],stage2_61[23],stage2_60[44],stage2_59[84],stage2_58[84]}
   );
   gpc606_5 gpc7046 (
      {stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97], stage1_59[98], stage1_59[99]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[24],stage2_60[45],stage2_59[85]}
   );
   gpc606_5 gpc7047 (
      {stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103], stage1_59[104], stage1_59[105]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[25],stage2_60[46],stage2_59[86]}
   );
   gpc606_5 gpc7048 (
      {stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109], stage1_59[110], stage1_59[111]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[26],stage2_60[47],stage2_59[87]}
   );
   gpc606_5 gpc7049 (
      {stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115], stage1_59[116], stage1_59[117]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[27],stage2_60[48],stage2_59[88]}
   );
   gpc606_5 gpc7050 (
      {stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121], stage1_59[122], stage1_59[123]},
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage2_63[4],stage2_62[9],stage2_61[28],stage2_60[49],stage2_59[89]}
   );
   gpc606_5 gpc7051 (
      {stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127], stage1_59[128], stage1_59[129]},
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage2_63[5],stage2_62[10],stage2_61[29],stage2_60[50],stage2_59[90]}
   );
   gpc606_5 gpc7052 (
      {stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133], stage1_59[134], stage1_59[135]},
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage2_63[6],stage2_62[11],stage2_61[30],stage2_60[51],stage2_59[91]}
   );
   gpc606_5 gpc7053 (
      {stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139], stage1_59[140], stage1_59[141]},
      {stage1_61[42], stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage2_63[7],stage2_62[12],stage2_61[31],stage2_60[52],stage2_59[92]}
   );
   gpc606_5 gpc7054 (
      {stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145], stage1_59[146], stage1_59[147]},
      {stage1_61[48], stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53]},
      {stage2_63[8],stage2_62[13],stage2_61[32],stage2_60[53],stage2_59[93]}
   );
   gpc606_5 gpc7055 (
      {stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151], stage1_59[152], stage1_59[153]},
      {stage1_61[54], stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59]},
      {stage2_63[9],stage2_62[14],stage2_61[33],stage2_60[54],stage2_59[94]}
   );
   gpc606_5 gpc7056 (
      {stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157], stage1_59[158], stage1_59[159]},
      {stage1_61[60], stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65]},
      {stage2_63[10],stage2_62[15],stage2_61[34],stage2_60[55],stage2_59[95]}
   );
   gpc606_5 gpc7057 (
      {stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163], stage1_59[164], stage1_59[165]},
      {stage1_61[66], stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71]},
      {stage2_63[11],stage2_62[16],stage2_61[35],stage2_60[56],stage2_59[96]}
   );
   gpc606_5 gpc7058 (
      {stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169], stage1_59[170], stage1_59[171]},
      {stage1_61[72], stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77]},
      {stage2_63[12],stage2_62[17],stage2_61[36],stage2_60[57],stage2_59[97]}
   );
   gpc606_5 gpc7059 (
      {stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175], stage1_59[176], stage1_59[177]},
      {stage1_61[78], stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83]},
      {stage2_63[13],stage2_62[18],stage2_61[37],stage2_60[58],stage2_59[98]}
   );
   gpc606_5 gpc7060 (
      {stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181], stage1_59[182], stage1_59[183]},
      {stage1_61[84], stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89]},
      {stage2_63[14],stage2_62[19],stage2_61[38],stage2_60[59],stage2_59[99]}
   );
   gpc606_5 gpc7061 (
      {stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187], stage1_59[188], stage1_59[189]},
      {stage1_61[90], stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95]},
      {stage2_63[15],stage2_62[20],stage2_61[39],stage2_60[60],stage2_59[100]}
   );
   gpc606_5 gpc7062 (
      {stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193], stage1_59[194], stage1_59[195]},
      {stage1_61[96], stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101]},
      {stage2_63[16],stage2_62[21],stage2_61[40],stage2_60[61],stage2_59[101]}
   );
   gpc606_5 gpc7063 (
      {stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199], stage1_59[200], stage1_59[201]},
      {stage1_61[102], stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107]},
      {stage2_63[17],stage2_62[22],stage2_61[41],stage2_60[62],stage2_59[102]}
   );
   gpc606_5 gpc7064 (
      {stage1_59[202], stage1_59[203], stage1_59[204], stage1_59[205], stage1_59[206], stage1_59[207]},
      {stage1_61[108], stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113]},
      {stage2_63[18],stage2_62[23],stage2_61[42],stage2_60[63],stage2_59[103]}
   );
   gpc606_5 gpc7065 (
      {stage1_59[208], stage1_59[209], stage1_59[210], stage1_59[211], stage1_59[212], stage1_59[213]},
      {stage1_61[114], stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119]},
      {stage2_63[19],stage2_62[24],stage2_61[43],stage2_60[64],stage2_59[104]}
   );
   gpc606_5 gpc7066 (
      {stage1_59[214], stage1_59[215], stage1_59[216], stage1_59[217], stage1_59[218], stage1_59[219]},
      {stage1_61[120], stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125]},
      {stage2_63[20],stage2_62[25],stage2_61[44],stage2_60[65],stage2_59[105]}
   );
   gpc606_5 gpc7067 (
      {stage1_59[220], stage1_59[221], stage1_59[222], stage1_59[223], stage1_59[224], stage1_59[225]},
      {stage1_61[126], stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131]},
      {stage2_63[21],stage2_62[26],stage2_61[45],stage2_60[66],stage2_59[106]}
   );
   gpc606_5 gpc7068 (
      {stage1_59[226], stage1_59[227], stage1_59[228], stage1_59[229], stage1_59[230], stage1_59[231]},
      {stage1_61[132], stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137]},
      {stage2_63[22],stage2_62[27],stage2_61[46],stage2_60[67],stage2_59[107]}
   );
   gpc606_5 gpc7069 (
      {stage1_59[232], stage1_59[233], stage1_59[234], stage1_59[235], stage1_59[236], stage1_59[237]},
      {stage1_61[138], stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143]},
      {stage2_63[23],stage2_62[28],stage2_61[47],stage2_60[68],stage2_59[108]}
   );
   gpc606_5 gpc7070 (
      {stage1_59[238], stage1_59[239], stage1_59[240], stage1_59[241], stage1_59[242], stage1_59[243]},
      {stage1_61[144], stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149]},
      {stage2_63[24],stage2_62[29],stage2_61[48],stage2_60[69],stage2_59[109]}
   );
   gpc606_5 gpc7071 (
      {stage1_59[244], stage1_59[245], stage1_59[246], stage1_59[247], stage1_59[248], stage1_59[249]},
      {stage1_61[150], stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155]},
      {stage2_63[25],stage2_62[30],stage2_61[49],stage2_60[70],stage2_59[110]}
   );
   gpc606_5 gpc7072 (
      {stage1_59[250], stage1_59[251], stage1_59[252], stage1_59[253], stage1_59[254], stage1_59[255]},
      {stage1_61[156], stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161]},
      {stage2_63[26],stage2_62[31],stage2_61[50],stage2_60[71],stage2_59[111]}
   );
   gpc606_5 gpc7073 (
      {stage1_59[256], stage1_59[257], stage1_59[258], stage1_59[259], stage1_59[260], stage1_59[261]},
      {stage1_61[162], stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167]},
      {stage2_63[27],stage2_62[32],stage2_61[51],stage2_60[72],stage2_59[112]}
   );
   gpc606_5 gpc7074 (
      {stage1_59[262], stage1_59[263], stage1_59[264], stage1_59[265], stage1_59[266], stage1_59[267]},
      {stage1_61[168], stage1_61[169], stage1_61[170], stage1_61[171], stage1_61[172], stage1_61[173]},
      {stage2_63[28],stage2_62[33],stage2_61[52],stage2_60[73],stage2_59[113]}
   );
   gpc1406_5 gpc7075 (
      {stage1_60[34], stage1_60[35], stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3]},
      {stage1_63[0]},
      {stage2_64[0],stage2_63[29],stage2_62[34],stage2_61[53],stage2_60[74]}
   );
   gpc606_5 gpc7076 (
      {stage1_60[40], stage1_60[41], stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45]},
      {stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9]},
      {stage2_64[1],stage2_63[30],stage2_62[35],stage2_61[54],stage2_60[75]}
   );
   gpc606_5 gpc7077 (
      {stage1_60[46], stage1_60[47], stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51]},
      {stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15]},
      {stage2_64[2],stage2_63[31],stage2_62[36],stage2_61[55],stage2_60[76]}
   );
   gpc606_5 gpc7078 (
      {stage1_60[52], stage1_60[53], stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57]},
      {stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21]},
      {stage2_64[3],stage2_63[32],stage2_62[37],stage2_61[56],stage2_60[77]}
   );
   gpc606_5 gpc7079 (
      {stage1_60[58], stage1_60[59], stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63]},
      {stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27]},
      {stage2_64[4],stage2_63[33],stage2_62[38],stage2_61[57],stage2_60[78]}
   );
   gpc606_5 gpc7080 (
      {stage1_60[64], stage1_60[65], stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69]},
      {stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33]},
      {stage2_64[5],stage2_63[34],stage2_62[39],stage2_61[58],stage2_60[79]}
   );
   gpc606_5 gpc7081 (
      {stage1_60[70], stage1_60[71], stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75]},
      {stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39]},
      {stage2_64[6],stage2_63[35],stage2_62[40],stage2_61[59],stage2_60[80]}
   );
   gpc606_5 gpc7082 (
      {stage1_60[76], stage1_60[77], stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81]},
      {stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage2_64[7],stage2_63[36],stage2_62[41],stage2_61[60],stage2_60[81]}
   );
   gpc606_5 gpc7083 (
      {stage1_60[82], stage1_60[83], stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87]},
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51]},
      {stage2_64[8],stage2_63[37],stage2_62[42],stage2_61[61],stage2_60[82]}
   );
   gpc606_5 gpc7084 (
      {stage1_60[88], stage1_60[89], stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93]},
      {stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57]},
      {stage2_64[9],stage2_63[38],stage2_62[43],stage2_61[62],stage2_60[83]}
   );
   gpc606_5 gpc7085 (
      {stage1_60[94], stage1_60[95], stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99]},
      {stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63]},
      {stage2_64[10],stage2_63[39],stage2_62[44],stage2_61[63],stage2_60[84]}
   );
   gpc606_5 gpc7086 (
      {stage1_60[100], stage1_60[101], stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105]},
      {stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69]},
      {stage2_64[11],stage2_63[40],stage2_62[45],stage2_61[64],stage2_60[85]}
   );
   gpc606_5 gpc7087 (
      {stage1_60[106], stage1_60[107], stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111]},
      {stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75]},
      {stage2_64[12],stage2_63[41],stage2_62[46],stage2_61[65],stage2_60[86]}
   );
   gpc606_5 gpc7088 (
      {stage1_60[112], stage1_60[113], stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117]},
      {stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79], stage1_62[80], stage1_62[81]},
      {stage2_64[13],stage2_63[42],stage2_62[47],stage2_61[66],stage2_60[87]}
   );
   gpc606_5 gpc7089 (
      {stage1_60[118], stage1_60[119], stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123]},
      {stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85], stage1_62[86], stage1_62[87]},
      {stage2_64[14],stage2_63[43],stage2_62[48],stage2_61[67],stage2_60[88]}
   );
   gpc606_5 gpc7090 (
      {stage1_60[124], stage1_60[125], stage1_60[126], stage1_60[127], stage1_60[128], stage1_60[129]},
      {stage1_62[88], stage1_62[89], stage1_62[90], stage1_62[91], stage1_62[92], stage1_62[93]},
      {stage2_64[15],stage2_63[44],stage2_62[49],stage2_61[68],stage2_60[89]}
   );
   gpc606_5 gpc7091 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[94], stage1_62[95], stage1_62[96], stage1_62[97], stage1_62[98], stage1_62[99]},
      {stage2_64[16],stage2_63[45],stage2_62[50],stage2_61[69],stage2_60[90]}
   );
   gpc606_5 gpc7092 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[100], stage1_62[101], stage1_62[102], stage1_62[103], stage1_62[104], stage1_62[105]},
      {stage2_64[17],stage2_63[46],stage2_62[51],stage2_61[70],stage2_60[91]}
   );
   gpc606_5 gpc7093 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[106], stage1_62[107], stage1_62[108], stage1_62[109], stage1_62[110], stage1_62[111]},
      {stage2_64[18],stage2_63[47],stage2_62[52],stage2_61[71],stage2_60[92]}
   );
   gpc606_5 gpc7094 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[112], stage1_62[113], stage1_62[114], stage1_62[115], stage1_62[116], stage1_62[117]},
      {stage2_64[19],stage2_63[48],stage2_62[53],stage2_61[72],stage2_60[93]}
   );
   gpc606_5 gpc7095 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[118], stage1_62[119], stage1_62[120], stage1_62[121], stage1_62[122], stage1_62[123]},
      {stage2_64[20],stage2_63[49],stage2_62[54],stage2_61[73],stage2_60[94]}
   );
   gpc615_5 gpc7096 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164]},
      {stage1_61[174]},
      {stage1_62[124], stage1_62[125], stage1_62[126], stage1_62[127], stage1_62[128], stage1_62[129]},
      {stage2_64[21],stage2_63[50],stage2_62[55],stage2_61[74],stage2_60[95]}
   );
   gpc615_5 gpc7097 (
      {stage1_60[165], stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169]},
      {stage1_61[175]},
      {stage1_62[130], stage1_62[131], stage1_62[132], stage1_62[133], stage1_62[134], stage1_62[135]},
      {stage2_64[22],stage2_63[51],stage2_62[56],stage2_61[75],stage2_60[96]}
   );
   gpc615_5 gpc7098 (
      {stage1_60[170], stage1_60[171], stage1_60[172], stage1_60[173], stage1_60[174]},
      {stage1_61[176]},
      {stage1_62[136], stage1_62[137], stage1_62[138], stage1_62[139], stage1_62[140], stage1_62[141]},
      {stage2_64[23],stage2_63[52],stage2_62[57],stage2_61[76],stage2_60[97]}
   );
   gpc615_5 gpc7099 (
      {stage1_60[175], stage1_60[176], stage1_60[177], stage1_60[178], stage1_60[179]},
      {stage1_61[177]},
      {stage1_62[142], stage1_62[143], stage1_62[144], stage1_62[145], stage1_62[146], stage1_62[147]},
      {stage2_64[24],stage2_63[53],stage2_62[58],stage2_61[77],stage2_60[98]}
   );
   gpc615_5 gpc7100 (
      {stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183], stage1_60[184]},
      {stage1_61[178]},
      {stage1_62[148], stage1_62[149], stage1_62[150], stage1_62[151], stage1_62[152], stage1_62[153]},
      {stage2_64[25],stage2_63[54],stage2_62[59],stage2_61[78],stage2_60[99]}
   );
   gpc615_5 gpc7101 (
      {stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188], stage1_60[189]},
      {stage1_61[179]},
      {stage1_62[154], stage1_62[155], stage1_62[156], stage1_62[157], stage1_62[158], stage1_62[159]},
      {stage2_64[26],stage2_63[55],stage2_62[60],stage2_61[79],stage2_60[100]}
   );
   gpc606_5 gpc7102 (
      {stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183], stage1_61[184], stage1_61[185]},
      {stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6]},
      {stage2_65[0],stage2_64[27],stage2_63[56],stage2_62[61],stage2_61[80]}
   );
   gpc606_5 gpc7103 (
      {stage1_61[186], stage1_61[187], stage1_61[188], stage1_61[189], stage1_61[190], stage1_61[191]},
      {stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12]},
      {stage2_65[1],stage2_64[28],stage2_63[57],stage2_62[62],stage2_61[81]}
   );
   gpc606_5 gpc7104 (
      {stage1_61[192], stage1_61[193], stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197]},
      {stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18]},
      {stage2_65[2],stage2_64[29],stage2_63[58],stage2_62[63],stage2_61[82]}
   );
   gpc1163_5 gpc7105 (
      {stage1_62[160], stage1_62[161], stage1_62[162]},
      {stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[3],stage2_64[30],stage2_63[59],stage2_62[64]}
   );
   gpc1163_5 gpc7106 (
      {stage1_62[163], stage1_62[164], stage1_62[165]},
      {stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29], stage1_63[30]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[4],stage2_64[31],stage2_63[60],stage2_62[65]}
   );
   gpc1163_5 gpc7107 (
      {stage1_62[166], stage1_62[167], stage1_62[168]},
      {stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35], stage1_63[36]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[5],stage2_64[32],stage2_63[61],stage2_62[66]}
   );
   gpc1163_5 gpc7108 (
      {stage1_62[169], stage1_62[170], stage1_62[171]},
      {stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41], stage1_63[42]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[6],stage2_64[33],stage2_63[62],stage2_62[67]}
   );
   gpc1163_5 gpc7109 (
      {stage1_62[172], stage1_62[173], stage1_62[174]},
      {stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47], stage1_63[48]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[7],stage2_64[34],stage2_63[63],stage2_62[68]}
   );
   gpc1163_5 gpc7110 (
      {stage1_62[175], stage1_62[176], stage1_62[177]},
      {stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53], stage1_63[54]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[8],stage2_64[35],stage2_63[64],stage2_62[69]}
   );
   gpc1163_5 gpc7111 (
      {stage1_62[178], stage1_62[179], stage1_62[180]},
      {stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59], stage1_63[60]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[9],stage2_64[36],stage2_63[65],stage2_62[70]}
   );
   gpc1163_5 gpc7112 (
      {stage1_62[181], stage1_62[182], stage1_62[183]},
      {stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65], stage1_63[66]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[10],stage2_64[37],stage2_63[66],stage2_62[71]}
   );
   gpc1163_5 gpc7113 (
      {stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71], stage1_63[72]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[11],stage2_64[38],stage2_63[67],stage2_62[72]}
   );
   gpc1163_5 gpc7114 (
      {stage1_62[187], stage1_62[188], stage1_62[189]},
      {stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77], stage1_63[78]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[12],stage2_64[39],stage2_63[68],stage2_62[73]}
   );
   gpc1163_5 gpc7115 (
      {stage1_62[190], stage1_62[191], stage1_62[192]},
      {stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83], stage1_63[84]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[13],stage2_64[40],stage2_63[69],stage2_62[74]}
   );
   gpc1163_5 gpc7116 (
      {stage1_62[193], stage1_62[194], stage1_62[195]},
      {stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89], stage1_63[90]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[14],stage2_64[41],stage2_63[70],stage2_62[75]}
   );
   gpc1163_5 gpc7117 (
      {stage1_62[196], stage1_62[197], stage1_62[198]},
      {stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95], stage1_63[96]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[15],stage2_64[42],stage2_63[71],stage2_62[76]}
   );
   gpc1163_5 gpc7118 (
      {stage1_62[199], stage1_62[200], stage1_62[201]},
      {stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101], stage1_63[102]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[16],stage2_64[43],stage2_63[72],stage2_62[77]}
   );
   gpc1163_5 gpc7119 (
      {stage1_62[202], stage1_62[203], stage1_62[204]},
      {stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107], stage1_63[108]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[17],stage2_64[44],stage2_63[73],stage2_62[78]}
   );
   gpc1163_5 gpc7120 (
      {stage1_62[205], stage1_62[206], stage1_62[207]},
      {stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113], stage1_63[114]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[18],stage2_64[45],stage2_63[74],stage2_62[79]}
   );
   gpc1163_5 gpc7121 (
      {stage1_62[208], stage1_62[209], stage1_62[210]},
      {stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119], stage1_63[120]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[19],stage2_64[46],stage2_63[75],stage2_62[80]}
   );
   gpc1163_5 gpc7122 (
      {stage1_62[211], stage1_62[212], stage1_62[213]},
      {stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125], stage1_63[126]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[20],stage2_64[47],stage2_63[76],stage2_62[81]}
   );
   gpc1163_5 gpc7123 (
      {stage1_62[214], stage1_62[215], stage1_62[216]},
      {stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131], stage1_63[132]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[21],stage2_64[48],stage2_63[77],stage2_62[82]}
   );
   gpc1163_5 gpc7124 (
      {stage1_62[217], stage1_62[218], stage1_62[219]},
      {stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137], stage1_63[138]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[22],stage2_64[49],stage2_63[78],stage2_62[83]}
   );
   gpc1163_5 gpc7125 (
      {stage1_62[220], stage1_62[221], stage1_62[222]},
      {stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143], stage1_63[144]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[23],stage2_64[50],stage2_63[79],stage2_62[84]}
   );
   gpc1163_5 gpc7126 (
      {stage1_62[223], stage1_62[224], stage1_62[225]},
      {stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149], stage1_63[150]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[24],stage2_64[51],stage2_63[80],stage2_62[85]}
   );
   gpc1163_5 gpc7127 (
      {stage1_62[226], stage1_62[227], stage1_62[228]},
      {stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155], stage1_63[156]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[25],stage2_64[52],stage2_63[81],stage2_62[86]}
   );
   gpc1163_5 gpc7128 (
      {stage1_62[229], stage1_62[230], stage1_62[231]},
      {stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161], stage1_63[162]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[26],stage2_64[53],stage2_63[82],stage2_62[87]}
   );
   gpc1163_5 gpc7129 (
      {stage1_62[232], stage1_62[233], stage1_62[234]},
      {stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167], stage1_63[168]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[27],stage2_64[54],stage2_63[83],stage2_62[88]}
   );
   gpc1163_5 gpc7130 (
      {stage1_62[235], stage1_62[236], stage1_62[237]},
      {stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173], stage1_63[174]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[28],stage2_64[55],stage2_63[84],stage2_62[89]}
   );
   gpc1163_5 gpc7131 (
      {stage1_62[238], stage1_62[239], stage1_62[240]},
      {stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179], stage1_63[180]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[29],stage2_64[56],stage2_63[85],stage2_62[90]}
   );
   gpc1163_5 gpc7132 (
      {stage1_62[241], stage1_62[242], stage1_62[243]},
      {stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185], stage1_63[186]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[30],stage2_64[57],stage2_63[86],stage2_62[91]}
   );
   gpc1163_5 gpc7133 (
      {stage1_62[244], stage1_62[245], stage1_62[246]},
      {stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191], stage1_63[192]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[31],stage2_64[58],stage2_63[87],stage2_62[92]}
   );
   gpc1163_5 gpc7134 (
      {stage1_62[247], stage1_62[248], stage1_62[249]},
      {stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197], stage1_63[198]},
      {stage1_64[29]},
      {stage1_65[29]},
      {stage2_66[29],stage2_65[32],stage2_64[59],stage2_63[88],stage2_62[93]}
   );
   gpc1163_5 gpc7135 (
      {stage1_62[250], stage1_62[251], stage1_62[252]},
      {stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203], stage1_63[204]},
      {stage1_64[30]},
      {stage1_65[30]},
      {stage2_66[30],stage2_65[33],stage2_64[60],stage2_63[89],stage2_62[94]}
   );
   gpc1163_5 gpc7136 (
      {stage1_62[253], stage1_62[254], stage1_62[255]},
      {stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209], stage1_63[210]},
      {stage1_64[31]},
      {stage1_65[31]},
      {stage2_66[31],stage2_65[34],stage2_64[61],stage2_63[90],stage2_62[95]}
   );
   gpc1163_5 gpc7137 (
      {stage1_62[256], stage1_62[257], stage1_62[258]},
      {stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215], stage1_63[216]},
      {stage1_64[32]},
      {stage1_65[32]},
      {stage2_66[32],stage2_65[35],stage2_64[62],stage2_63[91],stage2_62[96]}
   );
   gpc1163_5 gpc7138 (
      {stage1_62[259], stage1_62[260], stage1_62[261]},
      {stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221], stage1_63[222]},
      {stage1_64[33]},
      {stage1_65[33]},
      {stage2_66[33],stage2_65[36],stage2_64[63],stage2_63[92],stage2_62[97]}
   );
   gpc1163_5 gpc7139 (
      {stage1_62[262], stage1_62[263], stage1_62[264]},
      {stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227], stage1_63[228]},
      {stage1_64[34]},
      {stage1_65[34]},
      {stage2_66[34],stage2_65[37],stage2_64[64],stage2_63[93],stage2_62[98]}
   );
   gpc1163_5 gpc7140 (
      {stage1_62[265], stage1_62[266], stage1_62[267]},
      {stage1_63[229], stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[35]},
      {stage1_65[35]},
      {stage2_66[35],stage2_65[38],stage2_64[65],stage2_63[94],stage2_62[99]}
   );
   gpc1163_5 gpc7141 (
      {stage1_62[268], stage1_62[269], stage1_62[270]},
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239], stage1_63[240]},
      {stage1_64[36]},
      {stage1_65[36]},
      {stage2_66[36],stage2_65[39],stage2_64[66],stage2_63[95],stage2_62[100]}
   );
   gpc1163_5 gpc7142 (
      {stage1_62[271], stage1_62[272], stage1_62[273]},
      {stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_64[37]},
      {stage1_65[37]},
      {stage2_66[37],stage2_65[40],stage2_64[67],stage2_63[96],stage2_62[101]}
   );
   gpc1163_5 gpc7143 (
      {stage1_62[274], stage1_62[275], stage1_62[276]},
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252]},
      {stage1_64[38]},
      {stage1_65[38]},
      {stage2_66[38],stage2_65[41],stage2_64[68],stage2_63[97],stage2_62[102]}
   );
   gpc1163_5 gpc7144 (
      {stage1_62[277], stage1_62[278], stage1_62[279]},
      {stage1_63[253], stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258]},
      {stage1_64[39]},
      {stage1_65[39]},
      {stage2_66[39],stage2_65[42],stage2_64[69],stage2_63[98],stage2_62[103]}
   );
   gpc1163_5 gpc7145 (
      {stage1_62[280], stage1_62[281], stage1_62[282]},
      {stage1_63[259], stage1_63[260], stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264]},
      {stage1_64[40]},
      {stage1_65[40]},
      {stage2_66[40],stage2_65[43],stage2_64[70],stage2_63[99],stage2_62[104]}
   );
   gpc1163_5 gpc7146 (
      {stage1_62[283], stage1_62[284], stage1_62[285]},
      {stage1_63[265], stage1_63[266], stage1_63[267], stage1_63[268], stage1_63[269], stage1_63[270]},
      {stage1_64[41]},
      {stage1_65[41]},
      {stage2_66[41],stage2_65[44],stage2_64[71],stage2_63[100],stage2_62[105]}
   );
   gpc1163_5 gpc7147 (
      {stage1_62[286], stage1_62[287], stage1_62[288]},
      {stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274], stage1_63[275], stage1_63[276]},
      {stage1_64[42]},
      {stage1_65[42]},
      {stage2_66[42],stage2_65[45],stage2_64[72],stage2_63[101],stage2_62[106]}
   );
   gpc1163_5 gpc7148 (
      {stage1_62[289], stage1_62[290], stage1_62[291]},
      {stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281], stage1_63[282]},
      {stage1_64[43]},
      {stage1_65[43]},
      {stage2_66[43],stage2_65[46],stage2_64[73],stage2_63[102],stage2_62[107]}
   );
   gpc1163_5 gpc7149 (
      {stage1_62[292], stage1_62[293], stage1_62[294]},
      {stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_64[44]},
      {stage1_65[44]},
      {stage2_66[44],stage2_65[47],stage2_64[74],stage2_63[103],stage2_62[108]}
   );
   gpc1163_5 gpc7150 (
      {stage1_62[295], stage1_62[296], stage1_62[297]},
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294]},
      {stage1_64[45]},
      {stage1_65[45]},
      {stage2_66[45],stage2_65[48],stage2_64[75],stage2_63[104],stage2_62[109]}
   );
   gpc606_5 gpc7151 (
      {stage1_62[298], stage1_62[299], stage1_62[300], stage1_62[301], stage1_62[302], stage1_62[303]},
      {stage1_64[46], stage1_64[47], stage1_64[48], stage1_64[49], stage1_64[50], stage1_64[51]},
      {stage2_66[46],stage2_65[49],stage2_64[76],stage2_63[105],stage2_62[110]}
   );
   gpc606_5 gpc7152 (
      {stage1_62[304], stage1_62[305], stage1_62[306], stage1_62[307], stage1_62[308], stage1_62[309]},
      {stage1_64[52], stage1_64[53], stage1_64[54], stage1_64[55], stage1_64[56], stage1_64[57]},
      {stage2_66[47],stage2_65[50],stage2_64[77],stage2_63[106],stage2_62[111]}
   );
   gpc606_5 gpc7153 (
      {stage1_62[310], stage1_62[311], stage1_62[312], stage1_62[313], stage1_62[314], stage1_62[315]},
      {stage1_64[58], stage1_64[59], stage1_64[60], stage1_64[61], stage1_64[62], stage1_64[63]},
      {stage2_66[48],stage2_65[51],stage2_64[78],stage2_63[107],stage2_62[112]}
   );
   gpc606_5 gpc7154 (
      {stage1_62[316], stage1_62[317], stage1_62[318], stage1_62[319], stage1_62[320], stage1_62[321]},
      {stage1_64[64], stage1_64[65], stage1_64[66], stage1_64[67], stage1_64[68], stage1_64[69]},
      {stage2_66[49],stage2_65[52],stage2_64[79],stage2_63[108],stage2_62[113]}
   );
   gpc606_5 gpc7155 (
      {stage1_62[322], stage1_62[323], stage1_62[324], stage1_62[325], stage1_62[326], stage1_62[327]},
      {stage1_64[70], stage1_64[71], stage1_64[72], stage1_64[73], stage1_64[74], stage1_64[75]},
      {stage2_66[50],stage2_65[53],stage2_64[80],stage2_63[109],stage2_62[114]}
   );
   gpc606_5 gpc7156 (
      {stage1_62[328], stage1_62[329], stage1_62[330], stage1_62[331], stage1_62[332], stage1_62[333]},
      {stage1_64[76], stage1_64[77], stage1_64[78], stage1_64[79], stage1_64[80], stage1_64[81]},
      {stage2_66[51],stage2_65[54],stage2_64[81],stage2_63[110],stage2_62[115]}
   );
   gpc606_5 gpc7157 (
      {stage1_62[334], stage1_62[335], stage1_62[336], stage1_62[337], stage1_62[338], stage1_62[339]},
      {stage1_64[82], stage1_64[83], stage1_64[84], stage1_64[85], stage1_64[86], stage1_64[87]},
      {stage2_66[52],stage2_65[55],stage2_64[82],stage2_63[111],stage2_62[116]}
   );
   gpc606_5 gpc7158 (
      {stage1_62[340], stage1_62[341], stage1_62[342], stage1_62[343], stage1_62[344], stage1_62[345]},
      {stage1_64[88], stage1_64[89], stage1_64[90], stage1_64[91], stage1_64[92], stage1_64[93]},
      {stage2_66[53],stage2_65[56],stage2_64[83],stage2_63[112],stage2_62[117]}
   );
   gpc1_1 gpc7159 (
      {stage1_0[112]},
      {stage2_0[27]}
   );
   gpc1_1 gpc7160 (
      {stage1_0[113]},
      {stage2_0[28]}
   );
   gpc1_1 gpc7161 (
      {stage1_0[114]},
      {stage2_0[29]}
   );
   gpc1_1 gpc7162 (
      {stage1_0[115]},
      {stage2_0[30]}
   );
   gpc1_1 gpc7163 (
      {stage1_0[116]},
      {stage2_0[31]}
   );
   gpc1_1 gpc7164 (
      {stage1_0[117]},
      {stage2_0[32]}
   );
   gpc1_1 gpc7165 (
      {stage1_0[118]},
      {stage2_0[33]}
   );
   gpc1_1 gpc7166 (
      {stage1_2[208]},
      {stage2_2[60]}
   );
   gpc1_1 gpc7167 (
      {stage1_2[209]},
      {stage2_2[61]}
   );
   gpc1_1 gpc7168 (
      {stage1_2[210]},
      {stage2_2[62]}
   );
   gpc1_1 gpc7169 (
      {stage1_2[211]},
      {stage2_2[63]}
   );
   gpc1_1 gpc7170 (
      {stage1_2[212]},
      {stage2_2[64]}
   );
   gpc1_1 gpc7171 (
      {stage1_2[213]},
      {stage2_2[65]}
   );
   gpc1_1 gpc7172 (
      {stage1_2[214]},
      {stage2_2[66]}
   );
   gpc1_1 gpc7173 (
      {stage1_2[215]},
      {stage2_2[67]}
   );
   gpc1_1 gpc7174 (
      {stage1_2[216]},
      {stage2_2[68]}
   );
   gpc1_1 gpc7175 (
      {stage1_2[217]},
      {stage2_2[69]}
   );
   gpc1_1 gpc7176 (
      {stage1_2[218]},
      {stage2_2[70]}
   );
   gpc1_1 gpc7177 (
      {stage1_2[219]},
      {stage2_2[71]}
   );
   gpc1_1 gpc7178 (
      {stage1_2[220]},
      {stage2_2[72]}
   );
   gpc1_1 gpc7179 (
      {stage1_3[139]},
      {stage2_3[71]}
   );
   gpc1_1 gpc7180 (
      {stage1_3[140]},
      {stage2_3[72]}
   );
   gpc1_1 gpc7181 (
      {stage1_3[141]},
      {stage2_3[73]}
   );
   gpc1_1 gpc7182 (
      {stage1_3[142]},
      {stage2_3[74]}
   );
   gpc1_1 gpc7183 (
      {stage1_3[143]},
      {stage2_3[75]}
   );
   gpc1_1 gpc7184 (
      {stage1_3[144]},
      {stage2_3[76]}
   );
   gpc1_1 gpc7185 (
      {stage1_3[145]},
      {stage2_3[77]}
   );
   gpc1_1 gpc7186 (
      {stage1_3[146]},
      {stage2_3[78]}
   );
   gpc1_1 gpc7187 (
      {stage1_3[147]},
      {stage2_3[79]}
   );
   gpc1_1 gpc7188 (
      {stage1_3[148]},
      {stage2_3[80]}
   );
   gpc1_1 gpc7189 (
      {stage1_3[149]},
      {stage2_3[81]}
   );
   gpc1_1 gpc7190 (
      {stage1_3[150]},
      {stage2_3[82]}
   );
   gpc1_1 gpc7191 (
      {stage1_3[151]},
      {stage2_3[83]}
   );
   gpc1_1 gpc7192 (
      {stage1_3[152]},
      {stage2_3[84]}
   );
   gpc1_1 gpc7193 (
      {stage1_3[153]},
      {stage2_3[85]}
   );
   gpc1_1 gpc7194 (
      {stage1_3[154]},
      {stage2_3[86]}
   );
   gpc1_1 gpc7195 (
      {stage1_3[155]},
      {stage2_3[87]}
   );
   gpc1_1 gpc7196 (
      {stage1_3[156]},
      {stage2_3[88]}
   );
   gpc1_1 gpc7197 (
      {stage1_3[157]},
      {stage2_3[89]}
   );
   gpc1_1 gpc7198 (
      {stage1_3[158]},
      {stage2_3[90]}
   );
   gpc1_1 gpc7199 (
      {stage1_3[159]},
      {stage2_3[91]}
   );
   gpc1_1 gpc7200 (
      {stage1_3[160]},
      {stage2_3[92]}
   );
   gpc1_1 gpc7201 (
      {stage1_3[161]},
      {stage2_3[93]}
   );
   gpc1_1 gpc7202 (
      {stage1_3[162]},
      {stage2_3[94]}
   );
   gpc1_1 gpc7203 (
      {stage1_3[163]},
      {stage2_3[95]}
   );
   gpc1_1 gpc7204 (
      {stage1_3[164]},
      {stage2_3[96]}
   );
   gpc1_1 gpc7205 (
      {stage1_3[165]},
      {stage2_3[97]}
   );
   gpc1_1 gpc7206 (
      {stage1_3[166]},
      {stage2_3[98]}
   );
   gpc1_1 gpc7207 (
      {stage1_3[167]},
      {stage2_3[99]}
   );
   gpc1_1 gpc7208 (
      {stage1_3[168]},
      {stage2_3[100]}
   );
   gpc1_1 gpc7209 (
      {stage1_3[169]},
      {stage2_3[101]}
   );
   gpc1_1 gpc7210 (
      {stage1_3[170]},
      {stage2_3[102]}
   );
   gpc1_1 gpc7211 (
      {stage1_3[171]},
      {stage2_3[103]}
   );
   gpc1_1 gpc7212 (
      {stage1_3[172]},
      {stage2_3[104]}
   );
   gpc1_1 gpc7213 (
      {stage1_3[173]},
      {stage2_3[105]}
   );
   gpc1_1 gpc7214 (
      {stage1_3[174]},
      {stage2_3[106]}
   );
   gpc1_1 gpc7215 (
      {stage1_3[175]},
      {stage2_3[107]}
   );
   gpc1_1 gpc7216 (
      {stage1_3[176]},
      {stage2_3[108]}
   );
   gpc1_1 gpc7217 (
      {stage1_3[177]},
      {stage2_3[109]}
   );
   gpc1_1 gpc7218 (
      {stage1_3[178]},
      {stage2_3[110]}
   );
   gpc1_1 gpc7219 (
      {stage1_3[179]},
      {stage2_3[111]}
   );
   gpc1_1 gpc7220 (
      {stage1_3[180]},
      {stage2_3[112]}
   );
   gpc1_1 gpc7221 (
      {stage1_3[181]},
      {stage2_3[113]}
   );
   gpc1_1 gpc7222 (
      {stage1_3[182]},
      {stage2_3[114]}
   );
   gpc1_1 gpc7223 (
      {stage1_3[183]},
      {stage2_3[115]}
   );
   gpc1_1 gpc7224 (
      {stage1_3[184]},
      {stage2_3[116]}
   );
   gpc1_1 gpc7225 (
      {stage1_3[185]},
      {stage2_3[117]}
   );
   gpc1_1 gpc7226 (
      {stage1_3[186]},
      {stage2_3[118]}
   );
   gpc1_1 gpc7227 (
      {stage1_3[187]},
      {stage2_3[119]}
   );
   gpc1_1 gpc7228 (
      {stage1_3[188]},
      {stage2_3[120]}
   );
   gpc1_1 gpc7229 (
      {stage1_3[189]},
      {stage2_3[121]}
   );
   gpc1_1 gpc7230 (
      {stage1_3[190]},
      {stage2_3[122]}
   );
   gpc1_1 gpc7231 (
      {stage1_3[191]},
      {stage2_3[123]}
   );
   gpc1_1 gpc7232 (
      {stage1_3[192]},
      {stage2_3[124]}
   );
   gpc1_1 gpc7233 (
      {stage1_3[193]},
      {stage2_3[125]}
   );
   gpc1_1 gpc7234 (
      {stage1_3[194]},
      {stage2_3[126]}
   );
   gpc1_1 gpc7235 (
      {stage1_3[195]},
      {stage2_3[127]}
   );
   gpc1_1 gpc7236 (
      {stage1_3[196]},
      {stage2_3[128]}
   );
   gpc1_1 gpc7237 (
      {stage1_3[197]},
      {stage2_3[129]}
   );
   gpc1_1 gpc7238 (
      {stage1_3[198]},
      {stage2_3[130]}
   );
   gpc1_1 gpc7239 (
      {stage1_3[199]},
      {stage2_3[131]}
   );
   gpc1_1 gpc7240 (
      {stage1_3[200]},
      {stage2_3[132]}
   );
   gpc1_1 gpc7241 (
      {stage1_3[201]},
      {stage2_3[133]}
   );
   gpc1_1 gpc7242 (
      {stage1_3[202]},
      {stage2_3[134]}
   );
   gpc1_1 gpc7243 (
      {stage1_3[203]},
      {stage2_3[135]}
   );
   gpc1_1 gpc7244 (
      {stage1_3[204]},
      {stage2_3[136]}
   );
   gpc1_1 gpc7245 (
      {stage1_3[205]},
      {stage2_3[137]}
   );
   gpc1_1 gpc7246 (
      {stage1_3[206]},
      {stage2_3[138]}
   );
   gpc1_1 gpc7247 (
      {stage1_3[207]},
      {stage2_3[139]}
   );
   gpc1_1 gpc7248 (
      {stage1_3[208]},
      {stage2_3[140]}
   );
   gpc1_1 gpc7249 (
      {stage1_3[209]},
      {stage2_3[141]}
   );
   gpc1_1 gpc7250 (
      {stage1_3[210]},
      {stage2_3[142]}
   );
   gpc1_1 gpc7251 (
      {stage1_3[211]},
      {stage2_3[143]}
   );
   gpc1_1 gpc7252 (
      {stage1_3[212]},
      {stage2_3[144]}
   );
   gpc1_1 gpc7253 (
      {stage1_3[213]},
      {stage2_3[145]}
   );
   gpc1_1 gpc7254 (
      {stage1_3[214]},
      {stage2_3[146]}
   );
   gpc1_1 gpc7255 (
      {stage1_3[215]},
      {stage2_3[147]}
   );
   gpc1_1 gpc7256 (
      {stage1_3[216]},
      {stage2_3[148]}
   );
   gpc1_1 gpc7257 (
      {stage1_3[217]},
      {stage2_3[149]}
   );
   gpc1_1 gpc7258 (
      {stage1_3[218]},
      {stage2_3[150]}
   );
   gpc1_1 gpc7259 (
      {stage1_3[219]},
      {stage2_3[151]}
   );
   gpc1_1 gpc7260 (
      {stage1_3[220]},
      {stage2_3[152]}
   );
   gpc1_1 gpc7261 (
      {stage1_3[221]},
      {stage2_3[153]}
   );
   gpc1_1 gpc7262 (
      {stage1_3[222]},
      {stage2_3[154]}
   );
   gpc1_1 gpc7263 (
      {stage1_3[223]},
      {stage2_3[155]}
   );
   gpc1_1 gpc7264 (
      {stage1_3[224]},
      {stage2_3[156]}
   );
   gpc1_1 gpc7265 (
      {stage1_3[225]},
      {stage2_3[157]}
   );
   gpc1_1 gpc7266 (
      {stage1_3[226]},
      {stage2_3[158]}
   );
   gpc1_1 gpc7267 (
      {stage1_3[227]},
      {stage2_3[159]}
   );
   gpc1_1 gpc7268 (
      {stage1_3[228]},
      {stage2_3[160]}
   );
   gpc1_1 gpc7269 (
      {stage1_3[229]},
      {stage2_3[161]}
   );
   gpc1_1 gpc7270 (
      {stage1_3[230]},
      {stage2_3[162]}
   );
   gpc1_1 gpc7271 (
      {stage1_3[231]},
      {stage2_3[163]}
   );
   gpc1_1 gpc7272 (
      {stage1_3[232]},
      {stage2_3[164]}
   );
   gpc1_1 gpc7273 (
      {stage1_3[233]},
      {stage2_3[165]}
   );
   gpc1_1 gpc7274 (
      {stage1_3[234]},
      {stage2_3[166]}
   );
   gpc1_1 gpc7275 (
      {stage1_3[235]},
      {stage2_3[167]}
   );
   gpc1_1 gpc7276 (
      {stage1_3[236]},
      {stage2_3[168]}
   );
   gpc1_1 gpc7277 (
      {stage1_3[237]},
      {stage2_3[169]}
   );
   gpc1_1 gpc7278 (
      {stage1_3[238]},
      {stage2_3[170]}
   );
   gpc1_1 gpc7279 (
      {stage1_3[239]},
      {stage2_3[171]}
   );
   gpc1_1 gpc7280 (
      {stage1_3[240]},
      {stage2_3[172]}
   );
   gpc1_1 gpc7281 (
      {stage1_3[241]},
      {stage2_3[173]}
   );
   gpc1_1 gpc7282 (
      {stage1_3[242]},
      {stage2_3[174]}
   );
   gpc1_1 gpc7283 (
      {stage1_3[243]},
      {stage2_3[175]}
   );
   gpc1_1 gpc7284 (
      {stage1_3[244]},
      {stage2_3[176]}
   );
   gpc1_1 gpc7285 (
      {stage1_3[245]},
      {stage2_3[177]}
   );
   gpc1_1 gpc7286 (
      {stage1_3[246]},
      {stage2_3[178]}
   );
   gpc1_1 gpc7287 (
      {stage1_3[247]},
      {stage2_3[179]}
   );
   gpc1_1 gpc7288 (
      {stage1_3[248]},
      {stage2_3[180]}
   );
   gpc1_1 gpc7289 (
      {stage1_3[249]},
      {stage2_3[181]}
   );
   gpc1_1 gpc7290 (
      {stage1_3[250]},
      {stage2_3[182]}
   );
   gpc1_1 gpc7291 (
      {stage1_3[251]},
      {stage2_3[183]}
   );
   gpc1_1 gpc7292 (
      {stage1_3[252]},
      {stage2_3[184]}
   );
   gpc1_1 gpc7293 (
      {stage1_3[253]},
      {stage2_3[185]}
   );
   gpc1_1 gpc7294 (
      {stage1_3[254]},
      {stage2_3[186]}
   );
   gpc1_1 gpc7295 (
      {stage1_3[255]},
      {stage2_3[187]}
   );
   gpc1_1 gpc7296 (
      {stage1_3[256]},
      {stage2_3[188]}
   );
   gpc1_1 gpc7297 (
      {stage1_3[257]},
      {stage2_3[189]}
   );
   gpc1_1 gpc7298 (
      {stage1_3[258]},
      {stage2_3[190]}
   );
   gpc1_1 gpc7299 (
      {stage1_3[259]},
      {stage2_3[191]}
   );
   gpc1_1 gpc7300 (
      {stage1_3[260]},
      {stage2_3[192]}
   );
   gpc1_1 gpc7301 (
      {stage1_3[261]},
      {stage2_3[193]}
   );
   gpc1_1 gpc7302 (
      {stage1_3[262]},
      {stage2_3[194]}
   );
   gpc1_1 gpc7303 (
      {stage1_3[263]},
      {stage2_3[195]}
   );
   gpc1_1 gpc7304 (
      {stage1_3[264]},
      {stage2_3[196]}
   );
   gpc1_1 gpc7305 (
      {stage1_3[265]},
      {stage2_3[197]}
   );
   gpc1_1 gpc7306 (
      {stage1_3[266]},
      {stage2_3[198]}
   );
   gpc1_1 gpc7307 (
      {stage1_3[267]},
      {stage2_3[199]}
   );
   gpc1_1 gpc7308 (
      {stage1_3[268]},
      {stage2_3[200]}
   );
   gpc1_1 gpc7309 (
      {stage1_3[269]},
      {stage2_3[201]}
   );
   gpc1_1 gpc7310 (
      {stage1_3[270]},
      {stage2_3[202]}
   );
   gpc1_1 gpc7311 (
      {stage1_3[271]},
      {stage2_3[203]}
   );
   gpc1_1 gpc7312 (
      {stage1_3[272]},
      {stage2_3[204]}
   );
   gpc1_1 gpc7313 (
      {stage1_3[273]},
      {stage2_3[205]}
   );
   gpc1_1 gpc7314 (
      {stage1_3[274]},
      {stage2_3[206]}
   );
   gpc1_1 gpc7315 (
      {stage1_3[275]},
      {stage2_3[207]}
   );
   gpc1_1 gpc7316 (
      {stage1_3[276]},
      {stage2_3[208]}
   );
   gpc1_1 gpc7317 (
      {stage1_3[277]},
      {stage2_3[209]}
   );
   gpc1_1 gpc7318 (
      {stage1_3[278]},
      {stage2_3[210]}
   );
   gpc1_1 gpc7319 (
      {stage1_3[279]},
      {stage2_3[211]}
   );
   gpc1_1 gpc7320 (
      {stage1_3[280]},
      {stage2_3[212]}
   );
   gpc1_1 gpc7321 (
      {stage1_3[281]},
      {stage2_3[213]}
   );
   gpc1_1 gpc7322 (
      {stage1_3[282]},
      {stage2_3[214]}
   );
   gpc1_1 gpc7323 (
      {stage1_3[283]},
      {stage2_3[215]}
   );
   gpc1_1 gpc7324 (
      {stage1_3[284]},
      {stage2_3[216]}
   );
   gpc1_1 gpc7325 (
      {stage1_3[285]},
      {stage2_3[217]}
   );
   gpc1_1 gpc7326 (
      {stage1_3[286]},
      {stage2_3[218]}
   );
   gpc1_1 gpc7327 (
      {stage1_3[287]},
      {stage2_3[219]}
   );
   gpc1_1 gpc7328 (
      {stage1_3[288]},
      {stage2_3[220]}
   );
   gpc1_1 gpc7329 (
      {stage1_3[289]},
      {stage2_3[221]}
   );
   gpc1_1 gpc7330 (
      {stage1_3[290]},
      {stage2_3[222]}
   );
   gpc1_1 gpc7331 (
      {stage1_3[291]},
      {stage2_3[223]}
   );
   gpc1_1 gpc7332 (
      {stage1_3[292]},
      {stage2_3[224]}
   );
   gpc1_1 gpc7333 (
      {stage1_3[293]},
      {stage2_3[225]}
   );
   gpc1_1 gpc7334 (
      {stage1_3[294]},
      {stage2_3[226]}
   );
   gpc1_1 gpc7335 (
      {stage1_3[295]},
      {stage2_3[227]}
   );
   gpc1_1 gpc7336 (
      {stage1_3[296]},
      {stage2_3[228]}
   );
   gpc1_1 gpc7337 (
      {stage1_3[297]},
      {stage2_3[229]}
   );
   gpc1_1 gpc7338 (
      {stage1_3[298]},
      {stage2_3[230]}
   );
   gpc1_1 gpc7339 (
      {stage1_3[299]},
      {stage2_3[231]}
   );
   gpc1_1 gpc7340 (
      {stage1_3[300]},
      {stage2_3[232]}
   );
   gpc1_1 gpc7341 (
      {stage1_3[301]},
      {stage2_3[233]}
   );
   gpc1_1 gpc7342 (
      {stage1_3[302]},
      {stage2_3[234]}
   );
   gpc1_1 gpc7343 (
      {stage1_3[303]},
      {stage2_3[235]}
   );
   gpc1_1 gpc7344 (
      {stage1_3[304]},
      {stage2_3[236]}
   );
   gpc1_1 gpc7345 (
      {stage1_3[305]},
      {stage2_3[237]}
   );
   gpc1_1 gpc7346 (
      {stage1_3[306]},
      {stage2_3[238]}
   );
   gpc1_1 gpc7347 (
      {stage1_3[307]},
      {stage2_3[239]}
   );
   gpc1_1 gpc7348 (
      {stage1_3[308]},
      {stage2_3[240]}
   );
   gpc1_1 gpc7349 (
      {stage1_3[309]},
      {stage2_3[241]}
   );
   gpc1_1 gpc7350 (
      {stage1_3[310]},
      {stage2_3[242]}
   );
   gpc1_1 gpc7351 (
      {stage1_3[311]},
      {stage2_3[243]}
   );
   gpc1_1 gpc7352 (
      {stage1_3[312]},
      {stage2_3[244]}
   );
   gpc1_1 gpc7353 (
      {stage1_3[313]},
      {stage2_3[245]}
   );
   gpc1_1 gpc7354 (
      {stage1_3[314]},
      {stage2_3[246]}
   );
   gpc1_1 gpc7355 (
      {stage1_3[315]},
      {stage2_3[247]}
   );
   gpc1_1 gpc7356 (
      {stage1_3[316]},
      {stage2_3[248]}
   );
   gpc1_1 gpc7357 (
      {stage1_3[317]},
      {stage2_3[249]}
   );
   gpc1_1 gpc7358 (
      {stage1_3[318]},
      {stage2_3[250]}
   );
   gpc1_1 gpc7359 (
      {stage1_3[319]},
      {stage2_3[251]}
   );
   gpc1_1 gpc7360 (
      {stage1_3[320]},
      {stage2_3[252]}
   );
   gpc1_1 gpc7361 (
      {stage1_3[321]},
      {stage2_3[253]}
   );
   gpc1_1 gpc7362 (
      {stage1_4[247]},
      {stage2_4[89]}
   );
   gpc1_1 gpc7363 (
      {stage1_4[248]},
      {stage2_4[90]}
   );
   gpc1_1 gpc7364 (
      {stage1_4[249]},
      {stage2_4[91]}
   );
   gpc1_1 gpc7365 (
      {stage1_4[250]},
      {stage2_4[92]}
   );
   gpc1_1 gpc7366 (
      {stage1_5[188]},
      {stage2_5[83]}
   );
   gpc1_1 gpc7367 (
      {stage1_5[189]},
      {stage2_5[84]}
   );
   gpc1_1 gpc7368 (
      {stage1_5[190]},
      {stage2_5[85]}
   );
   gpc1_1 gpc7369 (
      {stage1_5[191]},
      {stage2_5[86]}
   );
   gpc1_1 gpc7370 (
      {stage1_5[192]},
      {stage2_5[87]}
   );
   gpc1_1 gpc7371 (
      {stage1_5[193]},
      {stage2_5[88]}
   );
   gpc1_1 gpc7372 (
      {stage1_5[194]},
      {stage2_5[89]}
   );
   gpc1_1 gpc7373 (
      {stage1_5[195]},
      {stage2_5[90]}
   );
   gpc1_1 gpc7374 (
      {stage1_5[196]},
      {stage2_5[91]}
   );
   gpc1_1 gpc7375 (
      {stage1_5[197]},
      {stage2_5[92]}
   );
   gpc1_1 gpc7376 (
      {stage1_5[198]},
      {stage2_5[93]}
   );
   gpc1_1 gpc7377 (
      {stage1_5[199]},
      {stage2_5[94]}
   );
   gpc1_1 gpc7378 (
      {stage1_5[200]},
      {stage2_5[95]}
   );
   gpc1_1 gpc7379 (
      {stage1_5[201]},
      {stage2_5[96]}
   );
   gpc1_1 gpc7380 (
      {stage1_5[202]},
      {stage2_5[97]}
   );
   gpc1_1 gpc7381 (
      {stage1_5[203]},
      {stage2_5[98]}
   );
   gpc1_1 gpc7382 (
      {stage1_5[204]},
      {stage2_5[99]}
   );
   gpc1_1 gpc7383 (
      {stage1_5[205]},
      {stage2_5[100]}
   );
   gpc1_1 gpc7384 (
      {stage1_5[206]},
      {stage2_5[101]}
   );
   gpc1_1 gpc7385 (
      {stage1_5[207]},
      {stage2_5[102]}
   );
   gpc1_1 gpc7386 (
      {stage1_5[208]},
      {stage2_5[103]}
   );
   gpc1_1 gpc7387 (
      {stage1_5[209]},
      {stage2_5[104]}
   );
   gpc1_1 gpc7388 (
      {stage1_5[210]},
      {stage2_5[105]}
   );
   gpc1_1 gpc7389 (
      {stage1_5[211]},
      {stage2_5[106]}
   );
   gpc1_1 gpc7390 (
      {stage1_5[212]},
      {stage2_5[107]}
   );
   gpc1_1 gpc7391 (
      {stage1_5[213]},
      {stage2_5[108]}
   );
   gpc1_1 gpc7392 (
      {stage1_5[214]},
      {stage2_5[109]}
   );
   gpc1_1 gpc7393 (
      {stage1_5[215]},
      {stage2_5[110]}
   );
   gpc1_1 gpc7394 (
      {stage1_5[216]},
      {stage2_5[111]}
   );
   gpc1_1 gpc7395 (
      {stage1_6[135]},
      {stage2_6[76]}
   );
   gpc1_1 gpc7396 (
      {stage1_6[136]},
      {stage2_6[77]}
   );
   gpc1_1 gpc7397 (
      {stage1_6[137]},
      {stage2_6[78]}
   );
   gpc1_1 gpc7398 (
      {stage1_6[138]},
      {stage2_6[79]}
   );
   gpc1_1 gpc7399 (
      {stage1_6[139]},
      {stage2_6[80]}
   );
   gpc1_1 gpc7400 (
      {stage1_6[140]},
      {stage2_6[81]}
   );
   gpc1_1 gpc7401 (
      {stage1_6[141]},
      {stage2_6[82]}
   );
   gpc1_1 gpc7402 (
      {stage1_6[142]},
      {stage2_6[83]}
   );
   gpc1_1 gpc7403 (
      {stage1_6[143]},
      {stage2_6[84]}
   );
   gpc1_1 gpc7404 (
      {stage1_6[144]},
      {stage2_6[85]}
   );
   gpc1_1 gpc7405 (
      {stage1_6[145]},
      {stage2_6[86]}
   );
   gpc1_1 gpc7406 (
      {stage1_6[146]},
      {stage2_6[87]}
   );
   gpc1_1 gpc7407 (
      {stage1_6[147]},
      {stage2_6[88]}
   );
   gpc1_1 gpc7408 (
      {stage1_6[148]},
      {stage2_6[89]}
   );
   gpc1_1 gpc7409 (
      {stage1_6[149]},
      {stage2_6[90]}
   );
   gpc1_1 gpc7410 (
      {stage1_6[150]},
      {stage2_6[91]}
   );
   gpc1_1 gpc7411 (
      {stage1_6[151]},
      {stage2_6[92]}
   );
   gpc1_1 gpc7412 (
      {stage1_6[152]},
      {stage2_6[93]}
   );
   gpc1_1 gpc7413 (
      {stage1_6[153]},
      {stage2_6[94]}
   );
   gpc1_1 gpc7414 (
      {stage1_6[154]},
      {stage2_6[95]}
   );
   gpc1_1 gpc7415 (
      {stage1_6[155]},
      {stage2_6[96]}
   );
   gpc1_1 gpc7416 (
      {stage1_6[156]},
      {stage2_6[97]}
   );
   gpc1_1 gpc7417 (
      {stage1_6[157]},
      {stage2_6[98]}
   );
   gpc1_1 gpc7418 (
      {stage1_6[158]},
      {stage2_6[99]}
   );
   gpc1_1 gpc7419 (
      {stage1_6[159]},
      {stage2_6[100]}
   );
   gpc1_1 gpc7420 (
      {stage1_6[160]},
      {stage2_6[101]}
   );
   gpc1_1 gpc7421 (
      {stage1_6[161]},
      {stage2_6[102]}
   );
   gpc1_1 gpc7422 (
      {stage1_6[162]},
      {stage2_6[103]}
   );
   gpc1_1 gpc7423 (
      {stage1_6[163]},
      {stage2_6[104]}
   );
   gpc1_1 gpc7424 (
      {stage1_6[164]},
      {stage2_6[105]}
   );
   gpc1_1 gpc7425 (
      {stage1_6[165]},
      {stage2_6[106]}
   );
   gpc1_1 gpc7426 (
      {stage1_6[166]},
      {stage2_6[107]}
   );
   gpc1_1 gpc7427 (
      {stage1_6[167]},
      {stage2_6[108]}
   );
   gpc1_1 gpc7428 (
      {stage1_6[168]},
      {stage2_6[109]}
   );
   gpc1_1 gpc7429 (
      {stage1_6[169]},
      {stage2_6[110]}
   );
   gpc1_1 gpc7430 (
      {stage1_6[170]},
      {stage2_6[111]}
   );
   gpc1_1 gpc7431 (
      {stage1_6[171]},
      {stage2_6[112]}
   );
   gpc1_1 gpc7432 (
      {stage1_6[172]},
      {stage2_6[113]}
   );
   gpc1_1 gpc7433 (
      {stage1_6[173]},
      {stage2_6[114]}
   );
   gpc1_1 gpc7434 (
      {stage1_6[174]},
      {stage2_6[115]}
   );
   gpc1_1 gpc7435 (
      {stage1_6[175]},
      {stage2_6[116]}
   );
   gpc1_1 gpc7436 (
      {stage1_6[176]},
      {stage2_6[117]}
   );
   gpc1_1 gpc7437 (
      {stage1_6[177]},
      {stage2_6[118]}
   );
   gpc1_1 gpc7438 (
      {stage1_6[178]},
      {stage2_6[119]}
   );
   gpc1_1 gpc7439 (
      {stage1_6[179]},
      {stage2_6[120]}
   );
   gpc1_1 gpc7440 (
      {stage1_8[168]},
      {stage2_8[102]}
   );
   gpc1_1 gpc7441 (
      {stage1_8[169]},
      {stage2_8[103]}
   );
   gpc1_1 gpc7442 (
      {stage1_8[170]},
      {stage2_8[104]}
   );
   gpc1_1 gpc7443 (
      {stage1_8[171]},
      {stage2_8[105]}
   );
   gpc1_1 gpc7444 (
      {stage1_8[172]},
      {stage2_8[106]}
   );
   gpc1_1 gpc7445 (
      {stage1_8[173]},
      {stage2_8[107]}
   );
   gpc1_1 gpc7446 (
      {stage1_8[174]},
      {stage2_8[108]}
   );
   gpc1_1 gpc7447 (
      {stage1_8[175]},
      {stage2_8[109]}
   );
   gpc1_1 gpc7448 (
      {stage1_8[176]},
      {stage2_8[110]}
   );
   gpc1_1 gpc7449 (
      {stage1_8[177]},
      {stage2_8[111]}
   );
   gpc1_1 gpc7450 (
      {stage1_8[178]},
      {stage2_8[112]}
   );
   gpc1_1 gpc7451 (
      {stage1_8[179]},
      {stage2_8[113]}
   );
   gpc1_1 gpc7452 (
      {stage1_8[180]},
      {stage2_8[114]}
   );
   gpc1_1 gpc7453 (
      {stage1_8[181]},
      {stage2_8[115]}
   );
   gpc1_1 gpc7454 (
      {stage1_8[182]},
      {stage2_8[116]}
   );
   gpc1_1 gpc7455 (
      {stage1_8[183]},
      {stage2_8[117]}
   );
   gpc1_1 gpc7456 (
      {stage1_8[184]},
      {stage2_8[118]}
   );
   gpc1_1 gpc7457 (
      {stage1_8[185]},
      {stage2_8[119]}
   );
   gpc1_1 gpc7458 (
      {stage1_8[186]},
      {stage2_8[120]}
   );
   gpc1_1 gpc7459 (
      {stage1_8[187]},
      {stage2_8[121]}
   );
   gpc1_1 gpc7460 (
      {stage1_8[188]},
      {stage2_8[122]}
   );
   gpc1_1 gpc7461 (
      {stage1_8[189]},
      {stage2_8[123]}
   );
   gpc1_1 gpc7462 (
      {stage1_8[190]},
      {stage2_8[124]}
   );
   gpc1_1 gpc7463 (
      {stage1_8[191]},
      {stage2_8[125]}
   );
   gpc1_1 gpc7464 (
      {stage1_8[192]},
      {stage2_8[126]}
   );
   gpc1_1 gpc7465 (
      {stage1_8[193]},
      {stage2_8[127]}
   );
   gpc1_1 gpc7466 (
      {stage1_8[194]},
      {stage2_8[128]}
   );
   gpc1_1 gpc7467 (
      {stage1_8[195]},
      {stage2_8[129]}
   );
   gpc1_1 gpc7468 (
      {stage1_8[196]},
      {stage2_8[130]}
   );
   gpc1_1 gpc7469 (
      {stage1_8[197]},
      {stage2_8[131]}
   );
   gpc1_1 gpc7470 (
      {stage1_8[198]},
      {stage2_8[132]}
   );
   gpc1_1 gpc7471 (
      {stage1_8[199]},
      {stage2_8[133]}
   );
   gpc1_1 gpc7472 (
      {stage1_8[200]},
      {stage2_8[134]}
   );
   gpc1_1 gpc7473 (
      {stage1_8[201]},
      {stage2_8[135]}
   );
   gpc1_1 gpc7474 (
      {stage1_8[202]},
      {stage2_8[136]}
   );
   gpc1_1 gpc7475 (
      {stage1_8[203]},
      {stage2_8[137]}
   );
   gpc1_1 gpc7476 (
      {stage1_8[204]},
      {stage2_8[138]}
   );
   gpc1_1 gpc7477 (
      {stage1_8[205]},
      {stage2_8[139]}
   );
   gpc1_1 gpc7478 (
      {stage1_8[206]},
      {stage2_8[140]}
   );
   gpc1_1 gpc7479 (
      {stage1_8[207]},
      {stage2_8[141]}
   );
   gpc1_1 gpc7480 (
      {stage1_8[208]},
      {stage2_8[142]}
   );
   gpc1_1 gpc7481 (
      {stage1_8[209]},
      {stage2_8[143]}
   );
   gpc1_1 gpc7482 (
      {stage1_8[210]},
      {stage2_8[144]}
   );
   gpc1_1 gpc7483 (
      {stage1_8[211]},
      {stage2_8[145]}
   );
   gpc1_1 gpc7484 (
      {stage1_8[212]},
      {stage2_8[146]}
   );
   gpc1_1 gpc7485 (
      {stage1_8[213]},
      {stage2_8[147]}
   );
   gpc1_1 gpc7486 (
      {stage1_8[214]},
      {stage2_8[148]}
   );
   gpc1_1 gpc7487 (
      {stage1_8[215]},
      {stage2_8[149]}
   );
   gpc1_1 gpc7488 (
      {stage1_8[216]},
      {stage2_8[150]}
   );
   gpc1_1 gpc7489 (
      {stage1_8[217]},
      {stage2_8[151]}
   );
   gpc1_1 gpc7490 (
      {stage1_8[218]},
      {stage2_8[152]}
   );
   gpc1_1 gpc7491 (
      {stage1_8[219]},
      {stage2_8[153]}
   );
   gpc1_1 gpc7492 (
      {stage1_8[220]},
      {stage2_8[154]}
   );
   gpc1_1 gpc7493 (
      {stage1_8[221]},
      {stage2_8[155]}
   );
   gpc1_1 gpc7494 (
      {stage1_8[222]},
      {stage2_8[156]}
   );
   gpc1_1 gpc7495 (
      {stage1_8[223]},
      {stage2_8[157]}
   );
   gpc1_1 gpc7496 (
      {stage1_8[224]},
      {stage2_8[158]}
   );
   gpc1_1 gpc7497 (
      {stage1_8[225]},
      {stage2_8[159]}
   );
   gpc1_1 gpc7498 (
      {stage1_8[226]},
      {stage2_8[160]}
   );
   gpc1_1 gpc7499 (
      {stage1_8[227]},
      {stage2_8[161]}
   );
   gpc1_1 gpc7500 (
      {stage1_8[228]},
      {stage2_8[162]}
   );
   gpc1_1 gpc7501 (
      {stage1_8[229]},
      {stage2_8[163]}
   );
   gpc1_1 gpc7502 (
      {stage1_8[230]},
      {stage2_8[164]}
   );
   gpc1_1 gpc7503 (
      {stage1_8[231]},
      {stage2_8[165]}
   );
   gpc1_1 gpc7504 (
      {stage1_8[232]},
      {stage2_8[166]}
   );
   gpc1_1 gpc7505 (
      {stage1_8[233]},
      {stage2_8[167]}
   );
   gpc1_1 gpc7506 (
      {stage1_8[234]},
      {stage2_8[168]}
   );
   gpc1_1 gpc7507 (
      {stage1_8[235]},
      {stage2_8[169]}
   );
   gpc1_1 gpc7508 (
      {stage1_8[236]},
      {stage2_8[170]}
   );
   gpc1_1 gpc7509 (
      {stage1_8[237]},
      {stage2_8[171]}
   );
   gpc1_1 gpc7510 (
      {stage1_8[238]},
      {stage2_8[172]}
   );
   gpc1_1 gpc7511 (
      {stage1_9[360]},
      {stage2_9[102]}
   );
   gpc1_1 gpc7512 (
      {stage1_9[361]},
      {stage2_9[103]}
   );
   gpc1_1 gpc7513 (
      {stage1_9[362]},
      {stage2_9[104]}
   );
   gpc1_1 gpc7514 (
      {stage1_10[101]},
      {stage2_10[82]}
   );
   gpc1_1 gpc7515 (
      {stage1_10[102]},
      {stage2_10[83]}
   );
   gpc1_1 gpc7516 (
      {stage1_10[103]},
      {stage2_10[84]}
   );
   gpc1_1 gpc7517 (
      {stage1_10[104]},
      {stage2_10[85]}
   );
   gpc1_1 gpc7518 (
      {stage1_10[105]},
      {stage2_10[86]}
   );
   gpc1_1 gpc7519 (
      {stage1_10[106]},
      {stage2_10[87]}
   );
   gpc1_1 gpc7520 (
      {stage1_10[107]},
      {stage2_10[88]}
   );
   gpc1_1 gpc7521 (
      {stage1_10[108]},
      {stage2_10[89]}
   );
   gpc1_1 gpc7522 (
      {stage1_10[109]},
      {stage2_10[90]}
   );
   gpc1_1 gpc7523 (
      {stage1_10[110]},
      {stage2_10[91]}
   );
   gpc1_1 gpc7524 (
      {stage1_10[111]},
      {stage2_10[92]}
   );
   gpc1_1 gpc7525 (
      {stage1_10[112]},
      {stage2_10[93]}
   );
   gpc1_1 gpc7526 (
      {stage1_10[113]},
      {stage2_10[94]}
   );
   gpc1_1 gpc7527 (
      {stage1_10[114]},
      {stage2_10[95]}
   );
   gpc1_1 gpc7528 (
      {stage1_10[115]},
      {stage2_10[96]}
   );
   gpc1_1 gpc7529 (
      {stage1_10[116]},
      {stage2_10[97]}
   );
   gpc1_1 gpc7530 (
      {stage1_10[117]},
      {stage2_10[98]}
   );
   gpc1_1 gpc7531 (
      {stage1_10[118]},
      {stage2_10[99]}
   );
   gpc1_1 gpc7532 (
      {stage1_10[119]},
      {stage2_10[100]}
   );
   gpc1_1 gpc7533 (
      {stage1_10[120]},
      {stage2_10[101]}
   );
   gpc1_1 gpc7534 (
      {stage1_10[121]},
      {stage2_10[102]}
   );
   gpc1_1 gpc7535 (
      {stage1_10[122]},
      {stage2_10[103]}
   );
   gpc1_1 gpc7536 (
      {stage1_10[123]},
      {stage2_10[104]}
   );
   gpc1_1 gpc7537 (
      {stage1_10[124]},
      {stage2_10[105]}
   );
   gpc1_1 gpc7538 (
      {stage1_10[125]},
      {stage2_10[106]}
   );
   gpc1_1 gpc7539 (
      {stage1_10[126]},
      {stage2_10[107]}
   );
   gpc1_1 gpc7540 (
      {stage1_10[127]},
      {stage2_10[108]}
   );
   gpc1_1 gpc7541 (
      {stage1_10[128]},
      {stage2_10[109]}
   );
   gpc1_1 gpc7542 (
      {stage1_10[129]},
      {stage2_10[110]}
   );
   gpc1_1 gpc7543 (
      {stage1_10[130]},
      {stage2_10[111]}
   );
   gpc1_1 gpc7544 (
      {stage1_10[131]},
      {stage2_10[112]}
   );
   gpc1_1 gpc7545 (
      {stage1_10[132]},
      {stage2_10[113]}
   );
   gpc1_1 gpc7546 (
      {stage1_10[133]},
      {stage2_10[114]}
   );
   gpc1_1 gpc7547 (
      {stage1_10[134]},
      {stage2_10[115]}
   );
   gpc1_1 gpc7548 (
      {stage1_10[135]},
      {stage2_10[116]}
   );
   gpc1_1 gpc7549 (
      {stage1_10[136]},
      {stage2_10[117]}
   );
   gpc1_1 gpc7550 (
      {stage1_10[137]},
      {stage2_10[118]}
   );
   gpc1_1 gpc7551 (
      {stage1_10[138]},
      {stage2_10[119]}
   );
   gpc1_1 gpc7552 (
      {stage1_10[139]},
      {stage2_10[120]}
   );
   gpc1_1 gpc7553 (
      {stage1_10[140]},
      {stage2_10[121]}
   );
   gpc1_1 gpc7554 (
      {stage1_10[141]},
      {stage2_10[122]}
   );
   gpc1_1 gpc7555 (
      {stage1_10[142]},
      {stage2_10[123]}
   );
   gpc1_1 gpc7556 (
      {stage1_10[143]},
      {stage2_10[124]}
   );
   gpc1_1 gpc7557 (
      {stage1_10[144]},
      {stage2_10[125]}
   );
   gpc1_1 gpc7558 (
      {stage1_10[145]},
      {stage2_10[126]}
   );
   gpc1_1 gpc7559 (
      {stage1_10[146]},
      {stage2_10[127]}
   );
   gpc1_1 gpc7560 (
      {stage1_10[147]},
      {stage2_10[128]}
   );
   gpc1_1 gpc7561 (
      {stage1_10[148]},
      {stage2_10[129]}
   );
   gpc1_1 gpc7562 (
      {stage1_10[149]},
      {stage2_10[130]}
   );
   gpc1_1 gpc7563 (
      {stage1_10[150]},
      {stage2_10[131]}
   );
   gpc1_1 gpc7564 (
      {stage1_10[151]},
      {stage2_10[132]}
   );
   gpc1_1 gpc7565 (
      {stage1_10[152]},
      {stage2_10[133]}
   );
   gpc1_1 gpc7566 (
      {stage1_11[307]},
      {stage2_11[125]}
   );
   gpc1_1 gpc7567 (
      {stage1_11[308]},
      {stage2_11[126]}
   );
   gpc1_1 gpc7568 (
      {stage1_11[309]},
      {stage2_11[127]}
   );
   gpc1_1 gpc7569 (
      {stage1_11[310]},
      {stage2_11[128]}
   );
   gpc1_1 gpc7570 (
      {stage1_11[311]},
      {stage2_11[129]}
   );
   gpc1_1 gpc7571 (
      {stage1_11[312]},
      {stage2_11[130]}
   );
   gpc1_1 gpc7572 (
      {stage1_11[313]},
      {stage2_11[131]}
   );
   gpc1_1 gpc7573 (
      {stage1_11[314]},
      {stage2_11[132]}
   );
   gpc1_1 gpc7574 (
      {stage1_11[315]},
      {stage2_11[133]}
   );
   gpc1_1 gpc7575 (
      {stage1_11[316]},
      {stage2_11[134]}
   );
   gpc1_1 gpc7576 (
      {stage1_11[317]},
      {stage2_11[135]}
   );
   gpc1_1 gpc7577 (
      {stage1_12[177]},
      {stage2_12[86]}
   );
   gpc1_1 gpc7578 (
      {stage1_12[178]},
      {stage2_12[87]}
   );
   gpc1_1 gpc7579 (
      {stage1_12[179]},
      {stage2_12[88]}
   );
   gpc1_1 gpc7580 (
      {stage1_12[180]},
      {stage2_12[89]}
   );
   gpc1_1 gpc7581 (
      {stage1_12[181]},
      {stage2_12[90]}
   );
   gpc1_1 gpc7582 (
      {stage1_12[182]},
      {stage2_12[91]}
   );
   gpc1_1 gpc7583 (
      {stage1_12[183]},
      {stage2_12[92]}
   );
   gpc1_1 gpc7584 (
      {stage1_12[184]},
      {stage2_12[93]}
   );
   gpc1_1 gpc7585 (
      {stage1_12[185]},
      {stage2_12[94]}
   );
   gpc1_1 gpc7586 (
      {stage1_12[186]},
      {stage2_12[95]}
   );
   gpc1_1 gpc7587 (
      {stage1_12[187]},
      {stage2_12[96]}
   );
   gpc1_1 gpc7588 (
      {stage1_12[188]},
      {stage2_12[97]}
   );
   gpc1_1 gpc7589 (
      {stage1_12[189]},
      {stage2_12[98]}
   );
   gpc1_1 gpc7590 (
      {stage1_12[190]},
      {stage2_12[99]}
   );
   gpc1_1 gpc7591 (
      {stage1_12[191]},
      {stage2_12[100]}
   );
   gpc1_1 gpc7592 (
      {stage1_12[192]},
      {stage2_12[101]}
   );
   gpc1_1 gpc7593 (
      {stage1_12[193]},
      {stage2_12[102]}
   );
   gpc1_1 gpc7594 (
      {stage1_12[194]},
      {stage2_12[103]}
   );
   gpc1_1 gpc7595 (
      {stage1_12[195]},
      {stage2_12[104]}
   );
   gpc1_1 gpc7596 (
      {stage1_12[196]},
      {stage2_12[105]}
   );
   gpc1_1 gpc7597 (
      {stage1_12[197]},
      {stage2_12[106]}
   );
   gpc1_1 gpc7598 (
      {stage1_12[198]},
      {stage2_12[107]}
   );
   gpc1_1 gpc7599 (
      {stage1_12[199]},
      {stage2_12[108]}
   );
   gpc1_1 gpc7600 (
      {stage1_12[200]},
      {stage2_12[109]}
   );
   gpc1_1 gpc7601 (
      {stage1_12[201]},
      {stage2_12[110]}
   );
   gpc1_1 gpc7602 (
      {stage1_12[202]},
      {stage2_12[111]}
   );
   gpc1_1 gpc7603 (
      {stage1_12[203]},
      {stage2_12[112]}
   );
   gpc1_1 gpc7604 (
      {stage1_12[204]},
      {stage2_12[113]}
   );
   gpc1_1 gpc7605 (
      {stage1_12[205]},
      {stage2_12[114]}
   );
   gpc1_1 gpc7606 (
      {stage1_12[206]},
      {stage2_12[115]}
   );
   gpc1_1 gpc7607 (
      {stage1_12[207]},
      {stage2_12[116]}
   );
   gpc1_1 gpc7608 (
      {stage1_12[208]},
      {stage2_12[117]}
   );
   gpc1_1 gpc7609 (
      {stage1_12[209]},
      {stage2_12[118]}
   );
   gpc1_1 gpc7610 (
      {stage1_12[210]},
      {stage2_12[119]}
   );
   gpc1_1 gpc7611 (
      {stage1_12[211]},
      {stage2_12[120]}
   );
   gpc1_1 gpc7612 (
      {stage1_12[212]},
      {stage2_12[121]}
   );
   gpc1_1 gpc7613 (
      {stage1_12[213]},
      {stage2_12[122]}
   );
   gpc1_1 gpc7614 (
      {stage1_12[214]},
      {stage2_12[123]}
   );
   gpc1_1 gpc7615 (
      {stage1_12[215]},
      {stage2_12[124]}
   );
   gpc1_1 gpc7616 (
      {stage1_12[216]},
      {stage2_12[125]}
   );
   gpc1_1 gpc7617 (
      {stage1_12[217]},
      {stage2_12[126]}
   );
   gpc1_1 gpc7618 (
      {stage1_12[218]},
      {stage2_12[127]}
   );
   gpc1_1 gpc7619 (
      {stage1_13[183]},
      {stage2_13[70]}
   );
   gpc1_1 gpc7620 (
      {stage1_13[184]},
      {stage2_13[71]}
   );
   gpc1_1 gpc7621 (
      {stage1_14[246]},
      {stage2_14[105]}
   );
   gpc1_1 gpc7622 (
      {stage1_14[247]},
      {stage2_14[106]}
   );
   gpc1_1 gpc7623 (
      {stage1_14[248]},
      {stage2_14[107]}
   );
   gpc1_1 gpc7624 (
      {stage1_14[249]},
      {stage2_14[108]}
   );
   gpc1_1 gpc7625 (
      {stage1_14[250]},
      {stage2_14[109]}
   );
   gpc1_1 gpc7626 (
      {stage1_14[251]},
      {stage2_14[110]}
   );
   gpc1_1 gpc7627 (
      {stage1_14[252]},
      {stage2_14[111]}
   );
   gpc1_1 gpc7628 (
      {stage1_14[253]},
      {stage2_14[112]}
   );
   gpc1_1 gpc7629 (
      {stage1_14[254]},
      {stage2_14[113]}
   );
   gpc1_1 gpc7630 (
      {stage1_14[255]},
      {stage2_14[114]}
   );
   gpc1_1 gpc7631 (
      {stage1_15[255]},
      {stage2_15[112]}
   );
   gpc1_1 gpc7632 (
      {stage1_15[256]},
      {stage2_15[113]}
   );
   gpc1_1 gpc7633 (
      {stage1_15[257]},
      {stage2_15[114]}
   );
   gpc1_1 gpc7634 (
      {stage1_16[182]},
      {stage2_16[68]}
   );
   gpc1_1 gpc7635 (
      {stage1_16[183]},
      {stage2_16[69]}
   );
   gpc1_1 gpc7636 (
      {stage1_16[184]},
      {stage2_16[70]}
   );
   gpc1_1 gpc7637 (
      {stage1_16[185]},
      {stage2_16[71]}
   );
   gpc1_1 gpc7638 (
      {stage1_16[186]},
      {stage2_16[72]}
   );
   gpc1_1 gpc7639 (
      {stage1_16[187]},
      {stage2_16[73]}
   );
   gpc1_1 gpc7640 (
      {stage1_16[188]},
      {stage2_16[74]}
   );
   gpc1_1 gpc7641 (
      {stage1_16[189]},
      {stage2_16[75]}
   );
   gpc1_1 gpc7642 (
      {stage1_16[190]},
      {stage2_16[76]}
   );
   gpc1_1 gpc7643 (
      {stage1_16[191]},
      {stage2_16[77]}
   );
   gpc1_1 gpc7644 (
      {stage1_16[192]},
      {stage2_16[78]}
   );
   gpc1_1 gpc7645 (
      {stage1_16[193]},
      {stage2_16[79]}
   );
   gpc1_1 gpc7646 (
      {stage1_16[194]},
      {stage2_16[80]}
   );
   gpc1_1 gpc7647 (
      {stage1_16[195]},
      {stage2_16[81]}
   );
   gpc1_1 gpc7648 (
      {stage1_16[196]},
      {stage2_16[82]}
   );
   gpc1_1 gpc7649 (
      {stage1_16[197]},
      {stage2_16[83]}
   );
   gpc1_1 gpc7650 (
      {stage1_16[198]},
      {stage2_16[84]}
   );
   gpc1_1 gpc7651 (
      {stage1_16[199]},
      {stage2_16[85]}
   );
   gpc1_1 gpc7652 (
      {stage1_16[200]},
      {stage2_16[86]}
   );
   gpc1_1 gpc7653 (
      {stage1_16[201]},
      {stage2_16[87]}
   );
   gpc1_1 gpc7654 (
      {stage1_16[202]},
      {stage2_16[88]}
   );
   gpc1_1 gpc7655 (
      {stage1_16[203]},
      {stage2_16[89]}
   );
   gpc1_1 gpc7656 (
      {stage1_16[204]},
      {stage2_16[90]}
   );
   gpc1_1 gpc7657 (
      {stage1_16[205]},
      {stage2_16[91]}
   );
   gpc1_1 gpc7658 (
      {stage1_16[206]},
      {stage2_16[92]}
   );
   gpc1_1 gpc7659 (
      {stage1_16[207]},
      {stage2_16[93]}
   );
   gpc1_1 gpc7660 (
      {stage1_16[208]},
      {stage2_16[94]}
   );
   gpc1_1 gpc7661 (
      {stage1_16[209]},
      {stage2_16[95]}
   );
   gpc1_1 gpc7662 (
      {stage1_16[210]},
      {stage2_16[96]}
   );
   gpc1_1 gpc7663 (
      {stage1_16[211]},
      {stage2_16[97]}
   );
   gpc1_1 gpc7664 (
      {stage1_16[212]},
      {stage2_16[98]}
   );
   gpc1_1 gpc7665 (
      {stage1_16[213]},
      {stage2_16[99]}
   );
   gpc1_1 gpc7666 (
      {stage1_16[214]},
      {stage2_16[100]}
   );
   gpc1_1 gpc7667 (
      {stage1_16[215]},
      {stage2_16[101]}
   );
   gpc1_1 gpc7668 (
      {stage1_16[216]},
      {stage2_16[102]}
   );
   gpc1_1 gpc7669 (
      {stage1_16[217]},
      {stage2_16[103]}
   );
   gpc1_1 gpc7670 (
      {stage1_16[218]},
      {stage2_16[104]}
   );
   gpc1_1 gpc7671 (
      {stage1_16[219]},
      {stage2_16[105]}
   );
   gpc1_1 gpc7672 (
      {stage1_16[220]},
      {stage2_16[106]}
   );
   gpc1_1 gpc7673 (
      {stage1_16[221]},
      {stage2_16[107]}
   );
   gpc1_1 gpc7674 (
      {stage1_16[222]},
      {stage2_16[108]}
   );
   gpc1_1 gpc7675 (
      {stage1_16[223]},
      {stage2_16[109]}
   );
   gpc1_1 gpc7676 (
      {stage1_18[204]},
      {stage2_18[124]}
   );
   gpc1_1 gpc7677 (
      {stage1_18[205]},
      {stage2_18[125]}
   );
   gpc1_1 gpc7678 (
      {stage1_18[206]},
      {stage2_18[126]}
   );
   gpc1_1 gpc7679 (
      {stage1_18[207]},
      {stage2_18[127]}
   );
   gpc1_1 gpc7680 (
      {stage1_18[208]},
      {stage2_18[128]}
   );
   gpc1_1 gpc7681 (
      {stage1_18[209]},
      {stage2_18[129]}
   );
   gpc1_1 gpc7682 (
      {stage1_18[210]},
      {stage2_18[130]}
   );
   gpc1_1 gpc7683 (
      {stage1_18[211]},
      {stage2_18[131]}
   );
   gpc1_1 gpc7684 (
      {stage1_18[212]},
      {stage2_18[132]}
   );
   gpc1_1 gpc7685 (
      {stage1_18[213]},
      {stage2_18[133]}
   );
   gpc1_1 gpc7686 (
      {stage1_18[214]},
      {stage2_18[134]}
   );
   gpc1_1 gpc7687 (
      {stage1_18[215]},
      {stage2_18[135]}
   );
   gpc1_1 gpc7688 (
      {stage1_18[216]},
      {stage2_18[136]}
   );
   gpc1_1 gpc7689 (
      {stage1_18[217]},
      {stage2_18[137]}
   );
   gpc1_1 gpc7690 (
      {stage1_18[218]},
      {stage2_18[138]}
   );
   gpc1_1 gpc7691 (
      {stage1_18[219]},
      {stage2_18[139]}
   );
   gpc1_1 gpc7692 (
      {stage1_18[220]},
      {stage2_18[140]}
   );
   gpc1_1 gpc7693 (
      {stage1_18[221]},
      {stage2_18[141]}
   );
   gpc1_1 gpc7694 (
      {stage1_18[222]},
      {stage2_18[142]}
   );
   gpc1_1 gpc7695 (
      {stage1_18[223]},
      {stage2_18[143]}
   );
   gpc1_1 gpc7696 (
      {stage1_18[224]},
      {stage2_18[144]}
   );
   gpc1_1 gpc7697 (
      {stage1_18[225]},
      {stage2_18[145]}
   );
   gpc1_1 gpc7698 (
      {stage1_18[226]},
      {stage2_18[146]}
   );
   gpc1_1 gpc7699 (
      {stage1_18[227]},
      {stage2_18[147]}
   );
   gpc1_1 gpc7700 (
      {stage1_18[228]},
      {stage2_18[148]}
   );
   gpc1_1 gpc7701 (
      {stage1_18[229]},
      {stage2_18[149]}
   );
   gpc1_1 gpc7702 (
      {stage1_18[230]},
      {stage2_18[150]}
   );
   gpc1_1 gpc7703 (
      {stage1_18[231]},
      {stage2_18[151]}
   );
   gpc1_1 gpc7704 (
      {stage1_18[232]},
      {stage2_18[152]}
   );
   gpc1_1 gpc7705 (
      {stage1_18[233]},
      {stage2_18[153]}
   );
   gpc1_1 gpc7706 (
      {stage1_18[234]},
      {stage2_18[154]}
   );
   gpc1_1 gpc7707 (
      {stage1_18[235]},
      {stage2_18[155]}
   );
   gpc1_1 gpc7708 (
      {stage1_18[236]},
      {stage2_18[156]}
   );
   gpc1_1 gpc7709 (
      {stage1_18[237]},
      {stage2_18[157]}
   );
   gpc1_1 gpc7710 (
      {stage1_18[238]},
      {stage2_18[158]}
   );
   gpc1_1 gpc7711 (
      {stage1_18[239]},
      {stage2_18[159]}
   );
   gpc1_1 gpc7712 (
      {stage1_18[240]},
      {stage2_18[160]}
   );
   gpc1_1 gpc7713 (
      {stage1_18[241]},
      {stage2_18[161]}
   );
   gpc1_1 gpc7714 (
      {stage1_19[201]},
      {stage2_19[76]}
   );
   gpc1_1 gpc7715 (
      {stage1_19[202]},
      {stage2_19[77]}
   );
   gpc1_1 gpc7716 (
      {stage1_19[203]},
      {stage2_19[78]}
   );
   gpc1_1 gpc7717 (
      {stage1_19[204]},
      {stage2_19[79]}
   );
   gpc1_1 gpc7718 (
      {stage1_19[205]},
      {stage2_19[80]}
   );
   gpc1_1 gpc7719 (
      {stage1_19[206]},
      {stage2_19[81]}
   );
   gpc1_1 gpc7720 (
      {stage1_19[207]},
      {stage2_19[82]}
   );
   gpc1_1 gpc7721 (
      {stage1_19[208]},
      {stage2_19[83]}
   );
   gpc1_1 gpc7722 (
      {stage1_19[209]},
      {stage2_19[84]}
   );
   gpc1_1 gpc7723 (
      {stage1_19[210]},
      {stage2_19[85]}
   );
   gpc1_1 gpc7724 (
      {stage1_19[211]},
      {stage2_19[86]}
   );
   gpc1_1 gpc7725 (
      {stage1_19[212]},
      {stage2_19[87]}
   );
   gpc1_1 gpc7726 (
      {stage1_19[213]},
      {stage2_19[88]}
   );
   gpc1_1 gpc7727 (
      {stage1_19[214]},
      {stage2_19[89]}
   );
   gpc1_1 gpc7728 (
      {stage1_19[215]},
      {stage2_19[90]}
   );
   gpc1_1 gpc7729 (
      {stage1_19[216]},
      {stage2_19[91]}
   );
   gpc1_1 gpc7730 (
      {stage1_19[217]},
      {stage2_19[92]}
   );
   gpc1_1 gpc7731 (
      {stage1_19[218]},
      {stage2_19[93]}
   );
   gpc1_1 gpc7732 (
      {stage1_20[227]},
      {stage2_20[71]}
   );
   gpc1_1 gpc7733 (
      {stage1_20[228]},
      {stage2_20[72]}
   );
   gpc1_1 gpc7734 (
      {stage1_20[229]},
      {stage2_20[73]}
   );
   gpc1_1 gpc7735 (
      {stage1_20[230]},
      {stage2_20[74]}
   );
   gpc1_1 gpc7736 (
      {stage1_20[231]},
      {stage2_20[75]}
   );
   gpc1_1 gpc7737 (
      {stage1_20[232]},
      {stage2_20[76]}
   );
   gpc1_1 gpc7738 (
      {stage1_20[233]},
      {stage2_20[77]}
   );
   gpc1_1 gpc7739 (
      {stage1_20[234]},
      {stage2_20[78]}
   );
   gpc1_1 gpc7740 (
      {stage1_20[235]},
      {stage2_20[79]}
   );
   gpc1_1 gpc7741 (
      {stage1_20[236]},
      {stage2_20[80]}
   );
   gpc1_1 gpc7742 (
      {stage1_20[237]},
      {stage2_20[81]}
   );
   gpc1_1 gpc7743 (
      {stage1_20[238]},
      {stage2_20[82]}
   );
   gpc1_1 gpc7744 (
      {stage1_20[239]},
      {stage2_20[83]}
   );
   gpc1_1 gpc7745 (
      {stage1_20[240]},
      {stage2_20[84]}
   );
   gpc1_1 gpc7746 (
      {stage1_20[241]},
      {stage2_20[85]}
   );
   gpc1_1 gpc7747 (
      {stage1_20[242]},
      {stage2_20[86]}
   );
   gpc1_1 gpc7748 (
      {stage1_20[243]},
      {stage2_20[87]}
   );
   gpc1_1 gpc7749 (
      {stage1_21[186]},
      {stage2_21[93]}
   );
   gpc1_1 gpc7750 (
      {stage1_21[187]},
      {stage2_21[94]}
   );
   gpc1_1 gpc7751 (
      {stage1_21[188]},
      {stage2_21[95]}
   );
   gpc1_1 gpc7752 (
      {stage1_21[189]},
      {stage2_21[96]}
   );
   gpc1_1 gpc7753 (
      {stage1_21[190]},
      {stage2_21[97]}
   );
   gpc1_1 gpc7754 (
      {stage1_21[191]},
      {stage2_21[98]}
   );
   gpc1_1 gpc7755 (
      {stage1_21[192]},
      {stage2_21[99]}
   );
   gpc1_1 gpc7756 (
      {stage1_21[193]},
      {stage2_21[100]}
   );
   gpc1_1 gpc7757 (
      {stage1_21[194]},
      {stage2_21[101]}
   );
   gpc1_1 gpc7758 (
      {stage1_21[195]},
      {stage2_21[102]}
   );
   gpc1_1 gpc7759 (
      {stage1_21[196]},
      {stage2_21[103]}
   );
   gpc1_1 gpc7760 (
      {stage1_21[197]},
      {stage2_21[104]}
   );
   gpc1_1 gpc7761 (
      {stage1_21[198]},
      {stage2_21[105]}
   );
   gpc1_1 gpc7762 (
      {stage1_21[199]},
      {stage2_21[106]}
   );
   gpc1_1 gpc7763 (
      {stage1_21[200]},
      {stage2_21[107]}
   );
   gpc1_1 gpc7764 (
      {stage1_21[201]},
      {stage2_21[108]}
   );
   gpc1_1 gpc7765 (
      {stage1_21[202]},
      {stage2_21[109]}
   );
   gpc1_1 gpc7766 (
      {stage1_21[203]},
      {stage2_21[110]}
   );
   gpc1_1 gpc7767 (
      {stage1_21[204]},
      {stage2_21[111]}
   );
   gpc1_1 gpc7768 (
      {stage1_22[194]},
      {stage2_22[103]}
   );
   gpc1_1 gpc7769 (
      {stage1_22[195]},
      {stage2_22[104]}
   );
   gpc1_1 gpc7770 (
      {stage1_22[196]},
      {stage2_22[105]}
   );
   gpc1_1 gpc7771 (
      {stage1_22[197]},
      {stage2_22[106]}
   );
   gpc1_1 gpc7772 (
      {stage1_22[198]},
      {stage2_22[107]}
   );
   gpc1_1 gpc7773 (
      {stage1_22[199]},
      {stage2_22[108]}
   );
   gpc1_1 gpc7774 (
      {stage1_22[200]},
      {stage2_22[109]}
   );
   gpc1_1 gpc7775 (
      {stage1_23[290]},
      {stage2_23[89]}
   );
   gpc1_1 gpc7776 (
      {stage1_23[291]},
      {stage2_23[90]}
   );
   gpc1_1 gpc7777 (
      {stage1_23[292]},
      {stage2_23[91]}
   );
   gpc1_1 gpc7778 (
      {stage1_23[293]},
      {stage2_23[92]}
   );
   gpc1_1 gpc7779 (
      {stage1_23[294]},
      {stage2_23[93]}
   );
   gpc1_1 gpc7780 (
      {stage1_23[295]},
      {stage2_23[94]}
   );
   gpc1_1 gpc7781 (
      {stage1_23[296]},
      {stage2_23[95]}
   );
   gpc1_1 gpc7782 (
      {stage1_23[297]},
      {stage2_23[96]}
   );
   gpc1_1 gpc7783 (
      {stage1_23[298]},
      {stage2_23[97]}
   );
   gpc1_1 gpc7784 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc7785 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc7786 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc7787 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc7788 (
      {stage1_25[184]},
      {stage2_25[96]}
   );
   gpc1_1 gpc7789 (
      {stage1_25[185]},
      {stage2_25[97]}
   );
   gpc1_1 gpc7790 (
      {stage1_25[186]},
      {stage2_25[98]}
   );
   gpc1_1 gpc7791 (
      {stage1_25[187]},
      {stage2_25[99]}
   );
   gpc1_1 gpc7792 (
      {stage1_25[188]},
      {stage2_25[100]}
   );
   gpc1_1 gpc7793 (
      {stage1_25[189]},
      {stage2_25[101]}
   );
   gpc1_1 gpc7794 (
      {stage1_25[190]},
      {stage2_25[102]}
   );
   gpc1_1 gpc7795 (
      {stage1_25[191]},
      {stage2_25[103]}
   );
   gpc1_1 gpc7796 (
      {stage1_25[192]},
      {stage2_25[104]}
   );
   gpc1_1 gpc7797 (
      {stage1_25[193]},
      {stage2_25[105]}
   );
   gpc1_1 gpc7798 (
      {stage1_25[194]},
      {stage2_25[106]}
   );
   gpc1_1 gpc7799 (
      {stage1_25[195]},
      {stage2_25[107]}
   );
   gpc1_1 gpc7800 (
      {stage1_25[196]},
      {stage2_25[108]}
   );
   gpc1_1 gpc7801 (
      {stage1_25[197]},
      {stage2_25[109]}
   );
   gpc1_1 gpc7802 (
      {stage1_25[198]},
      {stage2_25[110]}
   );
   gpc1_1 gpc7803 (
      {stage1_25[199]},
      {stage2_25[111]}
   );
   gpc1_1 gpc7804 (
      {stage1_25[200]},
      {stage2_25[112]}
   );
   gpc1_1 gpc7805 (
      {stage1_25[201]},
      {stage2_25[113]}
   );
   gpc1_1 gpc7806 (
      {stage1_25[202]},
      {stage2_25[114]}
   );
   gpc1_1 gpc7807 (
      {stage1_25[203]},
      {stage2_25[115]}
   );
   gpc1_1 gpc7808 (
      {stage1_25[204]},
      {stage2_25[116]}
   );
   gpc1_1 gpc7809 (
      {stage1_25[205]},
      {stage2_25[117]}
   );
   gpc1_1 gpc7810 (
      {stage1_25[206]},
      {stage2_25[118]}
   );
   gpc1_1 gpc7811 (
      {stage1_25[207]},
      {stage2_25[119]}
   );
   gpc1_1 gpc7812 (
      {stage1_25[208]},
      {stage2_25[120]}
   );
   gpc1_1 gpc7813 (
      {stage1_25[209]},
      {stage2_25[121]}
   );
   gpc1_1 gpc7814 (
      {stage1_25[210]},
      {stage2_25[122]}
   );
   gpc1_1 gpc7815 (
      {stage1_26[154]},
      {stage2_26[96]}
   );
   gpc1_1 gpc7816 (
      {stage1_26[155]},
      {stage2_26[97]}
   );
   gpc1_1 gpc7817 (
      {stage1_26[156]},
      {stage2_26[98]}
   );
   gpc1_1 gpc7818 (
      {stage1_26[157]},
      {stage2_26[99]}
   );
   gpc1_1 gpc7819 (
      {stage1_26[158]},
      {stage2_26[100]}
   );
   gpc1_1 gpc7820 (
      {stage1_26[159]},
      {stage2_26[101]}
   );
   gpc1_1 gpc7821 (
      {stage1_26[160]},
      {stage2_26[102]}
   );
   gpc1_1 gpc7822 (
      {stage1_26[161]},
      {stage2_26[103]}
   );
   gpc1_1 gpc7823 (
      {stage1_26[162]},
      {stage2_26[104]}
   );
   gpc1_1 gpc7824 (
      {stage1_26[163]},
      {stage2_26[105]}
   );
   gpc1_1 gpc7825 (
      {stage1_26[164]},
      {stage2_26[106]}
   );
   gpc1_1 gpc7826 (
      {stage1_26[165]},
      {stage2_26[107]}
   );
   gpc1_1 gpc7827 (
      {stage1_26[166]},
      {stage2_26[108]}
   );
   gpc1_1 gpc7828 (
      {stage1_26[167]},
      {stage2_26[109]}
   );
   gpc1_1 gpc7829 (
      {stage1_26[168]},
      {stage2_26[110]}
   );
   gpc1_1 gpc7830 (
      {stage1_26[169]},
      {stage2_26[111]}
   );
   gpc1_1 gpc7831 (
      {stage1_26[170]},
      {stage2_26[112]}
   );
   gpc1_1 gpc7832 (
      {stage1_26[171]},
      {stage2_26[113]}
   );
   gpc1_1 gpc7833 (
      {stage1_26[172]},
      {stage2_26[114]}
   );
   gpc1_1 gpc7834 (
      {stage1_26[173]},
      {stage2_26[115]}
   );
   gpc1_1 gpc7835 (
      {stage1_26[174]},
      {stage2_26[116]}
   );
   gpc1_1 gpc7836 (
      {stage1_26[175]},
      {stage2_26[117]}
   );
   gpc1_1 gpc7837 (
      {stage1_26[176]},
      {stage2_26[118]}
   );
   gpc1_1 gpc7838 (
      {stage1_26[177]},
      {stage2_26[119]}
   );
   gpc1_1 gpc7839 (
      {stage1_26[178]},
      {stage2_26[120]}
   );
   gpc1_1 gpc7840 (
      {stage1_26[179]},
      {stage2_26[121]}
   );
   gpc1_1 gpc7841 (
      {stage1_26[180]},
      {stage2_26[122]}
   );
   gpc1_1 gpc7842 (
      {stage1_26[181]},
      {stage2_26[123]}
   );
   gpc1_1 gpc7843 (
      {stage1_26[182]},
      {stage2_26[124]}
   );
   gpc1_1 gpc7844 (
      {stage1_26[183]},
      {stage2_26[125]}
   );
   gpc1_1 gpc7845 (
      {stage1_26[184]},
      {stage2_26[126]}
   );
   gpc1_1 gpc7846 (
      {stage1_26[185]},
      {stage2_26[127]}
   );
   gpc1_1 gpc7847 (
      {stage1_26[186]},
      {stage2_26[128]}
   );
   gpc1_1 gpc7848 (
      {stage1_26[187]},
      {stage2_26[129]}
   );
   gpc1_1 gpc7849 (
      {stage1_26[188]},
      {stage2_26[130]}
   );
   gpc1_1 gpc7850 (
      {stage1_27[211]},
      {stage2_27[85]}
   );
   gpc1_1 gpc7851 (
      {stage1_28[240]},
      {stage2_28[71]}
   );
   gpc1_1 gpc7852 (
      {stage1_28[241]},
      {stage2_28[72]}
   );
   gpc1_1 gpc7853 (
      {stage1_28[242]},
      {stage2_28[73]}
   );
   gpc1_1 gpc7854 (
      {stage1_28[243]},
      {stage2_28[74]}
   );
   gpc1_1 gpc7855 (
      {stage1_28[244]},
      {stage2_28[75]}
   );
   gpc1_1 gpc7856 (
      {stage1_28[245]},
      {stage2_28[76]}
   );
   gpc1_1 gpc7857 (
      {stage1_28[246]},
      {stage2_28[77]}
   );
   gpc1_1 gpc7858 (
      {stage1_28[247]},
      {stage2_28[78]}
   );
   gpc1_1 gpc7859 (
      {stage1_28[248]},
      {stage2_28[79]}
   );
   gpc1_1 gpc7860 (
      {stage1_29[186]},
      {stage2_29[77]}
   );
   gpc1_1 gpc7861 (
      {stage1_29[187]},
      {stage2_29[78]}
   );
   gpc1_1 gpc7862 (
      {stage1_29[188]},
      {stage2_29[79]}
   );
   gpc1_1 gpc7863 (
      {stage1_29[189]},
      {stage2_29[80]}
   );
   gpc1_1 gpc7864 (
      {stage1_29[190]},
      {stage2_29[81]}
   );
   gpc1_1 gpc7865 (
      {stage1_29[191]},
      {stage2_29[82]}
   );
   gpc1_1 gpc7866 (
      {stage1_29[192]},
      {stage2_29[83]}
   );
   gpc1_1 gpc7867 (
      {stage1_29[193]},
      {stage2_29[84]}
   );
   gpc1_1 gpc7868 (
      {stage1_29[194]},
      {stage2_29[85]}
   );
   gpc1_1 gpc7869 (
      {stage1_29[195]},
      {stage2_29[86]}
   );
   gpc1_1 gpc7870 (
      {stage1_29[196]},
      {stage2_29[87]}
   );
   gpc1_1 gpc7871 (
      {stage1_29[197]},
      {stage2_29[88]}
   );
   gpc1_1 gpc7872 (
      {stage1_29[198]},
      {stage2_29[89]}
   );
   gpc1_1 gpc7873 (
      {stage1_29[199]},
      {stage2_29[90]}
   );
   gpc1_1 gpc7874 (
      {stage1_29[200]},
      {stage2_29[91]}
   );
   gpc1_1 gpc7875 (
      {stage1_29[201]},
      {stage2_29[92]}
   );
   gpc1_1 gpc7876 (
      {stage1_29[202]},
      {stage2_29[93]}
   );
   gpc1_1 gpc7877 (
      {stage1_29[203]},
      {stage2_29[94]}
   );
   gpc1_1 gpc7878 (
      {stage1_29[204]},
      {stage2_29[95]}
   );
   gpc1_1 gpc7879 (
      {stage1_29[205]},
      {stage2_29[96]}
   );
   gpc1_1 gpc7880 (
      {stage1_29[206]},
      {stage2_29[97]}
   );
   gpc1_1 gpc7881 (
      {stage1_29[207]},
      {stage2_29[98]}
   );
   gpc1_1 gpc7882 (
      {stage1_29[208]},
      {stage2_29[99]}
   );
   gpc1_1 gpc7883 (
      {stage1_29[209]},
      {stage2_29[100]}
   );
   gpc1_1 gpc7884 (
      {stage1_29[210]},
      {stage2_29[101]}
   );
   gpc1_1 gpc7885 (
      {stage1_29[211]},
      {stage2_29[102]}
   );
   gpc1_1 gpc7886 (
      {stage1_29[212]},
      {stage2_29[103]}
   );
   gpc1_1 gpc7887 (
      {stage1_29[213]},
      {stage2_29[104]}
   );
   gpc1_1 gpc7888 (
      {stage1_29[214]},
      {stage2_29[105]}
   );
   gpc1_1 gpc7889 (
      {stage1_29[215]},
      {stage2_29[106]}
   );
   gpc1_1 gpc7890 (
      {stage1_29[216]},
      {stage2_29[107]}
   );
   gpc1_1 gpc7891 (
      {stage1_29[217]},
      {stage2_29[108]}
   );
   gpc1_1 gpc7892 (
      {stage1_29[218]},
      {stage2_29[109]}
   );
   gpc1_1 gpc7893 (
      {stage1_29[219]},
      {stage2_29[110]}
   );
   gpc1_1 gpc7894 (
      {stage1_29[220]},
      {stage2_29[111]}
   );
   gpc1_1 gpc7895 (
      {stage1_30[232]},
      {stage2_30[99]}
   );
   gpc1_1 gpc7896 (
      {stage1_31[180]},
      {stage2_31[96]}
   );
   gpc1_1 gpc7897 (
      {stage1_31[181]},
      {stage2_31[97]}
   );
   gpc1_1 gpc7898 (
      {stage1_31[182]},
      {stage2_31[98]}
   );
   gpc1_1 gpc7899 (
      {stage1_31[183]},
      {stage2_31[99]}
   );
   gpc1_1 gpc7900 (
      {stage1_31[184]},
      {stage2_31[100]}
   );
   gpc1_1 gpc7901 (
      {stage1_31[185]},
      {stage2_31[101]}
   );
   gpc1_1 gpc7902 (
      {stage1_31[186]},
      {stage2_31[102]}
   );
   gpc1_1 gpc7903 (
      {stage1_31[187]},
      {stage2_31[103]}
   );
   gpc1_1 gpc7904 (
      {stage1_31[188]},
      {stage2_31[104]}
   );
   gpc1_1 gpc7905 (
      {stage1_31[189]},
      {stage2_31[105]}
   );
   gpc1_1 gpc7906 (
      {stage1_31[190]},
      {stage2_31[106]}
   );
   gpc1_1 gpc7907 (
      {stage1_31[191]},
      {stage2_31[107]}
   );
   gpc1_1 gpc7908 (
      {stage1_31[192]},
      {stage2_31[108]}
   );
   gpc1_1 gpc7909 (
      {stage1_31[193]},
      {stage2_31[109]}
   );
   gpc1_1 gpc7910 (
      {stage1_31[194]},
      {stage2_31[110]}
   );
   gpc1_1 gpc7911 (
      {stage1_31[195]},
      {stage2_31[111]}
   );
   gpc1_1 gpc7912 (
      {stage1_31[196]},
      {stage2_31[112]}
   );
   gpc1_1 gpc7913 (
      {stage1_31[197]},
      {stage2_31[113]}
   );
   gpc1_1 gpc7914 (
      {stage1_31[198]},
      {stage2_31[114]}
   );
   gpc1_1 gpc7915 (
      {stage1_31[199]},
      {stage2_31[115]}
   );
   gpc1_1 gpc7916 (
      {stage1_31[200]},
      {stage2_31[116]}
   );
   gpc1_1 gpc7917 (
      {stage1_31[201]},
      {stage2_31[117]}
   );
   gpc1_1 gpc7918 (
      {stage1_31[202]},
      {stage2_31[118]}
   );
   gpc1_1 gpc7919 (
      {stage1_31[203]},
      {stage2_31[119]}
   );
   gpc1_1 gpc7920 (
      {stage1_31[204]},
      {stage2_31[120]}
   );
   gpc1_1 gpc7921 (
      {stage1_31[205]},
      {stage2_31[121]}
   );
   gpc1_1 gpc7922 (
      {stage1_31[206]},
      {stage2_31[122]}
   );
   gpc1_1 gpc7923 (
      {stage1_31[207]},
      {stage2_31[123]}
   );
   gpc1_1 gpc7924 (
      {stage1_31[208]},
      {stage2_31[124]}
   );
   gpc1_1 gpc7925 (
      {stage1_31[209]},
      {stage2_31[125]}
   );
   gpc1_1 gpc7926 (
      {stage1_31[210]},
      {stage2_31[126]}
   );
   gpc1_1 gpc7927 (
      {stage1_31[211]},
      {stage2_31[127]}
   );
   gpc1_1 gpc7928 (
      {stage1_32[404]},
      {stage2_32[107]}
   );
   gpc1_1 gpc7929 (
      {stage1_32[405]},
      {stage2_32[108]}
   );
   gpc1_1 gpc7930 (
      {stage1_32[406]},
      {stage2_32[109]}
   );
   gpc1_1 gpc7931 (
      {stage1_32[407]},
      {stage2_32[110]}
   );
   gpc1_1 gpc7932 (
      {stage1_32[408]},
      {stage2_32[111]}
   );
   gpc1_1 gpc7933 (
      {stage1_32[409]},
      {stage2_32[112]}
   );
   gpc1_1 gpc7934 (
      {stage1_32[410]},
      {stage2_32[113]}
   );
   gpc1_1 gpc7935 (
      {stage1_32[411]},
      {stage2_32[114]}
   );
   gpc1_1 gpc7936 (
      {stage1_32[412]},
      {stage2_32[115]}
   );
   gpc1_1 gpc7937 (
      {stage1_32[413]},
      {stage2_32[116]}
   );
   gpc1_1 gpc7938 (
      {stage1_32[414]},
      {stage2_32[117]}
   );
   gpc1_1 gpc7939 (
      {stage1_34[242]},
      {stage2_34[102]}
   );
   gpc1_1 gpc7940 (
      {stage1_34[243]},
      {stage2_34[103]}
   );
   gpc1_1 gpc7941 (
      {stage1_34[244]},
      {stage2_34[104]}
   );
   gpc1_1 gpc7942 (
      {stage1_34[245]},
      {stage2_34[105]}
   );
   gpc1_1 gpc7943 (
      {stage1_34[246]},
      {stage2_34[106]}
   );
   gpc1_1 gpc7944 (
      {stage1_34[247]},
      {stage2_34[107]}
   );
   gpc1_1 gpc7945 (
      {stage1_34[248]},
      {stage2_34[108]}
   );
   gpc1_1 gpc7946 (
      {stage1_34[249]},
      {stage2_34[109]}
   );
   gpc1_1 gpc7947 (
      {stage1_34[250]},
      {stage2_34[110]}
   );
   gpc1_1 gpc7948 (
      {stage1_34[251]},
      {stage2_34[111]}
   );
   gpc1_1 gpc7949 (
      {stage1_34[252]},
      {stage2_34[112]}
   );
   gpc1_1 gpc7950 (
      {stage1_34[253]},
      {stage2_34[113]}
   );
   gpc1_1 gpc7951 (
      {stage1_34[254]},
      {stage2_34[114]}
   );
   gpc1_1 gpc7952 (
      {stage1_34[255]},
      {stage2_34[115]}
   );
   gpc1_1 gpc7953 (
      {stage1_34[256]},
      {stage2_34[116]}
   );
   gpc1_1 gpc7954 (
      {stage1_34[257]},
      {stage2_34[117]}
   );
   gpc1_1 gpc7955 (
      {stage1_34[258]},
      {stage2_34[118]}
   );
   gpc1_1 gpc7956 (
      {stage1_34[259]},
      {stage2_34[119]}
   );
   gpc1_1 gpc7957 (
      {stage1_34[260]},
      {stage2_34[120]}
   );
   gpc1_1 gpc7958 (
      {stage1_34[261]},
      {stage2_34[121]}
   );
   gpc1_1 gpc7959 (
      {stage1_34[262]},
      {stage2_34[122]}
   );
   gpc1_1 gpc7960 (
      {stage1_34[263]},
      {stage2_34[123]}
   );
   gpc1_1 gpc7961 (
      {stage1_34[264]},
      {stage2_34[124]}
   );
   gpc1_1 gpc7962 (
      {stage1_34[265]},
      {stage2_34[125]}
   );
   gpc1_1 gpc7963 (
      {stage1_34[266]},
      {stage2_34[126]}
   );
   gpc1_1 gpc7964 (
      {stage1_34[267]},
      {stage2_34[127]}
   );
   gpc1_1 gpc7965 (
      {stage1_35[173]},
      {stage2_35[100]}
   );
   gpc1_1 gpc7966 (
      {stage1_35[174]},
      {stage2_35[101]}
   );
   gpc1_1 gpc7967 (
      {stage1_35[175]},
      {stage2_35[102]}
   );
   gpc1_1 gpc7968 (
      {stage1_35[176]},
      {stage2_35[103]}
   );
   gpc1_1 gpc7969 (
      {stage1_35[177]},
      {stage2_35[104]}
   );
   gpc1_1 gpc7970 (
      {stage1_35[178]},
      {stage2_35[105]}
   );
   gpc1_1 gpc7971 (
      {stage1_35[179]},
      {stage2_35[106]}
   );
   gpc1_1 gpc7972 (
      {stage1_35[180]},
      {stage2_35[107]}
   );
   gpc1_1 gpc7973 (
      {stage1_35[181]},
      {stage2_35[108]}
   );
   gpc1_1 gpc7974 (
      {stage1_35[182]},
      {stage2_35[109]}
   );
   gpc1_1 gpc7975 (
      {stage1_35[183]},
      {stage2_35[110]}
   );
   gpc1_1 gpc7976 (
      {stage1_35[184]},
      {stage2_35[111]}
   );
   gpc1_1 gpc7977 (
      {stage1_35[185]},
      {stage2_35[112]}
   );
   gpc1_1 gpc7978 (
      {stage1_35[186]},
      {stage2_35[113]}
   );
   gpc1_1 gpc7979 (
      {stage1_35[187]},
      {stage2_35[114]}
   );
   gpc1_1 gpc7980 (
      {stage1_35[188]},
      {stage2_35[115]}
   );
   gpc1_1 gpc7981 (
      {stage1_35[189]},
      {stage2_35[116]}
   );
   gpc1_1 gpc7982 (
      {stage1_35[190]},
      {stage2_35[117]}
   );
   gpc1_1 gpc7983 (
      {stage1_37[297]},
      {stage2_37[108]}
   );
   gpc1_1 gpc7984 (
      {stage1_37[298]},
      {stage2_37[109]}
   );
   gpc1_1 gpc7985 (
      {stage1_37[299]},
      {stage2_37[110]}
   );
   gpc1_1 gpc7986 (
      {stage1_37[300]},
      {stage2_37[111]}
   );
   gpc1_1 gpc7987 (
      {stage1_37[301]},
      {stage2_37[112]}
   );
   gpc1_1 gpc7988 (
      {stage1_37[302]},
      {stage2_37[113]}
   );
   gpc1_1 gpc7989 (
      {stage1_39[194]},
      {stage2_39[105]}
   );
   gpc1_1 gpc7990 (
      {stage1_39[195]},
      {stage2_39[106]}
   );
   gpc1_1 gpc7991 (
      {stage1_39[196]},
      {stage2_39[107]}
   );
   gpc1_1 gpc7992 (
      {stage1_40[203]},
      {stage2_40[113]}
   );
   gpc1_1 gpc7993 (
      {stage1_40[204]},
      {stage2_40[114]}
   );
   gpc1_1 gpc7994 (
      {stage1_40[205]},
      {stage2_40[115]}
   );
   gpc1_1 gpc7995 (
      {stage1_40[206]},
      {stage2_40[116]}
   );
   gpc1_1 gpc7996 (
      {stage1_40[207]},
      {stage2_40[117]}
   );
   gpc1_1 gpc7997 (
      {stage1_40[208]},
      {stage2_40[118]}
   );
   gpc1_1 gpc7998 (
      {stage1_40[209]},
      {stage2_40[119]}
   );
   gpc1_1 gpc7999 (
      {stage1_40[210]},
      {stage2_40[120]}
   );
   gpc1_1 gpc8000 (
      {stage1_40[211]},
      {stage2_40[121]}
   );
   gpc1_1 gpc8001 (
      {stage1_40[212]},
      {stage2_40[122]}
   );
   gpc1_1 gpc8002 (
      {stage1_40[213]},
      {stage2_40[123]}
   );
   gpc1_1 gpc8003 (
      {stage1_40[214]},
      {stage2_40[124]}
   );
   gpc1_1 gpc8004 (
      {stage1_40[215]},
      {stage2_40[125]}
   );
   gpc1_1 gpc8005 (
      {stage1_40[216]},
      {stage2_40[126]}
   );
   gpc1_1 gpc8006 (
      {stage1_40[217]},
      {stage2_40[127]}
   );
   gpc1_1 gpc8007 (
      {stage1_40[218]},
      {stage2_40[128]}
   );
   gpc1_1 gpc8008 (
      {stage1_40[219]},
      {stage2_40[129]}
   );
   gpc1_1 gpc8009 (
      {stage1_40[220]},
      {stage2_40[130]}
   );
   gpc1_1 gpc8010 (
      {stage1_40[221]},
      {stage2_40[131]}
   );
   gpc1_1 gpc8011 (
      {stage1_40[222]},
      {stage2_40[132]}
   );
   gpc1_1 gpc8012 (
      {stage1_40[223]},
      {stage2_40[133]}
   );
   gpc1_1 gpc8013 (
      {stage1_40[224]},
      {stage2_40[134]}
   );
   gpc1_1 gpc8014 (
      {stage1_40[225]},
      {stage2_40[135]}
   );
   gpc1_1 gpc8015 (
      {stage1_40[226]},
      {stage2_40[136]}
   );
   gpc1_1 gpc8016 (
      {stage1_40[227]},
      {stage2_40[137]}
   );
   gpc1_1 gpc8017 (
      {stage1_40[228]},
      {stage2_40[138]}
   );
   gpc1_1 gpc8018 (
      {stage1_40[229]},
      {stage2_40[139]}
   );
   gpc1_1 gpc8019 (
      {stage1_41[252]},
      {stage2_41[98]}
   );
   gpc1_1 gpc8020 (
      {stage1_41[253]},
      {stage2_41[99]}
   );
   gpc1_1 gpc8021 (
      {stage1_41[254]},
      {stage2_41[100]}
   );
   gpc1_1 gpc8022 (
      {stage1_41[255]},
      {stage2_41[101]}
   );
   gpc1_1 gpc8023 (
      {stage1_41[256]},
      {stage2_41[102]}
   );
   gpc1_1 gpc8024 (
      {stage1_41[257]},
      {stage2_41[103]}
   );
   gpc1_1 gpc8025 (
      {stage1_41[258]},
      {stage2_41[104]}
   );
   gpc1_1 gpc8026 (
      {stage1_41[259]},
      {stage2_41[105]}
   );
   gpc1_1 gpc8027 (
      {stage1_41[260]},
      {stage2_41[106]}
   );
   gpc1_1 gpc8028 (
      {stage1_41[261]},
      {stage2_41[107]}
   );
   gpc1_1 gpc8029 (
      {stage1_41[262]},
      {stage2_41[108]}
   );
   gpc1_1 gpc8030 (
      {stage1_41[263]},
      {stage2_41[109]}
   );
   gpc1_1 gpc8031 (
      {stage1_41[264]},
      {stage2_41[110]}
   );
   gpc1_1 gpc8032 (
      {stage1_41[265]},
      {stage2_41[111]}
   );
   gpc1_1 gpc8033 (
      {stage1_41[266]},
      {stage2_41[112]}
   );
   gpc1_1 gpc8034 (
      {stage1_41[267]},
      {stage2_41[113]}
   );
   gpc1_1 gpc8035 (
      {stage1_41[268]},
      {stage2_41[114]}
   );
   gpc1_1 gpc8036 (
      {stage1_41[269]},
      {stage2_41[115]}
   );
   gpc1_1 gpc8037 (
      {stage1_41[270]},
      {stage2_41[116]}
   );
   gpc1_1 gpc8038 (
      {stage1_41[271]},
      {stage2_41[117]}
   );
   gpc1_1 gpc8039 (
      {stage1_41[272]},
      {stage2_41[118]}
   );
   gpc1_1 gpc8040 (
      {stage1_41[273]},
      {stage2_41[119]}
   );
   gpc1_1 gpc8041 (
      {stage1_41[274]},
      {stage2_41[120]}
   );
   gpc1_1 gpc8042 (
      {stage1_41[275]},
      {stage2_41[121]}
   );
   gpc1_1 gpc8043 (
      {stage1_41[276]},
      {stage2_41[122]}
   );
   gpc1_1 gpc8044 (
      {stage1_42[228]},
      {stage2_42[81]}
   );
   gpc1_1 gpc8045 (
      {stage1_43[218]},
      {stage2_43[85]}
   );
   gpc1_1 gpc8046 (
      {stage1_43[219]},
      {stage2_43[86]}
   );
   gpc1_1 gpc8047 (
      {stage1_43[220]},
      {stage2_43[87]}
   );
   gpc1_1 gpc8048 (
      {stage1_43[221]},
      {stage2_43[88]}
   );
   gpc1_1 gpc8049 (
      {stage1_43[222]},
      {stage2_43[89]}
   );
   gpc1_1 gpc8050 (
      {stage1_43[223]},
      {stage2_43[90]}
   );
   gpc1_1 gpc8051 (
      {stage1_43[224]},
      {stage2_43[91]}
   );
   gpc1_1 gpc8052 (
      {stage1_43[225]},
      {stage2_43[92]}
   );
   gpc1_1 gpc8053 (
      {stage1_43[226]},
      {stage2_43[93]}
   );
   gpc1_1 gpc8054 (
      {stage1_43[227]},
      {stage2_43[94]}
   );
   gpc1_1 gpc8055 (
      {stage1_43[228]},
      {stage2_43[95]}
   );
   gpc1_1 gpc8056 (
      {stage1_43[229]},
      {stage2_43[96]}
   );
   gpc1_1 gpc8057 (
      {stage1_43[230]},
      {stage2_43[97]}
   );
   gpc1_1 gpc8058 (
      {stage1_43[231]},
      {stage2_43[98]}
   );
   gpc1_1 gpc8059 (
      {stage1_43[232]},
      {stage2_43[99]}
   );
   gpc1_1 gpc8060 (
      {stage1_43[233]},
      {stage2_43[100]}
   );
   gpc1_1 gpc8061 (
      {stage1_43[234]},
      {stage2_43[101]}
   );
   gpc1_1 gpc8062 (
      {stage1_43[235]},
      {stage2_43[102]}
   );
   gpc1_1 gpc8063 (
      {stage1_43[236]},
      {stage2_43[103]}
   );
   gpc1_1 gpc8064 (
      {stage1_43[237]},
      {stage2_43[104]}
   );
   gpc1_1 gpc8065 (
      {stage1_43[238]},
      {stage2_43[105]}
   );
   gpc1_1 gpc8066 (
      {stage1_43[239]},
      {stage2_43[106]}
   );
   gpc1_1 gpc8067 (
      {stage1_43[240]},
      {stage2_43[107]}
   );
   gpc1_1 gpc8068 (
      {stage1_43[241]},
      {stage2_43[108]}
   );
   gpc1_1 gpc8069 (
      {stage1_43[242]},
      {stage2_43[109]}
   );
   gpc1_1 gpc8070 (
      {stage1_43[243]},
      {stage2_43[110]}
   );
   gpc1_1 gpc8071 (
      {stage1_44[244]},
      {stage2_44[113]}
   );
   gpc1_1 gpc8072 (
      {stage1_44[245]},
      {stage2_44[114]}
   );
   gpc1_1 gpc8073 (
      {stage1_44[246]},
      {stage2_44[115]}
   );
   gpc1_1 gpc8074 (
      {stage1_44[247]},
      {stage2_44[116]}
   );
   gpc1_1 gpc8075 (
      {stage1_44[248]},
      {stage2_44[117]}
   );
   gpc1_1 gpc8076 (
      {stage1_44[249]},
      {stage2_44[118]}
   );
   gpc1_1 gpc8077 (
      {stage1_44[250]},
      {stage2_44[119]}
   );
   gpc1_1 gpc8078 (
      {stage1_44[251]},
      {stage2_44[120]}
   );
   gpc1_1 gpc8079 (
      {stage1_44[252]},
      {stage2_44[121]}
   );
   gpc1_1 gpc8080 (
      {stage1_44[253]},
      {stage2_44[122]}
   );
   gpc1_1 gpc8081 (
      {stage1_44[254]},
      {stage2_44[123]}
   );
   gpc1_1 gpc8082 (
      {stage1_44[255]},
      {stage2_44[124]}
   );
   gpc1_1 gpc8083 (
      {stage1_44[256]},
      {stage2_44[125]}
   );
   gpc1_1 gpc8084 (
      {stage1_44[257]},
      {stage2_44[126]}
   );
   gpc1_1 gpc8085 (
      {stage1_44[258]},
      {stage2_44[127]}
   );
   gpc1_1 gpc8086 (
      {stage1_44[259]},
      {stage2_44[128]}
   );
   gpc1_1 gpc8087 (
      {stage1_44[260]},
      {stage2_44[129]}
   );
   gpc1_1 gpc8088 (
      {stage1_44[261]},
      {stage2_44[130]}
   );
   gpc1_1 gpc8089 (
      {stage1_44[262]},
      {stage2_44[131]}
   );
   gpc1_1 gpc8090 (
      {stage1_44[263]},
      {stage2_44[132]}
   );
   gpc1_1 gpc8091 (
      {stage1_44[264]},
      {stage2_44[133]}
   );
   gpc1_1 gpc8092 (
      {stage1_44[265]},
      {stage2_44[134]}
   );
   gpc1_1 gpc8093 (
      {stage1_44[266]},
      {stage2_44[135]}
   );
   gpc1_1 gpc8094 (
      {stage1_44[267]},
      {stage2_44[136]}
   );
   gpc1_1 gpc8095 (
      {stage1_44[268]},
      {stage2_44[137]}
   );
   gpc1_1 gpc8096 (
      {stage1_45[157]},
      {stage2_45[100]}
   );
   gpc1_1 gpc8097 (
      {stage1_45[158]},
      {stage2_45[101]}
   );
   gpc1_1 gpc8098 (
      {stage1_45[159]},
      {stage2_45[102]}
   );
   gpc1_1 gpc8099 (
      {stage1_45[160]},
      {stage2_45[103]}
   );
   gpc1_1 gpc8100 (
      {stage1_45[161]},
      {stage2_45[104]}
   );
   gpc1_1 gpc8101 (
      {stage1_45[162]},
      {stage2_45[105]}
   );
   gpc1_1 gpc8102 (
      {stage1_45[163]},
      {stage2_45[106]}
   );
   gpc1_1 gpc8103 (
      {stage1_45[164]},
      {stage2_45[107]}
   );
   gpc1_1 gpc8104 (
      {stage1_45[165]},
      {stage2_45[108]}
   );
   gpc1_1 gpc8105 (
      {stage1_45[166]},
      {stage2_45[109]}
   );
   gpc1_1 gpc8106 (
      {stage1_45[167]},
      {stage2_45[110]}
   );
   gpc1_1 gpc8107 (
      {stage1_45[168]},
      {stage2_45[111]}
   );
   gpc1_1 gpc8108 (
      {stage1_45[169]},
      {stage2_45[112]}
   );
   gpc1_1 gpc8109 (
      {stage1_45[170]},
      {stage2_45[113]}
   );
   gpc1_1 gpc8110 (
      {stage1_45[171]},
      {stage2_45[114]}
   );
   gpc1_1 gpc8111 (
      {stage1_45[172]},
      {stage2_45[115]}
   );
   gpc1_1 gpc8112 (
      {stage1_45[173]},
      {stage2_45[116]}
   );
   gpc1_1 gpc8113 (
      {stage1_45[174]},
      {stage2_45[117]}
   );
   gpc1_1 gpc8114 (
      {stage1_45[175]},
      {stage2_45[118]}
   );
   gpc1_1 gpc8115 (
      {stage1_45[176]},
      {stage2_45[119]}
   );
   gpc1_1 gpc8116 (
      {stage1_45[177]},
      {stage2_45[120]}
   );
   gpc1_1 gpc8117 (
      {stage1_45[178]},
      {stage2_45[121]}
   );
   gpc1_1 gpc8118 (
      {stage1_45[179]},
      {stage2_45[122]}
   );
   gpc1_1 gpc8119 (
      {stage1_45[180]},
      {stage2_45[123]}
   );
   gpc1_1 gpc8120 (
      {stage1_45[181]},
      {stage2_45[124]}
   );
   gpc1_1 gpc8121 (
      {stage1_45[182]},
      {stage2_45[125]}
   );
   gpc1_1 gpc8122 (
      {stage1_45[183]},
      {stage2_45[126]}
   );
   gpc1_1 gpc8123 (
      {stage1_45[184]},
      {stage2_45[127]}
   );
   gpc1_1 gpc8124 (
      {stage1_45[185]},
      {stage2_45[128]}
   );
   gpc1_1 gpc8125 (
      {stage1_45[186]},
      {stage2_45[129]}
   );
   gpc1_1 gpc8126 (
      {stage1_45[187]},
      {stage2_45[130]}
   );
   gpc1_1 gpc8127 (
      {stage1_45[188]},
      {stage2_45[131]}
   );
   gpc1_1 gpc8128 (
      {stage1_46[285]},
      {stage2_46[78]}
   );
   gpc1_1 gpc8129 (
      {stage1_46[286]},
      {stage2_46[79]}
   );
   gpc1_1 gpc8130 (
      {stage1_46[287]},
      {stage2_46[80]}
   );
   gpc1_1 gpc8131 (
      {stage1_46[288]},
      {stage2_46[81]}
   );
   gpc1_1 gpc8132 (
      {stage1_46[289]},
      {stage2_46[82]}
   );
   gpc1_1 gpc8133 (
      {stage1_46[290]},
      {stage2_46[83]}
   );
   gpc1_1 gpc8134 (
      {stage1_46[291]},
      {stage2_46[84]}
   );
   gpc1_1 gpc8135 (
      {stage1_46[292]},
      {stage2_46[85]}
   );
   gpc1_1 gpc8136 (
      {stage1_46[293]},
      {stage2_46[86]}
   );
   gpc1_1 gpc8137 (
      {stage1_46[294]},
      {stage2_46[87]}
   );
   gpc1_1 gpc8138 (
      {stage1_46[295]},
      {stage2_46[88]}
   );
   gpc1_1 gpc8139 (
      {stage1_46[296]},
      {stage2_46[89]}
   );
   gpc1_1 gpc8140 (
      {stage1_46[297]},
      {stage2_46[90]}
   );
   gpc1_1 gpc8141 (
      {stage1_46[298]},
      {stage2_46[91]}
   );
   gpc1_1 gpc8142 (
      {stage1_46[299]},
      {stage2_46[92]}
   );
   gpc1_1 gpc8143 (
      {stage1_47[270]},
      {stage2_47[100]}
   );
   gpc1_1 gpc8144 (
      {stage1_47[271]},
      {stage2_47[101]}
   );
   gpc1_1 gpc8145 (
      {stage1_47[272]},
      {stage2_47[102]}
   );
   gpc1_1 gpc8146 (
      {stage1_47[273]},
      {stage2_47[103]}
   );
   gpc1_1 gpc8147 (
      {stage1_47[274]},
      {stage2_47[104]}
   );
   gpc1_1 gpc8148 (
      {stage1_47[275]},
      {stage2_47[105]}
   );
   gpc1_1 gpc8149 (
      {stage1_47[276]},
      {stage2_47[106]}
   );
   gpc1_1 gpc8150 (
      {stage1_47[277]},
      {stage2_47[107]}
   );
   gpc1_1 gpc8151 (
      {stage1_48[166]},
      {stage2_48[109]}
   );
   gpc1_1 gpc8152 (
      {stage1_48[167]},
      {stage2_48[110]}
   );
   gpc1_1 gpc8153 (
      {stage1_48[168]},
      {stage2_48[111]}
   );
   gpc1_1 gpc8154 (
      {stage1_48[169]},
      {stage2_48[112]}
   );
   gpc1_1 gpc8155 (
      {stage1_48[170]},
      {stage2_48[113]}
   );
   gpc1_1 gpc8156 (
      {stage1_48[171]},
      {stage2_48[114]}
   );
   gpc1_1 gpc8157 (
      {stage1_48[172]},
      {stage2_48[115]}
   );
   gpc1_1 gpc8158 (
      {stage1_48[173]},
      {stage2_48[116]}
   );
   gpc1_1 gpc8159 (
      {stage1_48[174]},
      {stage2_48[117]}
   );
   gpc1_1 gpc8160 (
      {stage1_48[175]},
      {stage2_48[118]}
   );
   gpc1_1 gpc8161 (
      {stage1_48[176]},
      {stage2_48[119]}
   );
   gpc1_1 gpc8162 (
      {stage1_48[177]},
      {stage2_48[120]}
   );
   gpc1_1 gpc8163 (
      {stage1_48[178]},
      {stage2_48[121]}
   );
   gpc1_1 gpc8164 (
      {stage1_48[179]},
      {stage2_48[122]}
   );
   gpc1_1 gpc8165 (
      {stage1_48[180]},
      {stage2_48[123]}
   );
   gpc1_1 gpc8166 (
      {stage1_48[181]},
      {stage2_48[124]}
   );
   gpc1_1 gpc8167 (
      {stage1_48[182]},
      {stage2_48[125]}
   );
   gpc1_1 gpc8168 (
      {stage1_48[183]},
      {stage2_48[126]}
   );
   gpc1_1 gpc8169 (
      {stage1_48[184]},
      {stage2_48[127]}
   );
   gpc1_1 gpc8170 (
      {stage1_48[185]},
      {stage2_48[128]}
   );
   gpc1_1 gpc8171 (
      {stage1_48[186]},
      {stage2_48[129]}
   );
   gpc1_1 gpc8172 (
      {stage1_48[187]},
      {stage2_48[130]}
   );
   gpc1_1 gpc8173 (
      {stage1_48[188]},
      {stage2_48[131]}
   );
   gpc1_1 gpc8174 (
      {stage1_48[189]},
      {stage2_48[132]}
   );
   gpc1_1 gpc8175 (
      {stage1_48[190]},
      {stage2_48[133]}
   );
   gpc1_1 gpc8176 (
      {stage1_48[191]},
      {stage2_48[134]}
   );
   gpc1_1 gpc8177 (
      {stage1_48[192]},
      {stage2_48[135]}
   );
   gpc1_1 gpc8178 (
      {stage1_48[193]},
      {stage2_48[136]}
   );
   gpc1_1 gpc8179 (
      {stage1_48[194]},
      {stage2_48[137]}
   );
   gpc1_1 gpc8180 (
      {stage1_48[195]},
      {stage2_48[138]}
   );
   gpc1_1 gpc8181 (
      {stage1_48[196]},
      {stage2_48[139]}
   );
   gpc1_1 gpc8182 (
      {stage1_48[197]},
      {stage2_48[140]}
   );
   gpc1_1 gpc8183 (
      {stage1_48[198]},
      {stage2_48[141]}
   );
   gpc1_1 gpc8184 (
      {stage1_48[199]},
      {stage2_48[142]}
   );
   gpc1_1 gpc8185 (
      {stage1_48[200]},
      {stage2_48[143]}
   );
   gpc1_1 gpc8186 (
      {stage1_48[201]},
      {stage2_48[144]}
   );
   gpc1_1 gpc8187 (
      {stage1_48[202]},
      {stage2_48[145]}
   );
   gpc1_1 gpc8188 (
      {stage1_48[203]},
      {stage2_48[146]}
   );
   gpc1_1 gpc8189 (
      {stage1_48[204]},
      {stage2_48[147]}
   );
   gpc1_1 gpc8190 (
      {stage1_48[205]},
      {stage2_48[148]}
   );
   gpc1_1 gpc8191 (
      {stage1_48[206]},
      {stage2_48[149]}
   );
   gpc1_1 gpc8192 (
      {stage1_48[207]},
      {stage2_48[150]}
   );
   gpc1_1 gpc8193 (
      {stage1_48[208]},
      {stage2_48[151]}
   );
   gpc1_1 gpc8194 (
      {stage1_48[209]},
      {stage2_48[152]}
   );
   gpc1_1 gpc8195 (
      {stage1_48[210]},
      {stage2_48[153]}
   );
   gpc1_1 gpc8196 (
      {stage1_49[203]},
      {stage2_49[77]}
   );
   gpc1_1 gpc8197 (
      {stage1_49[204]},
      {stage2_49[78]}
   );
   gpc1_1 gpc8198 (
      {stage1_49[205]},
      {stage2_49[79]}
   );
   gpc1_1 gpc8199 (
      {stage1_49[206]},
      {stage2_49[80]}
   );
   gpc1_1 gpc8200 (
      {stage1_49[207]},
      {stage2_49[81]}
   );
   gpc1_1 gpc8201 (
      {stage1_49[208]},
      {stage2_49[82]}
   );
   gpc1_1 gpc8202 (
      {stage1_49[209]},
      {stage2_49[83]}
   );
   gpc1_1 gpc8203 (
      {stage1_49[210]},
      {stage2_49[84]}
   );
   gpc1_1 gpc8204 (
      {stage1_49[211]},
      {stage2_49[85]}
   );
   gpc1_1 gpc8205 (
      {stage1_49[212]},
      {stage2_49[86]}
   );
   gpc1_1 gpc8206 (
      {stage1_49[213]},
      {stage2_49[87]}
   );
   gpc1_1 gpc8207 (
      {stage1_49[214]},
      {stage2_49[88]}
   );
   gpc1_1 gpc8208 (
      {stage1_49[215]},
      {stage2_49[89]}
   );
   gpc1_1 gpc8209 (
      {stage1_49[216]},
      {stage2_49[90]}
   );
   gpc1_1 gpc8210 (
      {stage1_49[217]},
      {stage2_49[91]}
   );
   gpc1_1 gpc8211 (
      {stage1_49[218]},
      {stage2_49[92]}
   );
   gpc1_1 gpc8212 (
      {stage1_49[219]},
      {stage2_49[93]}
   );
   gpc1_1 gpc8213 (
      {stage1_49[220]},
      {stage2_49[94]}
   );
   gpc1_1 gpc8214 (
      {stage1_49[221]},
      {stage2_49[95]}
   );
   gpc1_1 gpc8215 (
      {stage1_49[222]},
      {stage2_49[96]}
   );
   gpc1_1 gpc8216 (
      {stage1_49[223]},
      {stage2_49[97]}
   );
   gpc1_1 gpc8217 (
      {stage1_49[224]},
      {stage2_49[98]}
   );
   gpc1_1 gpc8218 (
      {stage1_49[225]},
      {stage2_49[99]}
   );
   gpc1_1 gpc8219 (
      {stage1_49[226]},
      {stage2_49[100]}
   );
   gpc1_1 gpc8220 (
      {stage1_49[227]},
      {stage2_49[101]}
   );
   gpc1_1 gpc8221 (
      {stage1_49[228]},
      {stage2_49[102]}
   );
   gpc1_1 gpc8222 (
      {stage1_49[229]},
      {stage2_49[103]}
   );
   gpc1_1 gpc8223 (
      {stage1_49[230]},
      {stage2_49[104]}
   );
   gpc1_1 gpc8224 (
      {stage1_49[231]},
      {stage2_49[105]}
   );
   gpc1_1 gpc8225 (
      {stage1_49[232]},
      {stage2_49[106]}
   );
   gpc1_1 gpc8226 (
      {stage1_49[233]},
      {stage2_49[107]}
   );
   gpc1_1 gpc8227 (
      {stage1_49[234]},
      {stage2_49[108]}
   );
   gpc1_1 gpc8228 (
      {stage1_49[235]},
      {stage2_49[109]}
   );
   gpc1_1 gpc8229 (
      {stage1_49[236]},
      {stage2_49[110]}
   );
   gpc1_1 gpc8230 (
      {stage1_49[237]},
      {stage2_49[111]}
   );
   gpc1_1 gpc8231 (
      {stage1_49[238]},
      {stage2_49[112]}
   );
   gpc1_1 gpc8232 (
      {stage1_49[239]},
      {stage2_49[113]}
   );
   gpc1_1 gpc8233 (
      {stage1_49[240]},
      {stage2_49[114]}
   );
   gpc1_1 gpc8234 (
      {stage1_49[241]},
      {stage2_49[115]}
   );
   gpc1_1 gpc8235 (
      {stage1_50[134]},
      {stage2_50[70]}
   );
   gpc1_1 gpc8236 (
      {stage1_50[135]},
      {stage2_50[71]}
   );
   gpc1_1 gpc8237 (
      {stage1_50[136]},
      {stage2_50[72]}
   );
   gpc1_1 gpc8238 (
      {stage1_50[137]},
      {stage2_50[73]}
   );
   gpc1_1 gpc8239 (
      {stage1_50[138]},
      {stage2_50[74]}
   );
   gpc1_1 gpc8240 (
      {stage1_50[139]},
      {stage2_50[75]}
   );
   gpc1_1 gpc8241 (
      {stage1_50[140]},
      {stage2_50[76]}
   );
   gpc1_1 gpc8242 (
      {stage1_50[141]},
      {stage2_50[77]}
   );
   gpc1_1 gpc8243 (
      {stage1_50[142]},
      {stage2_50[78]}
   );
   gpc1_1 gpc8244 (
      {stage1_50[143]},
      {stage2_50[79]}
   );
   gpc1_1 gpc8245 (
      {stage1_50[144]},
      {stage2_50[80]}
   );
   gpc1_1 gpc8246 (
      {stage1_50[145]},
      {stage2_50[81]}
   );
   gpc1_1 gpc8247 (
      {stage1_50[146]},
      {stage2_50[82]}
   );
   gpc1_1 gpc8248 (
      {stage1_50[147]},
      {stage2_50[83]}
   );
   gpc1_1 gpc8249 (
      {stage1_50[148]},
      {stage2_50[84]}
   );
   gpc1_1 gpc8250 (
      {stage1_50[149]},
      {stage2_50[85]}
   );
   gpc1_1 gpc8251 (
      {stage1_50[150]},
      {stage2_50[86]}
   );
   gpc1_1 gpc8252 (
      {stage1_50[151]},
      {stage2_50[87]}
   );
   gpc1_1 gpc8253 (
      {stage1_50[152]},
      {stage2_50[88]}
   );
   gpc1_1 gpc8254 (
      {stage1_50[153]},
      {stage2_50[89]}
   );
   gpc1_1 gpc8255 (
      {stage1_50[154]},
      {stage2_50[90]}
   );
   gpc1_1 gpc8256 (
      {stage1_50[155]},
      {stage2_50[91]}
   );
   gpc1_1 gpc8257 (
      {stage1_50[156]},
      {stage2_50[92]}
   );
   gpc1_1 gpc8258 (
      {stage1_50[157]},
      {stage2_50[93]}
   );
   gpc1_1 gpc8259 (
      {stage1_50[158]},
      {stage2_50[94]}
   );
   gpc1_1 gpc8260 (
      {stage1_50[159]},
      {stage2_50[95]}
   );
   gpc1_1 gpc8261 (
      {stage1_50[160]},
      {stage2_50[96]}
   );
   gpc1_1 gpc8262 (
      {stage1_50[161]},
      {stage2_50[97]}
   );
   gpc1_1 gpc8263 (
      {stage1_50[162]},
      {stage2_50[98]}
   );
   gpc1_1 gpc8264 (
      {stage1_50[163]},
      {stage2_50[99]}
   );
   gpc1_1 gpc8265 (
      {stage1_50[164]},
      {stage2_50[100]}
   );
   gpc1_1 gpc8266 (
      {stage1_50[165]},
      {stage2_50[101]}
   );
   gpc1_1 gpc8267 (
      {stage1_50[166]},
      {stage2_50[102]}
   );
   gpc1_1 gpc8268 (
      {stage1_50[167]},
      {stage2_50[103]}
   );
   gpc1_1 gpc8269 (
      {stage1_50[168]},
      {stage2_50[104]}
   );
   gpc1_1 gpc8270 (
      {stage1_50[169]},
      {stage2_50[105]}
   );
   gpc1_1 gpc8271 (
      {stage1_50[170]},
      {stage2_50[106]}
   );
   gpc1_1 gpc8272 (
      {stage1_50[171]},
      {stage2_50[107]}
   );
   gpc1_1 gpc8273 (
      {stage1_50[172]},
      {stage2_50[108]}
   );
   gpc1_1 gpc8274 (
      {stage1_50[173]},
      {stage2_50[109]}
   );
   gpc1_1 gpc8275 (
      {stage1_50[174]},
      {stage2_50[110]}
   );
   gpc1_1 gpc8276 (
      {stage1_50[175]},
      {stage2_50[111]}
   );
   gpc1_1 gpc8277 (
      {stage1_50[176]},
      {stage2_50[112]}
   );
   gpc1_1 gpc8278 (
      {stage1_50[177]},
      {stage2_50[113]}
   );
   gpc1_1 gpc8279 (
      {stage1_50[178]},
      {stage2_50[114]}
   );
   gpc1_1 gpc8280 (
      {stage1_50[179]},
      {stage2_50[115]}
   );
   gpc1_1 gpc8281 (
      {stage1_50[180]},
      {stage2_50[116]}
   );
   gpc1_1 gpc8282 (
      {stage1_50[181]},
      {stage2_50[117]}
   );
   gpc1_1 gpc8283 (
      {stage1_50[182]},
      {stage2_50[118]}
   );
   gpc1_1 gpc8284 (
      {stage1_50[183]},
      {stage2_50[119]}
   );
   gpc1_1 gpc8285 (
      {stage1_50[184]},
      {stage2_50[120]}
   );
   gpc1_1 gpc8286 (
      {stage1_50[185]},
      {stage2_50[121]}
   );
   gpc1_1 gpc8287 (
      {stage1_50[186]},
      {stage2_50[122]}
   );
   gpc1_1 gpc8288 (
      {stage1_50[187]},
      {stage2_50[123]}
   );
   gpc1_1 gpc8289 (
      {stage1_50[188]},
      {stage2_50[124]}
   );
   gpc1_1 gpc8290 (
      {stage1_50[189]},
      {stage2_50[125]}
   );
   gpc1_1 gpc8291 (
      {stage1_50[190]},
      {stage2_50[126]}
   );
   gpc1_1 gpc8292 (
      {stage1_50[191]},
      {stage2_50[127]}
   );
   gpc1_1 gpc8293 (
      {stage1_50[192]},
      {stage2_50[128]}
   );
   gpc1_1 gpc8294 (
      {stage1_50[193]},
      {stage2_50[129]}
   );
   gpc1_1 gpc8295 (
      {stage1_50[194]},
      {stage2_50[130]}
   );
   gpc1_1 gpc8296 (
      {stage1_50[195]},
      {stage2_50[131]}
   );
   gpc1_1 gpc8297 (
      {stage1_50[196]},
      {stage2_50[132]}
   );
   gpc1_1 gpc8298 (
      {stage1_50[197]},
      {stage2_50[133]}
   );
   gpc1_1 gpc8299 (
      {stage1_50[198]},
      {stage2_50[134]}
   );
   gpc1_1 gpc8300 (
      {stage1_50[199]},
      {stage2_50[135]}
   );
   gpc1_1 gpc8301 (
      {stage1_50[200]},
      {stage2_50[136]}
   );
   gpc1_1 gpc8302 (
      {stage1_50[201]},
      {stage2_50[137]}
   );
   gpc1_1 gpc8303 (
      {stage1_50[202]},
      {stage2_50[138]}
   );
   gpc1_1 gpc8304 (
      {stage1_50[203]},
      {stage2_50[139]}
   );
   gpc1_1 gpc8305 (
      {stage1_50[204]},
      {stage2_50[140]}
   );
   gpc1_1 gpc8306 (
      {stage1_50[205]},
      {stage2_50[141]}
   );
   gpc1_1 gpc8307 (
      {stage1_50[206]},
      {stage2_50[142]}
   );
   gpc1_1 gpc8308 (
      {stage1_50[207]},
      {stage2_50[143]}
   );
   gpc1_1 gpc8309 (
      {stage1_50[208]},
      {stage2_50[144]}
   );
   gpc1_1 gpc8310 (
      {stage1_50[209]},
      {stage2_50[145]}
   );
   gpc1_1 gpc8311 (
      {stage1_50[210]},
      {stage2_50[146]}
   );
   gpc1_1 gpc8312 (
      {stage1_50[211]},
      {stage2_50[147]}
   );
   gpc1_1 gpc8313 (
      {stage1_50[212]},
      {stage2_50[148]}
   );
   gpc1_1 gpc8314 (
      {stage1_50[213]},
      {stage2_50[149]}
   );
   gpc1_1 gpc8315 (
      {stage1_50[214]},
      {stage2_50[150]}
   );
   gpc1_1 gpc8316 (
      {stage1_50[215]},
      {stage2_50[151]}
   );
   gpc1_1 gpc8317 (
      {stage1_50[216]},
      {stage2_50[152]}
   );
   gpc1_1 gpc8318 (
      {stage1_51[224]},
      {stage2_51[85]}
   );
   gpc1_1 gpc8319 (
      {stage1_51[225]},
      {stage2_51[86]}
   );
   gpc1_1 gpc8320 (
      {stage1_51[226]},
      {stage2_51[87]}
   );
   gpc1_1 gpc8321 (
      {stage1_52[269]},
      {stage2_52[93]}
   );
   gpc1_1 gpc8322 (
      {stage1_52[270]},
      {stage2_52[94]}
   );
   gpc1_1 gpc8323 (
      {stage1_52[271]},
      {stage2_52[95]}
   );
   gpc1_1 gpc8324 (
      {stage1_52[272]},
      {stage2_52[96]}
   );
   gpc1_1 gpc8325 (
      {stage1_52[273]},
      {stage2_52[97]}
   );
   gpc1_1 gpc8326 (
      {stage1_52[274]},
      {stage2_52[98]}
   );
   gpc1_1 gpc8327 (
      {stage1_52[275]},
      {stage2_52[99]}
   );
   gpc1_1 gpc8328 (
      {stage1_52[276]},
      {stage2_52[100]}
   );
   gpc1_1 gpc8329 (
      {stage1_52[277]},
      {stage2_52[101]}
   );
   gpc1_1 gpc8330 (
      {stage1_52[278]},
      {stage2_52[102]}
   );
   gpc1_1 gpc8331 (
      {stage1_52[279]},
      {stage2_52[103]}
   );
   gpc1_1 gpc8332 (
      {stage1_52[280]},
      {stage2_52[104]}
   );
   gpc1_1 gpc8333 (
      {stage1_52[281]},
      {stage2_52[105]}
   );
   gpc1_1 gpc8334 (
      {stage1_52[282]},
      {stage2_52[106]}
   );
   gpc1_1 gpc8335 (
      {stage1_52[283]},
      {stage2_52[107]}
   );
   gpc1_1 gpc8336 (
      {stage1_52[284]},
      {stage2_52[108]}
   );
   gpc1_1 gpc8337 (
      {stage1_52[285]},
      {stage2_52[109]}
   );
   gpc1_1 gpc8338 (
      {stage1_52[286]},
      {stage2_52[110]}
   );
   gpc1_1 gpc8339 (
      {stage1_52[287]},
      {stage2_52[111]}
   );
   gpc1_1 gpc8340 (
      {stage1_52[288]},
      {stage2_52[112]}
   );
   gpc1_1 gpc8341 (
      {stage1_52[289]},
      {stage2_52[113]}
   );
   gpc1_1 gpc8342 (
      {stage1_52[290]},
      {stage2_52[114]}
   );
   gpc1_1 gpc8343 (
      {stage1_52[291]},
      {stage2_52[115]}
   );
   gpc1_1 gpc8344 (
      {stage1_52[292]},
      {stage2_52[116]}
   );
   gpc1_1 gpc8345 (
      {stage1_52[293]},
      {stage2_52[117]}
   );
   gpc1_1 gpc8346 (
      {stage1_52[294]},
      {stage2_52[118]}
   );
   gpc1_1 gpc8347 (
      {stage1_52[295]},
      {stage2_52[119]}
   );
   gpc1_1 gpc8348 (
      {stage1_52[296]},
      {stage2_52[120]}
   );
   gpc1_1 gpc8349 (
      {stage1_52[297]},
      {stage2_52[121]}
   );
   gpc1_1 gpc8350 (
      {stage1_52[298]},
      {stage2_52[122]}
   );
   gpc1_1 gpc8351 (
      {stage1_52[299]},
      {stage2_52[123]}
   );
   gpc1_1 gpc8352 (
      {stage1_52[300]},
      {stage2_52[124]}
   );
   gpc1_1 gpc8353 (
      {stage1_52[301]},
      {stage2_52[125]}
   );
   gpc1_1 gpc8354 (
      {stage1_52[302]},
      {stage2_52[126]}
   );
   gpc1_1 gpc8355 (
      {stage1_52[303]},
      {stage2_52[127]}
   );
   gpc1_1 gpc8356 (
      {stage1_53[173]},
      {stage2_53[83]}
   );
   gpc1_1 gpc8357 (
      {stage1_53[174]},
      {stage2_53[84]}
   );
   gpc1_1 gpc8358 (
      {stage1_53[175]},
      {stage2_53[85]}
   );
   gpc1_1 gpc8359 (
      {stage1_53[176]},
      {stage2_53[86]}
   );
   gpc1_1 gpc8360 (
      {stage1_53[177]},
      {stage2_53[87]}
   );
   gpc1_1 gpc8361 (
      {stage1_53[178]},
      {stage2_53[88]}
   );
   gpc1_1 gpc8362 (
      {stage1_53[179]},
      {stage2_53[89]}
   );
   gpc1_1 gpc8363 (
      {stage1_53[180]},
      {stage2_53[90]}
   );
   gpc1_1 gpc8364 (
      {stage1_53[181]},
      {stage2_53[91]}
   );
   gpc1_1 gpc8365 (
      {stage1_53[182]},
      {stage2_53[92]}
   );
   gpc1_1 gpc8366 (
      {stage1_53[183]},
      {stage2_53[93]}
   );
   gpc1_1 gpc8367 (
      {stage1_53[184]},
      {stage2_53[94]}
   );
   gpc1_1 gpc8368 (
      {stage1_53[185]},
      {stage2_53[95]}
   );
   gpc1_1 gpc8369 (
      {stage1_53[186]},
      {stage2_53[96]}
   );
   gpc1_1 gpc8370 (
      {stage1_54[216]},
      {stage2_54[77]}
   );
   gpc1_1 gpc8371 (
      {stage1_54[217]},
      {stage2_54[78]}
   );
   gpc1_1 gpc8372 (
      {stage1_54[218]},
      {stage2_54[79]}
   );
   gpc1_1 gpc8373 (
      {stage1_54[219]},
      {stage2_54[80]}
   );
   gpc1_1 gpc8374 (
      {stage1_54[220]},
      {stage2_54[81]}
   );
   gpc1_1 gpc8375 (
      {stage1_54[221]},
      {stage2_54[82]}
   );
   gpc1_1 gpc8376 (
      {stage1_54[222]},
      {stage2_54[83]}
   );
   gpc1_1 gpc8377 (
      {stage1_54[223]},
      {stage2_54[84]}
   );
   gpc1_1 gpc8378 (
      {stage1_54[224]},
      {stage2_54[85]}
   );
   gpc1_1 gpc8379 (
      {stage1_54[225]},
      {stage2_54[86]}
   );
   gpc1_1 gpc8380 (
      {stage1_54[226]},
      {stage2_54[87]}
   );
   gpc1_1 gpc8381 (
      {stage1_54[227]},
      {stage2_54[88]}
   );
   gpc1_1 gpc8382 (
      {stage1_54[228]},
      {stage2_54[89]}
   );
   gpc1_1 gpc8383 (
      {stage1_54[229]},
      {stage2_54[90]}
   );
   gpc1_1 gpc8384 (
      {stage1_54[230]},
      {stage2_54[91]}
   );
   gpc1_1 gpc8385 (
      {stage1_54[231]},
      {stage2_54[92]}
   );
   gpc1_1 gpc8386 (
      {stage1_54[232]},
      {stage2_54[93]}
   );
   gpc1_1 gpc8387 (
      {stage1_54[233]},
      {stage2_54[94]}
   );
   gpc1_1 gpc8388 (
      {stage1_54[234]},
      {stage2_54[95]}
   );
   gpc1_1 gpc8389 (
      {stage1_54[235]},
      {stage2_54[96]}
   );
   gpc1_1 gpc8390 (
      {stage1_54[236]},
      {stage2_54[97]}
   );
   gpc1_1 gpc8391 (
      {stage1_54[237]},
      {stage2_54[98]}
   );
   gpc1_1 gpc8392 (
      {stage1_54[238]},
      {stage2_54[99]}
   );
   gpc1_1 gpc8393 (
      {stage1_54[239]},
      {stage2_54[100]}
   );
   gpc1_1 gpc8394 (
      {stage1_54[240]},
      {stage2_54[101]}
   );
   gpc1_1 gpc8395 (
      {stage1_54[241]},
      {stage2_54[102]}
   );
   gpc1_1 gpc8396 (
      {stage1_54[242]},
      {stage2_54[103]}
   );
   gpc1_1 gpc8397 (
      {stage1_54[243]},
      {stage2_54[104]}
   );
   gpc1_1 gpc8398 (
      {stage1_54[244]},
      {stage2_54[105]}
   );
   gpc1_1 gpc8399 (
      {stage1_54[245]},
      {stage2_54[106]}
   );
   gpc1_1 gpc8400 (
      {stage1_54[246]},
      {stage2_54[107]}
   );
   gpc1_1 gpc8401 (
      {stage1_54[247]},
      {stage2_54[108]}
   );
   gpc1_1 gpc8402 (
      {stage1_54[248]},
      {stage2_54[109]}
   );
   gpc1_1 gpc8403 (
      {stage1_54[249]},
      {stage2_54[110]}
   );
   gpc1_1 gpc8404 (
      {stage1_54[250]},
      {stage2_54[111]}
   );
   gpc1_1 gpc8405 (
      {stage1_54[251]},
      {stage2_54[112]}
   );
   gpc1_1 gpc8406 (
      {stage1_54[252]},
      {stage2_54[113]}
   );
   gpc1_1 gpc8407 (
      {stage1_54[253]},
      {stage2_54[114]}
   );
   gpc1_1 gpc8408 (
      {stage1_54[254]},
      {stage2_54[115]}
   );
   gpc1_1 gpc8409 (
      {stage1_54[255]},
      {stage2_54[116]}
   );
   gpc1_1 gpc8410 (
      {stage1_54[256]},
      {stage2_54[117]}
   );
   gpc1_1 gpc8411 (
      {stage1_54[257]},
      {stage2_54[118]}
   );
   gpc1_1 gpc8412 (
      {stage1_54[258]},
      {stage2_54[119]}
   );
   gpc1_1 gpc8413 (
      {stage1_54[259]},
      {stage2_54[120]}
   );
   gpc1_1 gpc8414 (
      {stage1_54[260]},
      {stage2_54[121]}
   );
   gpc1_1 gpc8415 (
      {stage1_54[261]},
      {stage2_54[122]}
   );
   gpc1_1 gpc8416 (
      {stage1_54[262]},
      {stage2_54[123]}
   );
   gpc1_1 gpc8417 (
      {stage1_55[219]},
      {stage2_55[104]}
   );
   gpc1_1 gpc8418 (
      {stage1_55[220]},
      {stage2_55[105]}
   );
   gpc1_1 gpc8419 (
      {stage1_55[221]},
      {stage2_55[106]}
   );
   gpc1_1 gpc8420 (
      {stage1_55[222]},
      {stage2_55[107]}
   );
   gpc1_1 gpc8421 (
      {stage1_55[223]},
      {stage2_55[108]}
   );
   gpc1_1 gpc8422 (
      {stage1_55[224]},
      {stage2_55[109]}
   );
   gpc1_1 gpc8423 (
      {stage1_55[225]},
      {stage2_55[110]}
   );
   gpc1_1 gpc8424 (
      {stage1_56[225]},
      {stage2_56[100]}
   );
   gpc1_1 gpc8425 (
      {stage1_56[226]},
      {stage2_56[101]}
   );
   gpc1_1 gpc8426 (
      {stage1_56[227]},
      {stage2_56[102]}
   );
   gpc1_1 gpc8427 (
      {stage1_56[228]},
      {stage2_56[103]}
   );
   gpc1_1 gpc8428 (
      {stage1_56[229]},
      {stage2_56[104]}
   );
   gpc1_1 gpc8429 (
      {stage1_56[230]},
      {stage2_56[105]}
   );
   gpc1_1 gpc8430 (
      {stage1_56[231]},
      {stage2_56[106]}
   );
   gpc1_1 gpc8431 (
      {stage1_56[232]},
      {stage2_56[107]}
   );
   gpc1_1 gpc8432 (
      {stage1_56[233]},
      {stage2_56[108]}
   );
   gpc1_1 gpc8433 (
      {stage1_56[234]},
      {stage2_56[109]}
   );
   gpc1_1 gpc8434 (
      {stage1_56[235]},
      {stage2_56[110]}
   );
   gpc1_1 gpc8435 (
      {stage1_56[236]},
      {stage2_56[111]}
   );
   gpc1_1 gpc8436 (
      {stage1_56[237]},
      {stage2_56[112]}
   );
   gpc1_1 gpc8437 (
      {stage1_56[238]},
      {stage2_56[113]}
   );
   gpc1_1 gpc8438 (
      {stage1_56[239]},
      {stage2_56[114]}
   );
   gpc1_1 gpc8439 (
      {stage1_56[240]},
      {stage2_56[115]}
   );
   gpc1_1 gpc8440 (
      {stage1_56[241]},
      {stage2_56[116]}
   );
   gpc1_1 gpc8441 (
      {stage1_56[242]},
      {stage2_56[117]}
   );
   gpc1_1 gpc8442 (
      {stage1_56[243]},
      {stage2_56[118]}
   );
   gpc1_1 gpc8443 (
      {stage1_56[244]},
      {stage2_56[119]}
   );
   gpc1_1 gpc8444 (
      {stage1_56[245]},
      {stage2_56[120]}
   );
   gpc1_1 gpc8445 (
      {stage1_56[246]},
      {stage2_56[121]}
   );
   gpc1_1 gpc8446 (
      {stage1_56[247]},
      {stage2_56[122]}
   );
   gpc1_1 gpc8447 (
      {stage1_56[248]},
      {stage2_56[123]}
   );
   gpc1_1 gpc8448 (
      {stage1_56[249]},
      {stage2_56[124]}
   );
   gpc1_1 gpc8449 (
      {stage1_56[250]},
      {stage2_56[125]}
   );
   gpc1_1 gpc8450 (
      {stage1_56[251]},
      {stage2_56[126]}
   );
   gpc1_1 gpc8451 (
      {stage1_56[252]},
      {stage2_56[127]}
   );
   gpc1_1 gpc8452 (
      {stage1_56[253]},
      {stage2_56[128]}
   );
   gpc1_1 gpc8453 (
      {stage1_56[254]},
      {stage2_56[129]}
   );
   gpc1_1 gpc8454 (
      {stage1_56[255]},
      {stage2_56[130]}
   );
   gpc1_1 gpc8455 (
      {stage1_56[256]},
      {stage2_56[131]}
   );
   gpc1_1 gpc8456 (
      {stage1_59[268]},
      {stage2_59[114]}
   );
   gpc1_1 gpc8457 (
      {stage1_59[269]},
      {stage2_59[115]}
   );
   gpc1_1 gpc8458 (
      {stage1_59[270]},
      {stage2_59[116]}
   );
   gpc1_1 gpc8459 (
      {stage1_59[271]},
      {stage2_59[117]}
   );
   gpc1_1 gpc8460 (
      {stage1_59[272]},
      {stage2_59[118]}
   );
   gpc1_1 gpc8461 (
      {stage1_59[273]},
      {stage2_59[119]}
   );
   gpc1_1 gpc8462 (
      {stage1_59[274]},
      {stage2_59[120]}
   );
   gpc1_1 gpc8463 (
      {stage1_59[275]},
      {stage2_59[121]}
   );
   gpc1_1 gpc8464 (
      {stage1_59[276]},
      {stage2_59[122]}
   );
   gpc1_1 gpc8465 (
      {stage1_59[277]},
      {stage2_59[123]}
   );
   gpc1_1 gpc8466 (
      {stage1_59[278]},
      {stage2_59[124]}
   );
   gpc1_1 gpc8467 (
      {stage1_59[279]},
      {stage2_59[125]}
   );
   gpc1_1 gpc8468 (
      {stage1_59[280]},
      {stage2_59[126]}
   );
   gpc1_1 gpc8469 (
      {stage1_59[281]},
      {stage2_59[127]}
   );
   gpc1_1 gpc8470 (
      {stage1_59[282]},
      {stage2_59[128]}
   );
   gpc1_1 gpc8471 (
      {stage1_59[283]},
      {stage2_59[129]}
   );
   gpc1_1 gpc8472 (
      {stage1_59[284]},
      {stage2_59[130]}
   );
   gpc1_1 gpc8473 (
      {stage1_59[285]},
      {stage2_59[131]}
   );
   gpc1_1 gpc8474 (
      {stage1_59[286]},
      {stage2_59[132]}
   );
   gpc1_1 gpc8475 (
      {stage1_59[287]},
      {stage2_59[133]}
   );
   gpc1_1 gpc8476 (
      {stage1_59[288]},
      {stage2_59[134]}
   );
   gpc1_1 gpc8477 (
      {stage1_59[289]},
      {stage2_59[135]}
   );
   gpc1_1 gpc8478 (
      {stage1_59[290]},
      {stage2_59[136]}
   );
   gpc1_1 gpc8479 (
      {stage1_59[291]},
      {stage2_59[137]}
   );
   gpc1_1 gpc8480 (
      {stage1_59[292]},
      {stage2_59[138]}
   );
   gpc1_1 gpc8481 (
      {stage1_59[293]},
      {stage2_59[139]}
   );
   gpc1_1 gpc8482 (
      {stage1_60[190]},
      {stage2_60[101]}
   );
   gpc1_1 gpc8483 (
      {stage1_60[191]},
      {stage2_60[102]}
   );
   gpc1_1 gpc8484 (
      {stage1_60[192]},
      {stage2_60[103]}
   );
   gpc1_1 gpc8485 (
      {stage1_60[193]},
      {stage2_60[104]}
   );
   gpc1_1 gpc8486 (
      {stage1_60[194]},
      {stage2_60[105]}
   );
   gpc1_1 gpc8487 (
      {stage1_60[195]},
      {stage2_60[106]}
   );
   gpc1_1 gpc8488 (
      {stage1_60[196]},
      {stage2_60[107]}
   );
   gpc1_1 gpc8489 (
      {stage1_60[197]},
      {stage2_60[108]}
   );
   gpc1_1 gpc8490 (
      {stage1_60[198]},
      {stage2_60[109]}
   );
   gpc1_1 gpc8491 (
      {stage1_60[199]},
      {stage2_60[110]}
   );
   gpc1_1 gpc8492 (
      {stage1_61[198]},
      {stage2_61[83]}
   );
   gpc1_1 gpc8493 (
      {stage1_61[199]},
      {stage2_61[84]}
   );
   gpc1_1 gpc8494 (
      {stage1_61[200]},
      {stage2_61[85]}
   );
   gpc1_1 gpc8495 (
      {stage1_61[201]},
      {stage2_61[86]}
   );
   gpc1_1 gpc8496 (
      {stage1_61[202]},
      {stage2_61[87]}
   );
   gpc1_1 gpc8497 (
      {stage1_61[203]},
      {stage2_61[88]}
   );
   gpc1_1 gpc8498 (
      {stage1_61[204]},
      {stage2_61[89]}
   );
   gpc1_1 gpc8499 (
      {stage1_61[205]},
      {stage2_61[90]}
   );
   gpc1_1 gpc8500 (
      {stage1_61[206]},
      {stage2_61[91]}
   );
   gpc1_1 gpc8501 (
      {stage1_61[207]},
      {stage2_61[92]}
   );
   gpc1_1 gpc8502 (
      {stage1_61[208]},
      {stage2_61[93]}
   );
   gpc1_1 gpc8503 (
      {stage1_61[209]},
      {stage2_61[94]}
   );
   gpc1_1 gpc8504 (
      {stage1_61[210]},
      {stage2_61[95]}
   );
   gpc1_1 gpc8505 (
      {stage1_61[211]},
      {stage2_61[96]}
   );
   gpc1_1 gpc8506 (
      {stage1_61[212]},
      {stage2_61[97]}
   );
   gpc1_1 gpc8507 (
      {stage1_61[213]},
      {stage2_61[98]}
   );
   gpc1_1 gpc8508 (
      {stage1_61[214]},
      {stage2_61[99]}
   );
   gpc1_1 gpc8509 (
      {stage1_61[215]},
      {stage2_61[100]}
   );
   gpc1_1 gpc8510 (
      {stage1_61[216]},
      {stage2_61[101]}
   );
   gpc1_1 gpc8511 (
      {stage1_62[346]},
      {stage2_62[118]}
   );
   gpc1_1 gpc8512 (
      {stage1_62[347]},
      {stage2_62[119]}
   );
   gpc1_1 gpc8513 (
      {stage1_62[348]},
      {stage2_62[120]}
   );
   gpc1_1 gpc8514 (
      {stage1_62[349]},
      {stage2_62[121]}
   );
   gpc1_1 gpc8515 (
      {stage1_62[350]},
      {stage2_62[122]}
   );
   gpc1_1 gpc8516 (
      {stage1_62[351]},
      {stage2_62[123]}
   );
   gpc1_1 gpc8517 (
      {stage1_62[352]},
      {stage2_62[124]}
   );
   gpc1_1 gpc8518 (
      {stage1_62[353]},
      {stage2_62[125]}
   );
   gpc1_1 gpc8519 (
      {stage1_62[354]},
      {stage2_62[126]}
   );
   gpc1_1 gpc8520 (
      {stage1_62[355]},
      {stage2_62[127]}
   );
   gpc1_1 gpc8521 (
      {stage1_62[356]},
      {stage2_62[128]}
   );
   gpc1_1 gpc8522 (
      {stage1_62[357]},
      {stage2_62[129]}
   );
   gpc1_1 gpc8523 (
      {stage1_62[358]},
      {stage2_62[130]}
   );
   gpc1_1 gpc8524 (
      {stage1_62[359]},
      {stage2_62[131]}
   );
   gpc1_1 gpc8525 (
      {stage1_62[360]},
      {stage2_62[132]}
   );
   gpc1_1 gpc8526 (
      {stage1_62[361]},
      {stage2_62[133]}
   );
   gpc1_1 gpc8527 (
      {stage1_62[362]},
      {stage2_62[134]}
   );
   gpc1_1 gpc8528 (
      {stage1_62[363]},
      {stage2_62[135]}
   );
   gpc1_1 gpc8529 (
      {stage1_62[364]},
      {stage2_62[136]}
   );
   gpc1_1 gpc8530 (
      {stage1_62[365]},
      {stage2_62[137]}
   );
   gpc1_1 gpc8531 (
      {stage1_62[366]},
      {stage2_62[138]}
   );
   gpc1_1 gpc8532 (
      {stage1_62[367]},
      {stage2_62[139]}
   );
   gpc1_1 gpc8533 (
      {stage1_62[368]},
      {stage2_62[140]}
   );
   gpc1_1 gpc8534 (
      {stage1_62[369]},
      {stage2_62[141]}
   );
   gpc1_1 gpc8535 (
      {stage1_62[370]},
      {stage2_62[142]}
   );
   gpc1_1 gpc8536 (
      {stage1_62[371]},
      {stage2_62[143]}
   );
   gpc1_1 gpc8537 (
      {stage1_62[372]},
      {stage2_62[144]}
   );
   gpc1_1 gpc8538 (
      {stage1_64[94]},
      {stage2_64[84]}
   );
   gpc1_1 gpc8539 (
      {stage1_64[95]},
      {stage2_64[85]}
   );
   gpc1_1 gpc8540 (
      {stage1_64[96]},
      {stage2_64[86]}
   );
   gpc1_1 gpc8541 (
      {stage1_64[97]},
      {stage2_64[87]}
   );
   gpc1_1 gpc8542 (
      {stage1_64[98]},
      {stage2_64[88]}
   );
   gpc1_1 gpc8543 (
      {stage1_64[99]},
      {stage2_64[89]}
   );
   gpc1_1 gpc8544 (
      {stage1_64[100]},
      {stage2_64[90]}
   );
   gpc1_1 gpc8545 (
      {stage1_64[101]},
      {stage2_64[91]}
   );
   gpc1_1 gpc8546 (
      {stage1_64[102]},
      {stage2_64[92]}
   );
   gpc1_1 gpc8547 (
      {stage1_64[103]},
      {stage2_64[93]}
   );
   gpc1_1 gpc8548 (
      {stage1_64[104]},
      {stage2_64[94]}
   );
   gpc1_1 gpc8549 (
      {stage1_64[105]},
      {stage2_64[95]}
   );
   gpc1_1 gpc8550 (
      {stage1_64[106]},
      {stage2_64[96]}
   );
   gpc1_1 gpc8551 (
      {stage1_64[107]},
      {stage2_64[97]}
   );
   gpc1_1 gpc8552 (
      {stage1_64[108]},
      {stage2_64[98]}
   );
   gpc1_1 gpc8553 (
      {stage1_64[109]},
      {stage2_64[99]}
   );
   gpc1_1 gpc8554 (
      {stage1_64[110]},
      {stage2_64[100]}
   );
   gpc1_1 gpc8555 (
      {stage1_64[111]},
      {stage2_64[101]}
   );
   gpc1_1 gpc8556 (
      {stage1_65[46]},
      {stage2_65[57]}
   );
   gpc1_1 gpc8557 (
      {stage1_65[47]},
      {stage2_65[58]}
   );
   gpc1_1 gpc8558 (
      {stage1_65[48]},
      {stage2_65[59]}
   );
   gpc1_1 gpc8559 (
      {stage1_65[49]},
      {stage2_65[60]}
   );
   gpc1_1 gpc8560 (
      {stage1_65[50]},
      {stage2_65[61]}
   );
   gpc1_1 gpc8561 (
      {stage1_65[51]},
      {stage2_65[62]}
   );
   gpc1_1 gpc8562 (
      {stage1_65[52]},
      {stage2_65[63]}
   );
   gpc1_1 gpc8563 (
      {stage1_65[53]},
      {stage2_65[64]}
   );
   gpc1_1 gpc8564 (
      {stage1_65[54]},
      {stage2_65[65]}
   );
   gpc1_1 gpc8565 (
      {stage1_65[55]},
      {stage2_65[66]}
   );
   gpc1_1 gpc8566 (
      {stage1_65[56]},
      {stage2_65[67]}
   );
   gpc1163_5 gpc8567 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc8568 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc8569 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[6]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc8570 (
      {stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18]},
      {stage2_1[7]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc615_5 gpc8571 (
      {stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_1[8]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc615_5 gpc8572 (
      {stage2_0[24], stage2_0[25], stage2_0[26], stage2_0[27], stage2_0[28]},
      {stage2_1[9]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1343_5 gpc8573 (
      {stage2_1[10], stage2_1[11], stage2_1[12]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[1], stage2_3[2], stage2_3[3]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc1343_5 gpc8574 (
      {stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[1]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc8575 (
      {stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc8576 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage3_6[0],stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9]}
   );
   gpc606_5 gpc8577 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49], stage2_2[50]},
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage3_6[1],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc8578 (
      {stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54], stage2_2[55], stage2_2[56]},
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage3_6[2],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc606_5 gpc8579 (
      {stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60], stage2_2[61], stage2_2[62]},
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage3_6[3],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc8580 (
      {stage2_2[63], stage2_2[64], stage2_2[65], stage2_2[66], stage2_2[67], stage2_2[68]},
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage3_6[4],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc8581 (
      {stage2_2[69], stage2_2[70], stage2_2[71], stage2_2[72], 1'b0, 1'b0},
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage3_6[5],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc207_4 gpc8582 (
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_5[0], stage2_5[1]},
      {stage3_6[6],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc207_4 gpc8583 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26]},
      {stage2_5[2], stage2_5[3]},
      {stage3_6[7],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc207_4 gpc8584 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_5[4], stage2_5[5]},
      {stage3_6[8],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc207_4 gpc8585 (
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40]},
      {stage2_5[6], stage2_5[7]},
      {stage3_6[9],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc207_4 gpc8586 (
      {stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[8], stage2_5[9]},
      {stage3_6[10],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc207_4 gpc8587 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_5[10], stage2_5[11]},
      {stage3_6[11],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc207_4 gpc8588 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_5[12], stage2_5[13]},
      {stage3_6[12],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc207_4 gpc8589 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_5[14], stage2_5[15]},
      {stage3_6[13],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc207_4 gpc8590 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75]},
      {stage2_5[16], stage2_5[17]},
      {stage3_6[14],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc207_4 gpc8591 (
      {stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_5[18], stage2_5[19]},
      {stage3_6[15],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc207_4 gpc8592 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_5[20], stage2_5[21]},
      {stage3_6[16],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc207_4 gpc8593 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96]},
      {stage2_5[22], stage2_5[23]},
      {stage3_6[17],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc207_4 gpc8594 (
      {stage2_3[97], stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103]},
      {stage2_5[24], stage2_5[25]},
      {stage3_6[18],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc207_4 gpc8595 (
      {stage2_3[104], stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109], stage2_3[110]},
      {stage2_5[26], stage2_5[27]},
      {stage3_6[19],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc207_4 gpc8596 (
      {stage2_3[111], stage2_3[112], stage2_3[113], stage2_3[114], stage2_3[115], stage2_3[116], stage2_3[117]},
      {stage2_5[28], stage2_5[29]},
      {stage3_6[20],stage3_5[23],stage3_4[29],stage3_3[29]}
   );
   gpc207_4 gpc8597 (
      {stage2_3[118], stage2_3[119], stage2_3[120], stage2_3[121], stage2_3[122], stage2_3[123], stage2_3[124]},
      {stage2_5[30], stage2_5[31]},
      {stage3_6[21],stage3_5[24],stage3_4[30],stage3_3[30]}
   );
   gpc207_4 gpc8598 (
      {stage2_3[125], stage2_3[126], stage2_3[127], stage2_3[128], stage2_3[129], stage2_3[130], stage2_3[131]},
      {stage2_5[32], stage2_5[33]},
      {stage3_6[22],stage3_5[25],stage3_4[31],stage3_3[31]}
   );
   gpc207_4 gpc8599 (
      {stage2_3[132], stage2_3[133], stage2_3[134], stage2_3[135], stage2_3[136], stage2_3[137], stage2_3[138]},
      {stage2_5[34], stage2_5[35]},
      {stage3_6[23],stage3_5[26],stage3_4[32],stage3_3[32]}
   );
   gpc207_4 gpc8600 (
      {stage2_3[139], stage2_3[140], stage2_3[141], stage2_3[142], stage2_3[143], stage2_3[144], stage2_3[145]},
      {stage2_5[36], stage2_5[37]},
      {stage3_6[24],stage3_5[27],stage3_4[33],stage3_3[33]}
   );
   gpc207_4 gpc8601 (
      {stage2_3[146], stage2_3[147], stage2_3[148], stage2_3[149], stage2_3[150], stage2_3[151], stage2_3[152]},
      {stage2_5[38], stage2_5[39]},
      {stage3_6[25],stage3_5[28],stage3_4[34],stage3_3[34]}
   );
   gpc207_4 gpc8602 (
      {stage2_3[153], stage2_3[154], stage2_3[155], stage2_3[156], stage2_3[157], stage2_3[158], stage2_3[159]},
      {stage2_5[40], stage2_5[41]},
      {stage3_6[26],stage3_5[29],stage3_4[35],stage3_3[35]}
   );
   gpc207_4 gpc8603 (
      {stage2_3[160], stage2_3[161], stage2_3[162], stage2_3[163], stage2_3[164], stage2_3[165], stage2_3[166]},
      {stage2_5[42], stage2_5[43]},
      {stage3_6[27],stage3_5[30],stage3_4[36],stage3_3[36]}
   );
   gpc207_4 gpc8604 (
      {stage2_3[167], stage2_3[168], stage2_3[169], stage2_3[170], stage2_3[171], stage2_3[172], stage2_3[173]},
      {stage2_5[44], stage2_5[45]},
      {stage3_6[28],stage3_5[31],stage3_4[37],stage3_3[37]}
   );
   gpc207_4 gpc8605 (
      {stage2_3[174], stage2_3[175], stage2_3[176], stage2_3[177], stage2_3[178], stage2_3[179], stage2_3[180]},
      {stage2_5[46], stage2_5[47]},
      {stage3_6[29],stage3_5[32],stage3_4[38],stage3_3[38]}
   );
   gpc207_4 gpc8606 (
      {stage2_3[181], stage2_3[182], stage2_3[183], stage2_3[184], stage2_3[185], stage2_3[186], stage2_3[187]},
      {stage2_5[48], stage2_5[49]},
      {stage3_6[30],stage3_5[33],stage3_4[39],stage3_3[39]}
   );
   gpc207_4 gpc8607 (
      {stage2_3[188], stage2_3[189], stage2_3[190], stage2_3[191], stage2_3[192], stage2_3[193], stage2_3[194]},
      {stage2_5[50], stage2_5[51]},
      {stage3_6[31],stage3_5[34],stage3_4[40],stage3_3[40]}
   );
   gpc207_4 gpc8608 (
      {stage2_3[195], stage2_3[196], stage2_3[197], stage2_3[198], stage2_3[199], stage2_3[200], stage2_3[201]},
      {stage2_5[52], stage2_5[53]},
      {stage3_6[32],stage3_5[35],stage3_4[41],stage3_3[41]}
   );
   gpc207_4 gpc8609 (
      {stage2_3[202], stage2_3[203], stage2_3[204], stage2_3[205], stage2_3[206], stage2_3[207], stage2_3[208]},
      {stage2_5[54], stage2_5[55]},
      {stage3_6[33],stage3_5[36],stage3_4[42],stage3_3[42]}
   );
   gpc207_4 gpc8610 (
      {stage2_3[209], stage2_3[210], stage2_3[211], stage2_3[212], stage2_3[213], stage2_3[214], stage2_3[215]},
      {stage2_5[56], stage2_5[57]},
      {stage3_6[34],stage3_5[37],stage3_4[43],stage3_3[43]}
   );
   gpc615_5 gpc8611 (
      {stage2_3[216], stage2_3[217], stage2_3[218], stage2_3[219], stage2_3[220]},
      {stage2_4[38]},
      {stage2_5[58], stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63]},
      {stage3_7[0],stage3_6[35],stage3_5[38],stage3_4[44],stage3_3[44]}
   );
   gpc615_5 gpc8612 (
      {stage2_3[221], stage2_3[222], stage2_3[223], stage2_3[224], stage2_3[225]},
      {stage2_4[39]},
      {stage2_5[64], stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage3_7[1],stage3_6[36],stage3_5[39],stage3_4[45],stage3_3[45]}
   );
   gpc615_5 gpc8613 (
      {stage2_3[226], stage2_3[227], stage2_3[228], stage2_3[229], stage2_3[230]},
      {stage2_4[40]},
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75]},
      {stage3_7[2],stage3_6[37],stage3_5[40],stage3_4[46],stage3_3[46]}
   );
   gpc615_5 gpc8614 (
      {stage2_3[231], stage2_3[232], stage2_3[233], stage2_3[234], stage2_3[235]},
      {stage2_4[41]},
      {stage2_5[76], stage2_5[77], stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81]},
      {stage3_7[3],stage3_6[38],stage3_5[41],stage3_4[47],stage3_3[47]}
   );
   gpc615_5 gpc8615 (
      {stage2_3[236], stage2_3[237], stage2_3[238], stage2_3[239], stage2_3[240]},
      {stage2_4[42]},
      {stage2_5[82], stage2_5[83], stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87]},
      {stage3_7[4],stage3_6[39],stage3_5[42],stage3_4[48],stage3_3[48]}
   );
   gpc615_5 gpc8616 (
      {stage2_3[241], stage2_3[242], stage2_3[243], stage2_3[244], stage2_3[245]},
      {stage2_4[43]},
      {stage2_5[88], stage2_5[89], stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93]},
      {stage3_7[5],stage3_6[40],stage3_5[43],stage3_4[49],stage3_3[49]}
   );
   gpc615_5 gpc8617 (
      {stage2_3[246], stage2_3[247], stage2_3[248], stage2_3[249], stage2_3[250]},
      {stage2_4[44]},
      {stage2_5[94], stage2_5[95], stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99]},
      {stage3_7[6],stage3_6[41],stage3_5[44],stage3_4[50],stage3_3[50]}
   );
   gpc615_5 gpc8618 (
      {stage2_3[251], stage2_3[252], stage2_3[253], 1'b0, 1'b0},
      {stage2_4[45]},
      {stage2_5[100], stage2_5[101], stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105]},
      {stage3_7[7],stage3_6[42],stage3_5[45],stage3_4[51],stage3_3[51]}
   );
   gpc606_5 gpc8619 (
      {stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[43],stage3_5[46],stage3_4[52]}
   );
   gpc606_5 gpc8620 (
      {stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[44],stage3_5[47],stage3_4[53]}
   );
   gpc606_5 gpc8621 (
      {stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[45],stage3_5[48],stage3_4[54]}
   );
   gpc606_5 gpc8622 (
      {stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[46],stage3_5[49],stage3_4[55]}
   );
   gpc606_5 gpc8623 (
      {stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[47],stage3_5[50],stage3_4[56]}
   );
   gpc606_5 gpc8624 (
      {stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[48],stage3_5[51],stage3_4[57]}
   );
   gpc606_5 gpc8625 (
      {stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[14],stage3_6[49],stage3_5[52],stage3_4[58]}
   );
   gpc606_5 gpc8626 (
      {stage2_4[88], stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], 1'b0},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[15],stage3_6[50],stage3_5[53],stage3_4[59]}
   );
   gpc606_5 gpc8627 (
      {stage2_5[106], stage2_5[107], stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[16],stage3_6[51],stage3_5[54]}
   );
   gpc615_5 gpc8628 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[9],stage3_7[17],stage3_6[52]}
   );
   gpc615_5 gpc8629 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[7]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[10],stage3_7[18],stage3_6[53]}
   );
   gpc615_5 gpc8630 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[8]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[11],stage3_7[19],stage3_6[54]}
   );
   gpc615_5 gpc8631 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[9]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[4],stage3_8[12],stage3_7[20],stage3_6[55]}
   );
   gpc615_5 gpc8632 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[10]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[5],stage3_8[13],stage3_7[21],stage3_6[56]}
   );
   gpc615_5 gpc8633 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[11]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[6],stage3_8[14],stage3_7[22],stage3_6[57]}
   );
   gpc615_5 gpc8634 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[12]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[7],stage3_8[15],stage3_7[23],stage3_6[58]}
   );
   gpc615_5 gpc8635 (
      {stage2_6[83], stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87]},
      {stage2_7[13]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[8],stage3_8[16],stage3_7[24],stage3_6[59]}
   );
   gpc615_5 gpc8636 (
      {stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91], stage2_6[92]},
      {stage2_7[14]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[9],stage3_8[17],stage3_7[25],stage3_6[60]}
   );
   gpc615_5 gpc8637 (
      {stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_7[15]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[10],stage3_8[18],stage3_7[26],stage3_6[61]}
   );
   gpc615_5 gpc8638 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102]},
      {stage2_7[16]},
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage3_10[10],stage3_9[11],stage3_8[19],stage3_7[27],stage3_6[62]}
   );
   gpc615_5 gpc8639 (
      {stage2_6[103], stage2_6[104], stage2_6[105], stage2_6[106], stage2_6[107]},
      {stage2_7[17]},
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage3_10[11],stage3_9[12],stage3_8[20],stage3_7[28],stage3_6[63]}
   );
   gpc615_5 gpc8640 (
      {stage2_6[108], stage2_6[109], stage2_6[110], stage2_6[111], stage2_6[112]},
      {stage2_7[18]},
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage3_10[12],stage3_9[13],stage3_8[21],stage3_7[29],stage3_6[64]}
   );
   gpc615_5 gpc8641 (
      {stage2_6[113], stage2_6[114], stage2_6[115], stage2_6[116], stage2_6[117]},
      {stage2_7[19]},
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage3_10[13],stage3_9[14],stage3_8[22],stage3_7[30],stage3_6[65]}
   );
   gpc615_5 gpc8642 (
      {stage2_6[118], stage2_6[119], stage2_6[120], 1'b0, 1'b0},
      {stage2_7[20]},
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage3_10[14],stage3_9[15],stage3_8[23],stage3_7[31],stage3_6[66]}
   );
   gpc2116_5 gpc8643 (
      {stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[90]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[15],stage3_9[16],stage3_8[24],stage3_7[32]}
   );
   gpc2116_5 gpc8644 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[91]},
      {stage2_9[1]},
      {stage2_10[2], stage2_10[3]},
      {stage3_11[1],stage3_10[16],stage3_9[17],stage3_8[25],stage3_7[33]}
   );
   gpc2116_5 gpc8645 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[92]},
      {stage2_9[2]},
      {stage2_10[4], stage2_10[5]},
      {stage3_11[2],stage3_10[17],stage3_9[18],stage3_8[26],stage3_7[34]}
   );
   gpc2116_5 gpc8646 (
      {stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44]},
      {stage2_8[93]},
      {stage2_9[3]},
      {stage2_10[6], stage2_10[7]},
      {stage3_11[3],stage3_10[18],stage3_9[19],stage3_8[27],stage3_7[35]}
   );
   gpc2116_5 gpc8647 (
      {stage2_7[45], stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[94]},
      {stage2_9[4]},
      {stage2_10[8], stage2_10[9]},
      {stage3_11[4],stage3_10[19],stage3_9[20],stage3_8[28],stage3_7[36]}
   );
   gpc2116_5 gpc8648 (
      {stage2_7[51], stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[95]},
      {stage2_9[5]},
      {stage2_10[10], stage2_10[11]},
      {stage3_11[5],stage3_10[20],stage3_9[21],stage3_8[29],stage3_7[37]}
   );
   gpc2116_5 gpc8649 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62]},
      {stage2_8[96]},
      {stage2_9[6]},
      {stage2_10[12], stage2_10[13]},
      {stage3_11[6],stage3_10[21],stage3_9[22],stage3_8[30],stage3_7[38]}
   );
   gpc2116_5 gpc8650 (
      {stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[97]},
      {stage2_9[7]},
      {stage2_10[14], stage2_10[15]},
      {stage3_11[7],stage3_10[22],stage3_9[23],stage3_8[31],stage3_7[39]}
   );
   gpc2116_5 gpc8651 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73], stage2_7[74]},
      {stage2_8[98]},
      {stage2_9[8]},
      {stage2_10[16], stage2_10[17]},
      {stage3_11[8],stage3_10[23],stage3_9[24],stage3_8[32],stage3_7[40]}
   );
   gpc615_5 gpc8652 (
      {stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78], stage2_7[79]},
      {stage2_8[99]},
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage3_11[9],stage3_10[24],stage3_9[25],stage3_8[33],stage3_7[41]}
   );
   gpc615_5 gpc8653 (
      {stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83], stage2_7[84]},
      {stage2_8[100]},
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage3_11[10],stage3_10[25],stage3_9[26],stage3_8[34],stage3_7[42]}
   );
   gpc606_5 gpc8654 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[0],stage3_11[11],stage3_10[26],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc8655 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[1],stage3_11[12],stage3_10[27],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc8656 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[2],stage3_11[13],stage3_10[28],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc8657 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[3],stage3_11[14],stage3_10[29],stage3_9[30],stage3_8[38]}
   );
   gpc606_5 gpc8658 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[4],stage3_11[15],stage3_10[30],stage3_9[31],stage3_8[39]}
   );
   gpc606_5 gpc8659 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[5],stage3_11[16],stage3_10[31],stage3_9[32],stage3_8[40]}
   );
   gpc606_5 gpc8660 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[6],stage3_11[17],stage3_10[32],stage3_9[33],stage3_8[41]}
   );
   gpc606_5 gpc8661 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[7],stage3_11[18],stage3_10[33],stage3_9[34],stage3_8[42]}
   );
   gpc606_5 gpc8662 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[8],stage3_11[19],stage3_10[34],stage3_9[35],stage3_8[43]}
   );
   gpc606_5 gpc8663 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], stage2_8[160]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[9],stage3_11[20],stage3_10[35],stage3_9[36],stage3_8[44]}
   );
   gpc606_5 gpc8664 (
      {stage2_8[161], stage2_8[162], stage2_8[163], stage2_8[164], stage2_8[165], stage2_8[166]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[10],stage3_11[21],stage3_10[36],stage3_9[37],stage3_8[45]}
   );
   gpc606_5 gpc8665 (
      {stage2_8[167], stage2_8[168], stage2_8[169], stage2_8[170], stage2_8[171], stage2_8[172]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[11],stage3_11[22],stage3_10[37],stage3_9[38],stage3_8[46]}
   );
   gpc606_5 gpc8666 (
      {stage2_9[21], stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[12],stage3_11[23],stage3_10[38],stage3_9[39]}
   );
   gpc606_5 gpc8667 (
      {stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30], stage2_9[31], stage2_9[32]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[13],stage3_11[24],stage3_10[39],stage3_9[40]}
   );
   gpc606_5 gpc8668 (
      {stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37], stage2_9[38]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[14],stage3_11[25],stage3_10[40],stage3_9[41]}
   );
   gpc606_5 gpc8669 (
      {stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43], stage2_9[44]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[15],stage3_11[26],stage3_10[41],stage3_9[42]}
   );
   gpc606_5 gpc8670 (
      {stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49], stage2_9[50]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[16],stage3_11[27],stage3_10[42],stage3_9[43]}
   );
   gpc606_5 gpc8671 (
      {stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[17],stage3_11[28],stage3_10[43],stage3_9[44]}
   );
   gpc606_5 gpc8672 (
      {stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[18],stage3_11[29],stage3_10[44],stage3_9[45]}
   );
   gpc606_5 gpc8673 (
      {stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67], stage2_9[68]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[19],stage3_11[30],stage3_10[45],stage3_9[46]}
   );
   gpc606_5 gpc8674 (
      {stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[20],stage3_11[31],stage3_10[46],stage3_9[47]}
   );
   gpc606_5 gpc8675 (
      {stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[21],stage3_11[32],stage3_10[47],stage3_9[48]}
   );
   gpc606_5 gpc8676 (
      {stage2_9[81], stage2_9[82], stage2_9[83], stage2_9[84], stage2_9[85], stage2_9[86]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[22],stage3_11[33],stage3_10[48],stage3_9[49]}
   );
   gpc606_5 gpc8677 (
      {stage2_9[87], stage2_9[88], stage2_9[89], stage2_9[90], stage2_9[91], stage2_9[92]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[23],stage3_11[34],stage3_10[49],stage3_9[50]}
   );
   gpc606_5 gpc8678 (
      {stage2_9[93], stage2_9[94], stage2_9[95], stage2_9[96], stage2_9[97], stage2_9[98]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[24],stage3_11[35],stage3_10[50],stage3_9[51]}
   );
   gpc606_5 gpc8679 (
      {stage2_9[99], stage2_9[100], stage2_9[101], stage2_9[102], stage2_9[103], stage2_9[104]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[25],stage3_11[36],stage3_10[51],stage3_9[52]}
   );
   gpc215_4 gpc8680 (
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94]},
      {stage2_11[84]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[14],stage3_12[26],stage3_11[37],stage3_10[52]}
   );
   gpc215_4 gpc8681 (
      {stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99]},
      {stage2_11[85]},
      {stage2_12[2], stage2_12[3]},
      {stage3_13[15],stage3_12[27],stage3_11[38],stage3_10[53]}
   );
   gpc215_4 gpc8682 (
      {stage2_10[100], stage2_10[101], stage2_10[102], stage2_10[103], stage2_10[104]},
      {stage2_11[86]},
      {stage2_12[4], stage2_12[5]},
      {stage3_13[16],stage3_12[28],stage3_11[39],stage3_10[54]}
   );
   gpc615_5 gpc8683 (
      {stage2_10[105], stage2_10[106], stage2_10[107], stage2_10[108], stage2_10[109]},
      {stage2_11[87]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[0],stage3_13[17],stage3_12[29],stage3_11[40],stage3_10[55]}
   );
   gpc615_5 gpc8684 (
      {stage2_10[110], stage2_10[111], stage2_10[112], stage2_10[113], stage2_10[114]},
      {stage2_11[88]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[1],stage3_13[18],stage3_12[30],stage3_11[41],stage3_10[56]}
   );
   gpc615_5 gpc8685 (
      {stage2_10[115], stage2_10[116], stage2_10[117], stage2_10[118], stage2_10[119]},
      {stage2_11[89]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[2],stage3_13[19],stage3_12[31],stage3_11[42],stage3_10[57]}
   );
   gpc615_5 gpc8686 (
      {stage2_10[120], stage2_10[121], stage2_10[122], stage2_10[123], stage2_10[124]},
      {stage2_11[90]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[3],stage3_13[20],stage3_12[32],stage3_11[43],stage3_10[58]}
   );
   gpc606_5 gpc8687 (
      {stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[4],stage3_13[21],stage3_12[33],stage3_11[44]}
   );
   gpc606_5 gpc8688 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[5],stage3_13[22],stage3_12[34],stage3_11[45]}
   );
   gpc606_5 gpc8689 (
      {stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[6],stage3_13[23],stage3_12[35],stage3_11[46]}
   );
   gpc606_5 gpc8690 (
      {stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[7],stage3_13[24],stage3_12[36],stage3_11[47]}
   );
   gpc615_5 gpc8691 (
      {stage2_11[115], stage2_11[116], stage2_11[117], stage2_11[118], stage2_11[119]},
      {stage2_12[30]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[8],stage3_13[25],stage3_12[37],stage3_11[48]}
   );
   gpc615_5 gpc8692 (
      {stage2_11[120], stage2_11[121], stage2_11[122], stage2_11[123], stage2_11[124]},
      {stage2_12[31]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[9],stage3_13[26],stage3_12[38],stage3_11[49]}
   );
   gpc606_5 gpc8693 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[6],stage3_14[10],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc8694 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[7],stage3_14[11],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc8695 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[8],stage3_14[12],stage3_13[29],stage3_12[41]}
   );
   gpc606_5 gpc8696 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[9],stage3_14[13],stage3_13[30],stage3_12[42]}
   );
   gpc606_5 gpc8697 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[10],stage3_14[14],stage3_13[31],stage3_12[43]}
   );
   gpc606_5 gpc8698 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[11],stage3_14[15],stage3_13[32],stage3_12[44]}
   );
   gpc606_5 gpc8699 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[12],stage3_14[16],stage3_13[33],stage3_12[45]}
   );
   gpc606_5 gpc8700 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[13],stage3_14[17],stage3_13[34],stage3_12[46]}
   );
   gpc606_5 gpc8701 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[14],stage3_14[18],stage3_13[35],stage3_12[47]}
   );
   gpc606_5 gpc8702 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[15],stage3_14[19],stage3_13[36],stage3_12[48]}
   );
   gpc623_5 gpc8703 (
      {stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_13[36], stage2_13[37]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[16],stage3_14[20],stage3_13[37],stage3_12[49]}
   );
   gpc623_5 gpc8704 (
      {stage2_12[95], stage2_12[96], stage2_12[97]},
      {stage2_13[38], stage2_13[39]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[17],stage3_14[21],stage3_13[38],stage3_12[50]}
   );
   gpc615_5 gpc8705 (
      {stage2_13[40], stage2_13[41], stage2_13[42], stage2_13[43], stage2_13[44]},
      {stage2_14[72]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[18],stage3_14[22],stage3_13[39]}
   );
   gpc615_5 gpc8706 (
      {stage2_13[45], stage2_13[46], stage2_13[47], stage2_13[48], stage2_13[49]},
      {stage2_14[73]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[19],stage3_14[23],stage3_13[40]}
   );
   gpc615_5 gpc8707 (
      {stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53], stage2_13[54]},
      {stage2_14[74]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[20],stage3_14[24],stage3_13[41]}
   );
   gpc615_5 gpc8708 (
      {stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_14[75]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[21],stage3_14[25],stage3_13[42]}
   );
   gpc615_5 gpc8709 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64]},
      {stage2_14[76]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[22],stage3_14[26],stage3_13[43]}
   );
   gpc615_5 gpc8710 (
      {stage2_13[65], stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69]},
      {stage2_14[77]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[23],stage3_14[27],stage3_13[44]}
   );
   gpc606_5 gpc8711 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[18],stage3_15[24],stage3_14[28]}
   );
   gpc606_5 gpc8712 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[19],stage3_15[25],stage3_14[29]}
   );
   gpc615_5 gpc8713 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94]},
      {stage2_15[36]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[20],stage3_15[26],stage3_14[30]}
   );
   gpc615_5 gpc8714 (
      {stage2_14[95], stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99]},
      {stage2_15[37]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[21],stage3_15[27],stage3_14[31]}
   );
   gpc615_5 gpc8715 (
      {stage2_14[100], stage2_14[101], stage2_14[102], stage2_14[103], stage2_14[104]},
      {stage2_15[38]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[22],stage3_15[28],stage3_14[32]}
   );
   gpc615_5 gpc8716 (
      {stage2_14[105], stage2_14[106], stage2_14[107], stage2_14[108], stage2_14[109]},
      {stage2_15[39]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[23],stage3_15[29],stage3_14[33]}
   );
   gpc615_5 gpc8717 (
      {stage2_14[110], stage2_14[111], stage2_14[112], stage2_14[113], stage2_14[114]},
      {stage2_15[40]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[24],stage3_15[30],stage3_14[34]}
   );
   gpc207_4 gpc8718 (
      {stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[7],stage3_17[13],stage3_16[25],stage3_15[31]}
   );
   gpc615_5 gpc8719 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[42]},
      {stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7]},
      {stage3_19[0],stage3_18[8],stage3_17[14],stage3_16[26],stage3_15[32]}
   );
   gpc615_5 gpc8720 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[43]},
      {stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13]},
      {stage3_19[1],stage3_18[9],stage3_17[15],stage3_16[27],stage3_15[33]}
   );
   gpc615_5 gpc8721 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[44]},
      {stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19]},
      {stage3_19[2],stage3_18[10],stage3_17[16],stage3_16[28],stage3_15[34]}
   );
   gpc615_5 gpc8722 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[45]},
      {stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25]},
      {stage3_19[3],stage3_18[11],stage3_17[17],stage3_16[29],stage3_15[35]}
   );
   gpc615_5 gpc8723 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[46]},
      {stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31]},
      {stage3_19[4],stage3_18[12],stage3_17[18],stage3_16[30],stage3_15[36]}
   );
   gpc615_5 gpc8724 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[47]},
      {stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37]},
      {stage3_19[5],stage3_18[13],stage3_17[19],stage3_16[31],stage3_15[37]}
   );
   gpc615_5 gpc8725 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[48]},
      {stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43]},
      {stage3_19[6],stage3_18[14],stage3_17[20],stage3_16[32],stage3_15[38]}
   );
   gpc615_5 gpc8726 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[49]},
      {stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49]},
      {stage3_19[7],stage3_18[15],stage3_17[21],stage3_16[33],stage3_15[39]}
   );
   gpc615_5 gpc8727 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[50]},
      {stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55]},
      {stage3_19[8],stage3_18[16],stage3_17[22],stage3_16[34],stage3_15[40]}
   );
   gpc615_5 gpc8728 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[51]},
      {stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61]},
      {stage3_19[9],stage3_18[17],stage3_17[23],stage3_16[35],stage3_15[41]}
   );
   gpc615_5 gpc8729 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[52]},
      {stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67]},
      {stage3_19[10],stage3_18[18],stage3_17[24],stage3_16[36],stage3_15[42]}
   );
   gpc615_5 gpc8730 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[53]},
      {stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73]},
      {stage3_19[11],stage3_18[19],stage3_17[25],stage3_16[37],stage3_15[43]}
   );
   gpc606_5 gpc8731 (
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[12],stage3_18[20],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc8732 (
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[13],stage3_18[21],stage3_17[27],stage3_16[39]}
   );
   gpc606_5 gpc8733 (
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[14],stage3_18[22],stage3_17[28],stage3_16[40]}
   );
   gpc606_5 gpc8734 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[15],stage3_18[23],stage3_17[29],stage3_16[41]}
   );
   gpc606_5 gpc8735 (
      {stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[16],stage3_18[24],stage3_17[30],stage3_16[42]}
   );
   gpc606_5 gpc8736 (
      {stage2_16[84], stage2_16[85], stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89]},
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage3_20[5],stage3_19[17],stage3_18[25],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc8737 (
      {stage2_16[90], stage2_16[91], stage2_16[92], stage2_16[93], stage2_16[94], stage2_16[95]},
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41]},
      {stage3_20[6],stage3_19[18],stage3_18[26],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc8738 (
      {stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[7],stage3_19[19],stage3_18[27],stage3_17[33]}
   );
   gpc2135_5 gpc8739 (
      {stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[1],stage3_20[8],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc8740 (
      {stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50], stage2_18[51]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[2],stage3_20[9],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc8741 (
      {stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55], stage2_18[56]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[3],stage3_20[10],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc8742 (
      {stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60], stage2_18[61]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[4],stage3_20[11],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc8743 (
      {stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[5],stage3_20[12],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc8744 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[6],stage3_20[13],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc8745 (
      {stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75], stage2_18[76]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[7],stage3_20[14],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc8746 (
      {stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80], stage2_18[81]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[8],stage3_20[15],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc8747 (
      {stage2_18[82], stage2_18[83], stage2_18[84], stage2_18[85], stage2_18[86]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[9],stage3_20[16],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc8748 (
      {stage2_18[87], stage2_18[88], stage2_18[89], stage2_18[90], stage2_18[91]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[10],stage3_20[17],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc8749 (
      {stage2_18[92], stage2_18[93], stage2_18[94], stage2_18[95], stage2_18[96]},
      {stage2_19[36], stage2_19[37], stage2_19[38]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[11],stage3_20[18],stage3_19[30],stage3_18[38]}
   );
   gpc2135_5 gpc8750 (
      {stage2_18[97], stage2_18[98], stage2_18[99], stage2_18[100], stage2_18[101]},
      {stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[12],stage3_20[19],stage3_19[31],stage3_18[39]}
   );
   gpc2135_5 gpc8751 (
      {stage2_18[102], stage2_18[103], stage2_18[104], stage2_18[105], stage2_18[106]},
      {stage2_19[42], stage2_19[43], stage2_19[44]},
      {stage2_20[12]},
      {stage2_21[24], stage2_21[25]},
      {stage3_22[12],stage3_21[13],stage3_20[20],stage3_19[32],stage3_18[40]}
   );
   gpc2135_5 gpc8752 (
      {stage2_18[107], stage2_18[108], stage2_18[109], stage2_18[110], stage2_18[111]},
      {stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[13]},
      {stage2_21[26], stage2_21[27]},
      {stage3_22[13],stage3_21[14],stage3_20[21],stage3_19[33],stage3_18[41]}
   );
   gpc2135_5 gpc8753 (
      {stage2_18[112], stage2_18[113], stage2_18[114], stage2_18[115], stage2_18[116]},
      {stage2_19[48], stage2_19[49], stage2_19[50]},
      {stage2_20[14]},
      {stage2_21[28], stage2_21[29]},
      {stage3_22[14],stage3_21[15],stage3_20[22],stage3_19[34],stage3_18[42]}
   );
   gpc2135_5 gpc8754 (
      {stage2_18[117], stage2_18[118], stage2_18[119], stage2_18[120], stage2_18[121]},
      {stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_20[15]},
      {stage2_21[30], stage2_21[31]},
      {stage3_22[15],stage3_21[16],stage3_20[23],stage3_19[35],stage3_18[43]}
   );
   gpc2135_5 gpc8755 (
      {stage2_18[122], stage2_18[123], stage2_18[124], stage2_18[125], stage2_18[126]},
      {stage2_19[54], stage2_19[55], stage2_19[56]},
      {stage2_20[16]},
      {stage2_21[32], stage2_21[33]},
      {stage3_22[16],stage3_21[17],stage3_20[24],stage3_19[36],stage3_18[44]}
   );
   gpc2135_5 gpc8756 (
      {stage2_18[127], stage2_18[128], stage2_18[129], stage2_18[130], stage2_18[131]},
      {stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage2_20[17]},
      {stage2_21[34], stage2_21[35]},
      {stage3_22[17],stage3_21[18],stage3_20[25],stage3_19[37],stage3_18[45]}
   );
   gpc2135_5 gpc8757 (
      {stage2_18[132], stage2_18[133], stage2_18[134], stage2_18[135], stage2_18[136]},
      {stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[18]},
      {stage2_21[36], stage2_21[37]},
      {stage3_22[18],stage3_21[19],stage3_20[26],stage3_19[38],stage3_18[46]}
   );
   gpc2135_5 gpc8758 (
      {stage2_18[137], stage2_18[138], stage2_18[139], stage2_18[140], stage2_18[141]},
      {stage2_19[63], stage2_19[64], stage2_19[65]},
      {stage2_20[19]},
      {stage2_21[38], stage2_21[39]},
      {stage3_22[19],stage3_21[20],stage3_20[27],stage3_19[39],stage3_18[47]}
   );
   gpc2135_5 gpc8759 (
      {stage2_18[142], stage2_18[143], stage2_18[144], stage2_18[145], stage2_18[146]},
      {stage2_19[66], stage2_19[67], stage2_19[68]},
      {stage2_20[20]},
      {stage2_21[40], stage2_21[41]},
      {stage3_22[20],stage3_21[21],stage3_20[28],stage3_19[40],stage3_18[48]}
   );
   gpc615_5 gpc8760 (
      {stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72], stage2_19[73]},
      {stage2_20[21]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[0],stage3_22[21],stage3_21[22],stage3_20[29],stage3_19[41]}
   );
   gpc615_5 gpc8761 (
      {stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77], stage2_19[78]},
      {stage2_20[22]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[1],stage3_22[22],stage3_21[23],stage3_20[30],stage3_19[42]}
   );
   gpc615_5 gpc8762 (
      {stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82], stage2_19[83]},
      {stage2_20[23]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[2],stage3_22[23],stage3_21[24],stage3_20[31],stage3_19[43]}
   );
   gpc615_5 gpc8763 (
      {stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87], stage2_19[88]},
      {stage2_20[24]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[3],stage3_22[24],stage3_21[25],stage3_20[32],stage3_19[44]}
   );
   gpc615_5 gpc8764 (
      {stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92], stage2_19[93]},
      {stage2_20[25]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[4],stage3_22[25],stage3_21[26],stage3_20[33],stage3_19[45]}
   );
   gpc606_5 gpc8765 (
      {stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30], stage2_20[31]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[26],stage3_21[27],stage3_20[34]}
   );
   gpc606_5 gpc8766 (
      {stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35], stage2_20[36], stage2_20[37]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[27],stage3_21[28],stage3_20[35]}
   );
   gpc606_5 gpc8767 (
      {stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[28],stage3_21[29],stage3_20[36]}
   );
   gpc606_5 gpc8768 (
      {stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47], stage2_20[48], stage2_20[49]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[8],stage3_22[29],stage3_21[30],stage3_20[37]}
   );
   gpc606_5 gpc8769 (
      {stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53], stage2_20[54], stage2_20[55]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[9],stage3_22[30],stage3_21[31],stage3_20[38]}
   );
   gpc606_5 gpc8770 (
      {stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59], stage2_20[60], stage2_20[61]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[10],stage3_22[31],stage3_21[32],stage3_20[39]}
   );
   gpc615_5 gpc8771 (
      {stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65], stage2_20[66]},
      {stage2_21[72]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[11],stage3_22[32],stage3_21[33],stage3_20[40]}
   );
   gpc615_5 gpc8772 (
      {stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage2_21[73]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage3_24[7],stage3_23[12],stage3_22[33],stage3_21[34],stage3_20[41]}
   );
   gpc606_5 gpc8773 (
      {stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77], stage2_21[78], stage2_21[79]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[8],stage3_23[13],stage3_22[34],stage3_21[35]}
   );
   gpc606_5 gpc8774 (
      {stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83], stage2_21[84], stage2_21[85]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[9],stage3_23[14],stage3_22[35],stage3_21[36]}
   );
   gpc615_5 gpc8775 (
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[10],stage3_23[15],stage3_22[36]}
   );
   gpc615_5 gpc8776 (
      {stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[11],stage3_23[16],stage3_22[37]}
   );
   gpc615_5 gpc8777 (
      {stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61], stage2_22[62]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[12],stage3_23[17],stage3_22[38]}
   );
   gpc615_5 gpc8778 (
      {stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66], stage2_22[67]},
      {stage2_23[15]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[5],stage3_24[13],stage3_23[18],stage3_22[39]}
   );
   gpc615_5 gpc8779 (
      {stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71], stage2_22[72]},
      {stage2_23[16]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[6],stage3_24[14],stage3_23[19],stage3_22[40]}
   );
   gpc615_5 gpc8780 (
      {stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76], stage2_22[77]},
      {stage2_23[17]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[7],stage3_24[15],stage3_23[20],stage3_22[41]}
   );
   gpc615_5 gpc8781 (
      {stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81], stage2_22[82]},
      {stage2_23[18]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[8],stage3_24[16],stage3_23[21],stage3_22[42]}
   );
   gpc615_5 gpc8782 (
      {stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86], stage2_22[87]},
      {stage2_23[19]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[9],stage3_24[17],stage3_23[22],stage3_22[43]}
   );
   gpc615_5 gpc8783 (
      {stage2_22[88], stage2_22[89], stage2_22[90], stage2_22[91], stage2_22[92]},
      {stage2_23[20]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[10],stage3_24[18],stage3_23[23],stage3_22[44]}
   );
   gpc615_5 gpc8784 (
      {stage2_22[93], stage2_22[94], stage2_22[95], stage2_22[96], stage2_22[97]},
      {stage2_23[21]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[11],stage3_24[19],stage3_23[24],stage3_22[45]}
   );
   gpc615_5 gpc8785 (
      {stage2_22[98], stage2_22[99], stage2_22[100], stage2_22[101], stage2_22[102]},
      {stage2_23[22]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[12],stage3_24[20],stage3_23[25],stage3_22[46]}
   );
   gpc615_5 gpc8786 (
      {stage2_22[103], stage2_22[104], stage2_22[105], stage2_22[106], stage2_22[107]},
      {stage2_23[23]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[13],stage3_24[21],stage3_23[26],stage3_22[47]}
   );
   gpc615_5 gpc8787 (
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28]},
      {stage2_24[72]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[12],stage3_25[14],stage3_24[22],stage3_23[27]}
   );
   gpc615_5 gpc8788 (
      {stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33]},
      {stage2_24[73]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[13],stage3_25[15],stage3_24[23],stage3_23[28]}
   );
   gpc615_5 gpc8789 (
      {stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage2_24[74]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[14],stage3_25[16],stage3_24[24],stage3_23[29]}
   );
   gpc615_5 gpc8790 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43]},
      {stage2_24[75]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[15],stage3_25[17],stage3_24[25],stage3_23[30]}
   );
   gpc615_5 gpc8791 (
      {stage2_23[44], stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48]},
      {stage2_24[76]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[16],stage3_25[18],stage3_24[26],stage3_23[31]}
   );
   gpc615_5 gpc8792 (
      {stage2_23[49], stage2_23[50], stage2_23[51], stage2_23[52], stage2_23[53]},
      {stage2_24[77]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[17],stage3_25[19],stage3_24[27],stage3_23[32]}
   );
   gpc615_5 gpc8793 (
      {stage2_23[54], stage2_23[55], stage2_23[56], stage2_23[57], stage2_23[58]},
      {stage2_24[78]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[18],stage3_25[20],stage3_24[28],stage3_23[33]}
   );
   gpc615_5 gpc8794 (
      {stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62], stage2_23[63]},
      {stage2_24[79]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[19],stage3_25[21],stage3_24[29],stage3_23[34]}
   );
   gpc615_5 gpc8795 (
      {stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_24[80]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[20],stage3_25[22],stage3_24[30],stage3_23[35]}
   );
   gpc615_5 gpc8796 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73]},
      {stage2_24[81]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[21],stage3_25[23],stage3_24[31],stage3_23[36]}
   );
   gpc615_5 gpc8797 (
      {stage2_23[74], stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78]},
      {stage2_24[82]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[22],stage3_25[24],stage3_24[32],stage3_23[37]}
   );
   gpc615_5 gpc8798 (
      {stage2_23[79], stage2_23[80], stage2_23[81], stage2_23[82], stage2_23[83]},
      {stage2_24[83]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[23],stage3_25[25],stage3_24[33],stage3_23[38]}
   );
   gpc615_5 gpc8799 (
      {stage2_23[84], stage2_23[85], stage2_23[86], stage2_23[87], stage2_23[88]},
      {stage2_24[84]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[24],stage3_25[26],stage3_24[34],stage3_23[39]}
   );
   gpc606_5 gpc8800 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[13],stage3_26[25],stage3_25[27]}
   );
   gpc606_5 gpc8801 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[1],stage3_27[14],stage3_26[26],stage3_25[28]}
   );
   gpc606_5 gpc8802 (
      {stage2_25[90], stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[2],stage3_27[15],stage3_26[27],stage3_25[29]}
   );
   gpc606_5 gpc8803 (
      {stage2_25[96], stage2_25[97], stage2_25[98], stage2_25[99], stage2_25[100], stage2_25[101]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[3],stage3_27[16],stage3_26[28],stage3_25[30]}
   );
   gpc117_4 gpc8804 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6]},
      {stage2_27[24]},
      {stage2_28[0]},
      {stage3_29[4],stage3_28[4],stage3_27[17],stage3_26[29]}
   );
   gpc117_4 gpc8805 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12], stage2_26[13]},
      {stage2_27[25]},
      {stage2_28[1]},
      {stage3_29[5],stage3_28[5],stage3_27[18],stage3_26[30]}
   );
   gpc117_4 gpc8806 (
      {stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_27[26]},
      {stage2_28[2]},
      {stage3_29[6],stage3_28[6],stage3_27[19],stage3_26[31]}
   );
   gpc117_4 gpc8807 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[27]},
      {stage2_28[3]},
      {stage3_29[7],stage3_28[7],stage3_27[20],stage3_26[32]}
   );
   gpc117_4 gpc8808 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34]},
      {stage2_27[28]},
      {stage2_28[4]},
      {stage3_29[8],stage3_28[8],stage3_27[21],stage3_26[33]}
   );
   gpc117_4 gpc8809 (
      {stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage2_27[29]},
      {stage2_28[5]},
      {stage3_29[9],stage3_28[9],stage3_27[22],stage3_26[34]}
   );
   gpc117_4 gpc8810 (
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48]},
      {stage2_27[30]},
      {stage2_28[6]},
      {stage3_29[10],stage3_28[10],stage3_27[23],stage3_26[35]}
   );
   gpc117_4 gpc8811 (
      {stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55]},
      {stage2_27[31]},
      {stage2_28[7]},
      {stage3_29[11],stage3_28[11],stage3_27[24],stage3_26[36]}
   );
   gpc117_4 gpc8812 (
      {stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[32]},
      {stage2_28[8]},
      {stage3_29[12],stage3_28[12],stage3_27[25],stage3_26[37]}
   );
   gpc117_4 gpc8813 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69]},
      {stage2_27[33]},
      {stage2_28[9]},
      {stage3_29[13],stage3_28[13],stage3_27[26],stage3_26[38]}
   );
   gpc117_4 gpc8814 (
      {stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76]},
      {stage2_27[34]},
      {stage2_28[10]},
      {stage3_29[14],stage3_28[14],stage3_27[27],stage3_26[39]}
   );
   gpc117_4 gpc8815 (
      {stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage2_27[35]},
      {stage2_28[11]},
      {stage3_29[15],stage3_28[15],stage3_27[28],stage3_26[40]}
   );
   gpc117_4 gpc8816 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88], stage2_26[89], stage2_26[90]},
      {stage2_27[36]},
      {stage2_28[12]},
      {stage3_29[16],stage3_28[16],stage3_27[29],stage3_26[41]}
   );
   gpc117_4 gpc8817 (
      {stage2_26[91], stage2_26[92], stage2_26[93], stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97]},
      {stage2_27[37]},
      {stage2_28[13]},
      {stage3_29[17],stage3_28[17],stage3_27[30],stage3_26[42]}
   );
   gpc117_4 gpc8818 (
      {stage2_26[98], stage2_26[99], stage2_26[100], stage2_26[101], stage2_26[102], stage2_26[103], stage2_26[104]},
      {stage2_27[38]},
      {stage2_28[14]},
      {stage3_29[18],stage3_28[18],stage3_27[31],stage3_26[43]}
   );
   gpc117_4 gpc8819 (
      {stage2_26[105], stage2_26[106], stage2_26[107], stage2_26[108], stage2_26[109], stage2_26[110], stage2_26[111]},
      {stage2_27[39]},
      {stage2_28[15]},
      {stage3_29[19],stage3_28[19],stage3_27[32],stage3_26[44]}
   );
   gpc117_4 gpc8820 (
      {stage2_26[112], stage2_26[113], stage2_26[114], stage2_26[115], stage2_26[116], stage2_26[117], stage2_26[118]},
      {stage2_27[40]},
      {stage2_28[16]},
      {stage3_29[20],stage3_28[20],stage3_27[33],stage3_26[45]}
   );
   gpc117_4 gpc8821 (
      {stage2_26[119], stage2_26[120], stage2_26[121], stage2_26[122], stage2_26[123], stage2_26[124], stage2_26[125]},
      {stage2_27[41]},
      {stage2_28[17]},
      {stage3_29[21],stage3_28[21],stage3_27[34],stage3_26[46]}
   );
   gpc7_3 gpc8822 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48]},
      {stage3_29[22],stage3_28[22],stage3_27[35]}
   );
   gpc7_3 gpc8823 (
      {stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55]},
      {stage3_29[23],stage3_28[23],stage3_27[36]}
   );
   gpc207_4 gpc8824 (
      {stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_29[0], stage2_29[1]},
      {stage3_30[0],stage3_29[24],stage3_28[24],stage3_27[37]}
   );
   gpc207_4 gpc8825 (
      {stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_29[2], stage2_29[3]},
      {stage3_30[1],stage3_29[25],stage3_28[25],stage3_27[38]}
   );
   gpc606_5 gpc8826 (
      {stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73], stage2_27[74], stage2_27[75]},
      {stage2_29[4], stage2_29[5], stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9]},
      {stage3_31[0],stage3_30[2],stage3_29[26],stage3_28[26],stage3_27[39]}
   );
   gpc606_5 gpc8827 (
      {stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80], stage2_27[81]},
      {stage2_29[10], stage2_29[11], stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15]},
      {stage3_31[1],stage3_30[3],stage3_29[27],stage3_28[27],stage3_27[40]}
   );
   gpc615_5 gpc8828 (
      {stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], 1'b0},
      {stage2_28[18]},
      {stage2_29[16], stage2_29[17], stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage3_31[2],stage3_30[4],stage3_29[28],stage3_28[28],stage3_27[41]}
   );
   gpc615_5 gpc8829 (
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_29[22]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[5],stage3_29[29],stage3_28[29]}
   );
   gpc615_5 gpc8830 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[23]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[6],stage3_29[30],stage3_28[30]}
   );
   gpc615_5 gpc8831 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[24]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[7],stage3_29[31],stage3_28[31]}
   );
   gpc615_5 gpc8832 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[25]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[8],stage3_29[32],stage3_28[32]}
   );
   gpc615_5 gpc8833 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[26]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[7],stage3_30[9],stage3_29[33],stage3_28[33]}
   );
   gpc1163_5 gpc8834 (
      {stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[5],stage3_31[8],stage3_30[10],stage3_29[34]}
   );
   gpc1163_5 gpc8835 (
      {stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[6],stage3_31[9],stage3_30[11],stage3_29[35]}
   );
   gpc1163_5 gpc8836 (
      {stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[7],stage3_31[10],stage3_30[12],stage3_29[36]}
   );
   gpc1163_5 gpc8837 (
      {stage2_29[36], stage2_29[37], stage2_29[38]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[8],stage3_31[11],stage3_30[13],stage3_29[37]}
   );
   gpc1163_5 gpc8838 (
      {stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[9],stage3_31[12],stage3_30[14],stage3_29[38]}
   );
   gpc606_5 gpc8839 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[10],stage3_31[13],stage3_30[15],stage3_29[39]}
   );
   gpc606_5 gpc8840 (
      {stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[11],stage3_31[14],stage3_30[16],stage3_29[40]}
   );
   gpc606_5 gpc8841 (
      {stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[12],stage3_31[15],stage3_30[17],stage3_29[41]}
   );
   gpc606_5 gpc8842 (
      {stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[13],stage3_31[16],stage3_30[18],stage3_29[42]}
   );
   gpc606_5 gpc8843 (
      {stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[14],stage3_31[17],stage3_30[19],stage3_29[43]}
   );
   gpc606_5 gpc8844 (
      {stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[15],stage3_31[18],stage3_30[20],stage3_29[44]}
   );
   gpc606_5 gpc8845 (
      {stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[16],stage3_31[19],stage3_30[21],stage3_29[45]}
   );
   gpc606_5 gpc8846 (
      {stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[17],stage3_31[20],stage3_30[22],stage3_29[46]}
   );
   gpc606_5 gpc8847 (
      {stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[18],stage3_31[21],stage3_30[23],stage3_29[47]}
   );
   gpc606_5 gpc8848 (
      {stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101]},
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage3_33[14],stage3_32[19],stage3_31[22],stage3_30[24],stage3_29[48]}
   );
   gpc1163_5 gpc8849 (
      {stage2_30[60], stage2_30[61], stage2_30[62]},
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_32[5]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[15],stage3_32[20],stage3_31[23],stage3_30[25]}
   );
   gpc615_5 gpc8850 (
      {stage2_30[63], stage2_30[64], stage2_30[65], stage2_30[66], stage2_30[67]},
      {stage2_31[71]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[16],stage3_32[21],stage3_31[24],stage3_30[26]}
   );
   gpc615_5 gpc8851 (
      {stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71], stage2_30[72]},
      {stage2_31[72]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[17],stage3_32[22],stage3_31[25],stage3_30[27]}
   );
   gpc615_5 gpc8852 (
      {stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[73]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[18],stage3_32[23],stage3_31[26],stage3_30[28]}
   );
   gpc615_5 gpc8853 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82]},
      {stage2_31[74]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[19],stage3_32[24],stage3_31[27],stage3_30[29]}
   );
   gpc615_5 gpc8854 (
      {stage2_30[83], stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87]},
      {stage2_31[75]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[20],stage3_32[25],stage3_31[28],stage3_30[30]}
   );
   gpc615_5 gpc8855 (
      {stage2_30[88], stage2_30[89], stage2_30[90], stage2_30[91], stage2_30[92]},
      {stage2_31[76]},
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40], stage2_32[41]},
      {stage3_34[6],stage3_33[21],stage3_32[26],stage3_31[29],stage3_30[31]}
   );
   gpc606_5 gpc8856 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[0],stage3_34[7],stage3_33[22],stage3_32[27],stage3_31[30]}
   );
   gpc606_5 gpc8857 (
      {stage2_31[83], stage2_31[84], stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88]},
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12]},
      {stage3_35[1],stage3_34[8],stage3_33[23],stage3_32[28],stage3_31[31]}
   );
   gpc606_5 gpc8858 (
      {stage2_31[89], stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18]},
      {stage3_35[2],stage3_34[9],stage3_33[24],stage3_32[29],stage3_31[32]}
   );
   gpc606_5 gpc8859 (
      {stage2_31[95], stage2_31[96], stage2_31[97], stage2_31[98], stage2_31[99], stage2_31[100]},
      {stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24]},
      {stage3_35[3],stage3_34[10],stage3_33[25],stage3_32[30],stage3_31[33]}
   );
   gpc606_5 gpc8860 (
      {stage2_31[101], stage2_31[102], stage2_31[103], stage2_31[104], stage2_31[105], stage2_31[106]},
      {stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29], stage2_33[30]},
      {stage3_35[4],stage3_34[11],stage3_33[26],stage3_32[31],stage3_31[34]}
   );
   gpc606_5 gpc8861 (
      {stage2_31[107], stage2_31[108], stage2_31[109], stage2_31[110], stage2_31[111], stage2_31[112]},
      {stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35], stage2_33[36]},
      {stage3_35[5],stage3_34[12],stage3_33[27],stage3_32[32],stage3_31[35]}
   );
   gpc606_5 gpc8862 (
      {stage2_31[113], stage2_31[114], stage2_31[115], stage2_31[116], stage2_31[117], stage2_31[118]},
      {stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41], stage2_33[42]},
      {stage3_35[6],stage3_34[13],stage3_33[28],stage3_32[33],stage3_31[36]}
   );
   gpc615_5 gpc8863 (
      {stage2_31[119], stage2_31[120], stage2_31[121], stage2_31[122], stage2_31[123]},
      {stage2_32[42]},
      {stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48]},
      {stage3_35[7],stage3_34[14],stage3_33[29],stage3_32[34],stage3_31[37]}
   );
   gpc1163_5 gpc8864 (
      {stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54]},
      {stage2_34[0]},
      {stage2_35[0]},
      {stage3_36[0],stage3_35[8],stage3_34[15],stage3_33[30],stage3_32[35]}
   );
   gpc1163_5 gpc8865 (
      {stage2_32[46], stage2_32[47], stage2_32[48]},
      {stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59], stage2_33[60]},
      {stage2_34[1]},
      {stage2_35[1]},
      {stage3_36[1],stage3_35[9],stage3_34[16],stage3_33[31],stage3_32[36]}
   );
   gpc1163_5 gpc8866 (
      {stage2_32[49], stage2_32[50], stage2_32[51]},
      {stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65], stage2_33[66]},
      {stage2_34[2]},
      {stage2_35[2]},
      {stage3_36[2],stage3_35[10],stage3_34[17],stage3_33[32],stage3_32[37]}
   );
   gpc1163_5 gpc8867 (
      {stage2_32[52], stage2_32[53], stage2_32[54]},
      {stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71], stage2_33[72]},
      {stage2_34[3]},
      {stage2_35[3]},
      {stage3_36[3],stage3_35[11],stage3_34[18],stage3_33[33],stage3_32[38]}
   );
   gpc1163_5 gpc8868 (
      {stage2_32[55], stage2_32[56], stage2_32[57]},
      {stage2_33[73], stage2_33[74], stage2_33[75], stage2_33[76], stage2_33[77], stage2_33[78]},
      {stage2_34[4]},
      {stage2_35[4]},
      {stage3_36[4],stage3_35[12],stage3_34[19],stage3_33[34],stage3_32[39]}
   );
   gpc1163_5 gpc8869 (
      {stage2_32[58], stage2_32[59], stage2_32[60]},
      {stage2_33[79], stage2_33[80], stage2_33[81], stage2_33[82], stage2_33[83], stage2_33[84]},
      {stage2_34[5]},
      {stage2_35[5]},
      {stage3_36[5],stage3_35[13],stage3_34[20],stage3_33[35],stage3_32[40]}
   );
   gpc1163_5 gpc8870 (
      {stage2_32[61], stage2_32[62], stage2_32[63]},
      {stage2_33[85], stage2_33[86], stage2_33[87], stage2_33[88], stage2_33[89], stage2_33[90]},
      {stage2_34[6]},
      {stage2_35[6]},
      {stage3_36[6],stage3_35[14],stage3_34[21],stage3_33[36],stage3_32[41]}
   );
   gpc606_5 gpc8871 (
      {stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68], stage2_32[69]},
      {stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11], stage2_34[12]},
      {stage3_36[7],stage3_35[15],stage3_34[22],stage3_33[37],stage3_32[42]}
   );
   gpc606_5 gpc8872 (
      {stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74], stage2_32[75]},
      {stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17], stage2_34[18]},
      {stage3_36[8],stage3_35[16],stage3_34[23],stage3_33[38],stage3_32[43]}
   );
   gpc606_5 gpc8873 (
      {stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80], stage2_32[81]},
      {stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23], stage2_34[24]},
      {stage3_36[9],stage3_35[17],stage3_34[24],stage3_33[39],stage3_32[44]}
   );
   gpc606_5 gpc8874 (
      {stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86], stage2_32[87]},
      {stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29], stage2_34[30]},
      {stage3_36[10],stage3_35[18],stage3_34[25],stage3_33[40],stage3_32[45]}
   );
   gpc606_5 gpc8875 (
      {stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92], stage2_32[93]},
      {stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35], stage2_34[36]},
      {stage3_36[11],stage3_35[19],stage3_34[26],stage3_33[41],stage3_32[46]}
   );
   gpc606_5 gpc8876 (
      {stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98], stage2_32[99]},
      {stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41], stage2_34[42]},
      {stage3_36[12],stage3_35[20],stage3_34[27],stage3_33[42],stage3_32[47]}
   );
   gpc606_5 gpc8877 (
      {stage2_32[100], stage2_32[101], stage2_32[102], stage2_32[103], stage2_32[104], stage2_32[105]},
      {stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47], stage2_34[48]},
      {stage3_36[13],stage3_35[21],stage3_34[28],stage3_33[43],stage3_32[48]}
   );
   gpc606_5 gpc8878 (
      {stage2_32[106], stage2_32[107], stage2_32[108], stage2_32[109], stage2_32[110], stage2_32[111]},
      {stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53], stage2_34[54]},
      {stage3_36[14],stage3_35[22],stage3_34[29],stage3_33[44],stage3_32[49]}
   );
   gpc615_5 gpc8879 (
      {stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage2_35[7]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[15],stage3_35[23],stage3_34[30]}
   );
   gpc615_5 gpc8880 (
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64]},
      {stage2_35[8]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[1],stage3_36[16],stage3_35[24],stage3_34[31]}
   );
   gpc615_5 gpc8881 (
      {stage2_34[65], stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69]},
      {stage2_35[9]},
      {stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage3_38[2],stage3_37[2],stage3_36[17],stage3_35[25],stage3_34[32]}
   );
   gpc615_5 gpc8882 (
      {stage2_34[70], stage2_34[71], stage2_34[72], stage2_34[73], stage2_34[74]},
      {stage2_35[10]},
      {stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21], stage2_36[22], stage2_36[23]},
      {stage3_38[3],stage3_37[3],stage3_36[18],stage3_35[26],stage3_34[33]}
   );
   gpc615_5 gpc8883 (
      {stage2_34[75], stage2_34[76], stage2_34[77], stage2_34[78], stage2_34[79]},
      {stage2_35[11]},
      {stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27], stage2_36[28], stage2_36[29]},
      {stage3_38[4],stage3_37[4],stage3_36[19],stage3_35[27],stage3_34[34]}
   );
   gpc615_5 gpc8884 (
      {stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83], stage2_34[84]},
      {stage2_35[12]},
      {stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35]},
      {stage3_38[5],stage3_37[5],stage3_36[20],stage3_35[28],stage3_34[35]}
   );
   gpc615_5 gpc8885 (
      {stage2_34[85], stage2_34[86], stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[13]},
      {stage2_36[36], stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41]},
      {stage3_38[6],stage3_37[6],stage3_36[21],stage3_35[29],stage3_34[36]}
   );
   gpc615_5 gpc8886 (
      {stage2_34[90], stage2_34[91], stage2_34[92], stage2_34[93], stage2_34[94]},
      {stage2_35[14]},
      {stage2_36[42], stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47]},
      {stage3_38[7],stage3_37[7],stage3_36[22],stage3_35[30],stage3_34[37]}
   );
   gpc615_5 gpc8887 (
      {stage2_34[95], stage2_34[96], stage2_34[97], stage2_34[98], stage2_34[99]},
      {stage2_35[15]},
      {stage2_36[48], stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53]},
      {stage3_38[8],stage3_37[8],stage3_36[23],stage3_35[31],stage3_34[38]}
   );
   gpc615_5 gpc8888 (
      {stage2_34[100], stage2_34[101], stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[16]},
      {stage2_36[54], stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59]},
      {stage3_38[9],stage3_37[9],stage3_36[24],stage3_35[32],stage3_34[39]}
   );
   gpc615_5 gpc8889 (
      {stage2_34[105], stage2_34[106], stage2_34[107], stage2_34[108], stage2_34[109]},
      {stage2_35[17]},
      {stage2_36[60], stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65]},
      {stage3_38[10],stage3_37[10],stage3_36[25],stage3_35[33],stage3_34[40]}
   );
   gpc615_5 gpc8890 (
      {stage2_34[110], stage2_34[111], stage2_34[112], stage2_34[113], stage2_34[114]},
      {stage2_35[18]},
      {stage2_36[66], stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71]},
      {stage3_38[11],stage3_37[11],stage3_36[26],stage3_35[34],stage3_34[41]}
   );
   gpc615_5 gpc8891 (
      {stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118], stage2_34[119]},
      {stage2_35[19]},
      {stage2_36[72], stage2_36[73], stage2_36[74], stage2_36[75], stage2_36[76], stage2_36[77]},
      {stage3_38[12],stage3_37[12],stage3_36[27],stage3_35[35],stage3_34[42]}
   );
   gpc615_5 gpc8892 (
      {stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123], stage2_34[124]},
      {stage2_35[20]},
      {stage2_36[78], stage2_36[79], stage2_36[80], stage2_36[81], stage2_36[82], stage2_36[83]},
      {stage3_38[13],stage3_37[13],stage3_36[28],stage3_35[36],stage3_34[43]}
   );
   gpc615_5 gpc8893 (
      {stage2_34[125], stage2_34[126], stage2_34[127], 1'b0, 1'b0},
      {stage2_35[21]},
      {stage2_36[84], stage2_36[85], stage2_36[86], stage2_36[87], stage2_36[88], stage2_36[89]},
      {stage3_38[14],stage3_37[14],stage3_36[29],stage3_35[37],stage3_34[44]}
   );
   gpc606_5 gpc8894 (
      {stage2_35[22], stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[15],stage3_37[15],stage3_36[30],stage3_35[38]}
   );
   gpc615_5 gpc8895 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[90]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[16],stage3_37[16],stage3_36[31],stage3_35[39]}
   );
   gpc615_5 gpc8896 (
      {stage2_35[33], stage2_35[34], stage2_35[35], stage2_35[36], stage2_35[37]},
      {stage2_36[91]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[17],stage3_37[17],stage3_36[32],stage3_35[40]}
   );
   gpc615_5 gpc8897 (
      {stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41], stage2_35[42]},
      {stage2_36[92]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[18],stage3_37[18],stage3_36[33],stage3_35[41]}
   );
   gpc615_5 gpc8898 (
      {stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[93]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[19],stage3_37[19],stage3_36[34],stage3_35[42]}
   );
   gpc615_5 gpc8899 (
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52]},
      {stage2_36[94]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[20],stage3_37[20],stage3_36[35],stage3_35[43]}
   );
   gpc615_5 gpc8900 (
      {stage2_35[53], stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57]},
      {stage2_36[95]},
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage3_39[6],stage3_38[21],stage3_37[21],stage3_36[36],stage3_35[44]}
   );
   gpc615_5 gpc8901 (
      {stage2_35[58], stage2_35[59], stage2_35[60], stage2_35[61], stage2_35[62]},
      {stage2_36[96]},
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage3_39[7],stage3_38[22],stage3_37[22],stage3_36[37],stage3_35[45]}
   );
   gpc615_5 gpc8902 (
      {stage2_35[63], stage2_35[64], stage2_35[65], stage2_35[66], stage2_35[67]},
      {stage2_36[97]},
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage3_39[8],stage3_38[23],stage3_37[23],stage3_36[38],stage3_35[46]}
   );
   gpc615_5 gpc8903 (
      {stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71], stage2_35[72]},
      {stage2_36[98]},
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58], stage2_37[59]},
      {stage3_39[9],stage3_38[24],stage3_37[24],stage3_36[39],stage3_35[47]}
   );
   gpc615_5 gpc8904 (
      {stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[99]},
      {stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63], stage2_37[64], stage2_37[65]},
      {stage3_39[10],stage3_38[25],stage3_37[25],stage3_36[40],stage3_35[48]}
   );
   gpc615_5 gpc8905 (
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82]},
      {stage2_36[100]},
      {stage2_37[66], stage2_37[67], stage2_37[68], stage2_37[69], stage2_37[70], stage2_37[71]},
      {stage3_39[11],stage3_38[26],stage3_37[26],stage3_36[41],stage3_35[49]}
   );
   gpc615_5 gpc8906 (
      {stage2_35[83], stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87]},
      {stage2_36[101]},
      {stage2_37[72], stage2_37[73], stage2_37[74], stage2_37[75], stage2_37[76], stage2_37[77]},
      {stage3_39[12],stage3_38[27],stage3_37[27],stage3_36[42],stage3_35[50]}
   );
   gpc615_5 gpc8907 (
      {stage2_35[88], stage2_35[89], stage2_35[90], stage2_35[91], stage2_35[92]},
      {stage2_36[102]},
      {stage2_37[78], stage2_37[79], stage2_37[80], stage2_37[81], stage2_37[82], stage2_37[83]},
      {stage3_39[13],stage3_38[28],stage3_37[28],stage3_36[43],stage3_35[51]}
   );
   gpc615_5 gpc8908 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97]},
      {stage2_36[103]},
      {stage2_37[84], stage2_37[85], stage2_37[86], stage2_37[87], stage2_37[88], stage2_37[89]},
      {stage3_39[14],stage3_38[29],stage3_37[29],stage3_36[44],stage3_35[52]}
   );
   gpc615_5 gpc8909 (
      {stage2_35[98], stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102]},
      {stage2_36[104]},
      {stage2_37[90], stage2_37[91], stage2_37[92], stage2_37[93], stage2_37[94], stage2_37[95]},
      {stage3_39[15],stage3_38[30],stage3_37[30],stage3_36[45],stage3_35[53]}
   );
   gpc615_5 gpc8910 (
      {stage2_35[103], stage2_35[104], stage2_35[105], stage2_35[106], stage2_35[107]},
      {stage2_36[105]},
      {stage2_37[96], stage2_37[97], stage2_37[98], stage2_37[99], stage2_37[100], stage2_37[101]},
      {stage3_39[16],stage3_38[31],stage3_37[31],stage3_36[46],stage3_35[54]}
   );
   gpc615_5 gpc8911 (
      {stage2_35[108], stage2_35[109], stage2_35[110], stage2_35[111], stage2_35[112]},
      {stage2_36[106]},
      {stage2_37[102], stage2_37[103], stage2_37[104], stage2_37[105], stage2_37[106], stage2_37[107]},
      {stage3_39[17],stage3_38[32],stage3_37[32],stage3_36[47],stage3_35[55]}
   );
   gpc615_5 gpc8912 (
      {stage2_35[113], stage2_35[114], stage2_35[115], stage2_35[116], stage2_35[117]},
      {stage2_36[107]},
      {stage2_37[108], stage2_37[109], stage2_37[110], stage2_37[111], stage2_37[112], stage2_37[113]},
      {stage3_39[18],stage3_38[33],stage3_37[33],stage3_36[48],stage3_35[56]}
   );
   gpc606_5 gpc8913 (
      {stage2_36[108], stage2_36[109], stage2_36[110], stage2_36[111], stage2_36[112], stage2_36[113]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[19],stage3_38[34],stage3_37[34],stage3_36[49]}
   );
   gpc615_5 gpc8914 (
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10]},
      {stage2_39[0]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[1],stage3_39[20],stage3_38[35]}
   );
   gpc615_5 gpc8915 (
      {stage2_38[11], stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15]},
      {stage2_39[1]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[1],stage3_40[2],stage3_39[21],stage3_38[36]}
   );
   gpc615_5 gpc8916 (
      {stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_39[2]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[2],stage3_40[3],stage3_39[22],stage3_38[37]}
   );
   gpc615_5 gpc8917 (
      {stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage2_39[3]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[3],stage3_40[4],stage3_39[23],stage3_38[38]}
   );
   gpc615_5 gpc8918 (
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30]},
      {stage2_39[4]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[4],stage3_40[5],stage3_39[24],stage3_38[39]}
   );
   gpc615_5 gpc8919 (
      {stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage2_39[5]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[5],stage3_40[6],stage3_39[25],stage3_38[40]}
   );
   gpc615_5 gpc8920 (
      {stage2_38[36], stage2_38[37], stage2_38[38], stage2_38[39], stage2_38[40]},
      {stage2_39[6]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[6],stage3_40[7],stage3_39[26],stage3_38[41]}
   );
   gpc615_5 gpc8921 (
      {stage2_38[41], stage2_38[42], stage2_38[43], stage2_38[44], stage2_38[45]},
      {stage2_39[7]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[7],stage3_40[8],stage3_39[27],stage3_38[42]}
   );
   gpc615_5 gpc8922 (
      {stage2_38[46], stage2_38[47], stage2_38[48], stage2_38[49], stage2_38[50]},
      {stage2_39[8]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[8],stage3_40[9],stage3_39[28],stage3_38[43]}
   );
   gpc615_5 gpc8923 (
      {stage2_38[51], stage2_38[52], stage2_38[53], stage2_38[54], stage2_38[55]},
      {stage2_39[9]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[9],stage3_40[10],stage3_39[29],stage3_38[44]}
   );
   gpc615_5 gpc8924 (
      {stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59], stage2_38[60]},
      {stage2_39[10]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[10],stage3_40[11],stage3_39[30],stage3_38[45]}
   );
   gpc615_5 gpc8925 (
      {stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_39[11]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[11],stage3_40[12],stage3_39[31],stage3_38[46]}
   );
   gpc615_5 gpc8926 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70]},
      {stage2_39[12]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[12],stage3_40[13],stage3_39[32],stage3_38[47]}
   );
   gpc615_5 gpc8927 (
      {stage2_38[71], stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75]},
      {stage2_39[13]},
      {stage2_40[78], stage2_40[79], stage2_40[80], stage2_40[81], stage2_40[82], stage2_40[83]},
      {stage3_42[13],stage3_41[13],stage3_40[14],stage3_39[33],stage3_38[48]}
   );
   gpc615_5 gpc8928 (
      {stage2_38[76], stage2_38[77], stage2_38[78], stage2_38[79], stage2_38[80]},
      {stage2_39[14]},
      {stage2_40[84], stage2_40[85], stage2_40[86], stage2_40[87], stage2_40[88], stage2_40[89]},
      {stage3_42[14],stage3_41[14],stage3_40[15],stage3_39[34],stage3_38[49]}
   );
   gpc615_5 gpc8929 (
      {stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_40[90]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[15],stage3_41[15],stage3_40[16],stage3_39[35]}
   );
   gpc615_5 gpc8930 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24]},
      {stage2_40[91]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[16],stage3_41[16],stage3_40[17],stage3_39[36]}
   );
   gpc615_5 gpc8931 (
      {stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage2_40[92]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[17],stage3_41[17],stage3_40[18],stage3_39[37]}
   );
   gpc615_5 gpc8932 (
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34]},
      {stage2_40[93]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[18],stage3_41[18],stage3_40[19],stage3_39[38]}
   );
   gpc615_5 gpc8933 (
      {stage2_39[35], stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39]},
      {stage2_40[94]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[19],stage3_41[19],stage3_40[20],stage3_39[39]}
   );
   gpc615_5 gpc8934 (
      {stage2_39[40], stage2_39[41], stage2_39[42], stage2_39[43], stage2_39[44]},
      {stage2_40[95]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[20],stage3_41[20],stage3_40[21],stage3_39[40]}
   );
   gpc615_5 gpc8935 (
      {stage2_39[45], stage2_39[46], stage2_39[47], stage2_39[48], stage2_39[49]},
      {stage2_40[96]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[21],stage3_41[21],stage3_40[22],stage3_39[41]}
   );
   gpc615_5 gpc8936 (
      {stage2_39[50], stage2_39[51], stage2_39[52], stage2_39[53], stage2_39[54]},
      {stage2_40[97]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[22],stage3_41[22],stage3_40[23],stage3_39[42]}
   );
   gpc615_5 gpc8937 (
      {stage2_39[55], stage2_39[56], stage2_39[57], stage2_39[58], stage2_39[59]},
      {stage2_40[98]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[23],stage3_41[23],stage3_40[24],stage3_39[43]}
   );
   gpc615_5 gpc8938 (
      {stage2_39[60], stage2_39[61], stage2_39[62], stage2_39[63], stage2_39[64]},
      {stage2_40[99]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[24],stage3_41[24],stage3_40[25],stage3_39[44]}
   );
   gpc615_5 gpc8939 (
      {stage2_39[65], stage2_39[66], stage2_39[67], stage2_39[68], stage2_39[69]},
      {stage2_40[100]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[25],stage3_41[25],stage3_40[26],stage3_39[45]}
   );
   gpc615_5 gpc8940 (
      {stage2_39[70], stage2_39[71], stage2_39[72], stage2_39[73], stage2_39[74]},
      {stage2_40[101]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[26],stage3_41[26],stage3_40[27],stage3_39[46]}
   );
   gpc615_5 gpc8941 (
      {stage2_39[75], stage2_39[76], stage2_39[77], stage2_39[78], stage2_39[79]},
      {stage2_40[102]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[27],stage3_41[27],stage3_40[28],stage3_39[47]}
   );
   gpc615_5 gpc8942 (
      {stage2_39[80], stage2_39[81], stage2_39[82], stage2_39[83], stage2_39[84]},
      {stage2_40[103]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[28],stage3_41[28],stage3_40[29],stage3_39[48]}
   );
   gpc615_5 gpc8943 (
      {stage2_39[85], stage2_39[86], stage2_39[87], stage2_39[88], stage2_39[89]},
      {stage2_40[104]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[29],stage3_41[29],stage3_40[30],stage3_39[49]}
   );
   gpc615_5 gpc8944 (
      {stage2_39[90], stage2_39[91], stage2_39[92], stage2_39[93], stage2_39[94]},
      {stage2_40[105]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[30],stage3_41[30],stage3_40[31],stage3_39[50]}
   );
   gpc615_5 gpc8945 (
      {stage2_39[95], stage2_39[96], stage2_39[97], stage2_39[98], stage2_39[99]},
      {stage2_40[106]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[31],stage3_41[31],stage3_40[32],stage3_39[51]}
   );
   gpc606_5 gpc8946 (
      {stage2_40[107], stage2_40[108], stage2_40[109], stage2_40[110], stage2_40[111], stage2_40[112]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[32],stage3_41[32],stage3_40[33]}
   );
   gpc606_5 gpc8947 (
      {stage2_40[113], stage2_40[114], stage2_40[115], stage2_40[116], stage2_40[117], stage2_40[118]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[33],stage3_41[33],stage3_40[34]}
   );
   gpc606_5 gpc8948 (
      {stage2_40[119], stage2_40[120], stage2_40[121], stage2_40[122], stage2_40[123], stage2_40[124]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[19],stage3_42[34],stage3_41[34],stage3_40[35]}
   );
   gpc606_5 gpc8949 (
      {stage2_40[125], stage2_40[126], stage2_40[127], stage2_40[128], stage2_40[129], stage2_40[130]},
      {stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21], stage2_42[22], stage2_42[23]},
      {stage3_44[3],stage3_43[20],stage3_42[35],stage3_41[35],stage3_40[36]}
   );
   gpc615_5 gpc8950 (
      {stage2_42[24], stage2_42[25], stage2_42[26], stage2_42[27], stage2_42[28]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[21],stage3_42[36]}
   );
   gpc615_5 gpc8951 (
      {stage2_42[29], stage2_42[30], stage2_42[31], stage2_42[32], stage2_42[33]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[22],stage3_42[37]}
   );
   gpc615_5 gpc8952 (
      {stage2_42[34], stage2_42[35], stage2_42[36], stage2_42[37], stage2_42[38]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[6],stage3_43[23],stage3_42[38]}
   );
   gpc615_5 gpc8953 (
      {stage2_42[39], stage2_42[40], stage2_42[41], stage2_42[42], stage2_42[43]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[7],stage3_43[24],stage3_42[39]}
   );
   gpc615_5 gpc8954 (
      {stage2_42[44], stage2_42[45], stage2_42[46], stage2_42[47], stage2_42[48]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[8],stage3_43[25],stage3_42[40]}
   );
   gpc615_5 gpc8955 (
      {stage2_42[49], stage2_42[50], stage2_42[51], stage2_42[52], stage2_42[53]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[9],stage3_43[26],stage3_42[41]}
   );
   gpc615_5 gpc8956 (
      {stage2_42[54], stage2_42[55], stage2_42[56], stage2_42[57], stage2_42[58]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[10],stage3_43[27],stage3_42[42]}
   );
   gpc615_5 gpc8957 (
      {stage2_42[59], stage2_42[60], stage2_42[61], stage2_42[62], stage2_42[63]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[11],stage3_43[28],stage3_42[43]}
   );
   gpc615_5 gpc8958 (
      {stage2_42[64], stage2_42[65], stage2_42[66], stage2_42[67], stage2_42[68]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[12],stage3_43[29],stage3_42[44]}
   );
   gpc615_5 gpc8959 (
      {stage2_42[69], stage2_42[70], stage2_42[71], stage2_42[72], stage2_42[73]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[13],stage3_43[30],stage3_42[45]}
   );
   gpc606_5 gpc8960 (
      {stage2_43[10], stage2_43[11], stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[10],stage3_45[10],stage3_44[14],stage3_43[31]}
   );
   gpc606_5 gpc8961 (
      {stage2_43[16], stage2_43[17], stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[11],stage3_45[11],stage3_44[15],stage3_43[32]}
   );
   gpc606_5 gpc8962 (
      {stage2_43[22], stage2_43[23], stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[12],stage3_45[12],stage3_44[16],stage3_43[33]}
   );
   gpc606_5 gpc8963 (
      {stage2_43[28], stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[13],stage3_45[13],stage3_44[17],stage3_43[34]}
   );
   gpc606_5 gpc8964 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38], stage2_43[39]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[14],stage3_45[14],stage3_44[18],stage3_43[35]}
   );
   gpc606_5 gpc8965 (
      {stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[15],stage3_45[15],stage3_44[19],stage3_43[36]}
   );
   gpc606_5 gpc8966 (
      {stage2_43[46], stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[16],stage3_45[16],stage3_44[20],stage3_43[37]}
   );
   gpc606_5 gpc8967 (
      {stage2_43[52], stage2_43[53], stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[17],stage3_45[17],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc8968 (
      {stage2_43[58], stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62]},
      {stage2_44[60]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[18],stage3_45[18],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc8969 (
      {stage2_43[63], stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67]},
      {stage2_44[61]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[19],stage3_45[19],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc8970 (
      {stage2_43[68], stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72]},
      {stage2_44[62]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[20],stage3_45[20],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc8971 (
      {stage2_43[73], stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77]},
      {stage2_44[63]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[21],stage3_45[21],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc8972 (
      {stage2_43[78], stage2_43[79], stage2_43[80], stage2_43[81], stage2_43[82]},
      {stage2_44[64]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[22],stage3_45[22],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc8973 (
      {stage2_43[83], stage2_43[84], stage2_43[85], stage2_43[86], stage2_43[87]},
      {stage2_44[65]},
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage3_47[13],stage3_46[23],stage3_45[23],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc8974 (
      {stage2_43[88], stage2_43[89], stage2_43[90], stage2_43[91], stage2_43[92]},
      {stage2_44[66]},
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage3_47[14],stage3_46[24],stage3_45[24],stage3_44[28],stage3_43[45]}
   );
   gpc615_5 gpc8975 (
      {stage2_43[93], stage2_43[94], stage2_43[95], stage2_43[96], stage2_43[97]},
      {stage2_44[67]},
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage3_47[15],stage3_46[25],stage3_45[25],stage3_44[29],stage3_43[46]}
   );
   gpc606_5 gpc8976 (
      {stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71], stage2_44[72], stage2_44[73]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[16],stage3_46[26],stage3_45[26],stage3_44[30]}
   );
   gpc606_5 gpc8977 (
      {stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77], stage2_44[78], stage2_44[79]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[17],stage3_46[27],stage3_45[27],stage3_44[31]}
   );
   gpc606_5 gpc8978 (
      {stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83], stage2_44[84], stage2_44[85]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[18],stage3_46[28],stage3_45[28],stage3_44[32]}
   );
   gpc606_5 gpc8979 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[3],stage3_47[19],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc8980 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[4],stage3_47[20],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc8981 (
      {stage2_45[108], stage2_45[109], stage2_45[110], stage2_45[111], stage2_45[112], stage2_45[113]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[5],stage3_47[21],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc8982 (
      {stage2_45[114], stage2_45[115], stage2_45[116], stage2_45[117], stage2_45[118], stage2_45[119]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[6],stage3_47[22],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc8983 (
      {stage2_45[120], stage2_45[121], stage2_45[122], stage2_45[123], stage2_45[124], stage2_45[125]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[7],stage3_47[23],stage3_46[33],stage3_45[33]}
   );
   gpc615_5 gpc8984 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[30]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[5],stage3_48[8],stage3_47[24],stage3_46[34]}
   );
   gpc615_5 gpc8985 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[31]},
      {stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage3_50[1],stage3_49[6],stage3_48[9],stage3_47[25],stage3_46[35]}
   );
   gpc615_5 gpc8986 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[32]},
      {stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17]},
      {stage3_50[2],stage3_49[7],stage3_48[10],stage3_47[26],stage3_46[36]}
   );
   gpc615_5 gpc8987 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[33]},
      {stage2_48[18], stage2_48[19], stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23]},
      {stage3_50[3],stage3_49[8],stage3_48[11],stage3_47[27],stage3_46[37]}
   );
   gpc615_5 gpc8988 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[34]},
      {stage2_48[24], stage2_48[25], stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29]},
      {stage3_50[4],stage3_49[9],stage3_48[12],stage3_47[28],stage3_46[38]}
   );
   gpc615_5 gpc8989 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[35]},
      {stage2_48[30], stage2_48[31], stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35]},
      {stage3_50[5],stage3_49[10],stage3_48[13],stage3_47[29],stage3_46[39]}
   );
   gpc615_5 gpc8990 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[36]},
      {stage2_48[36], stage2_48[37], stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41]},
      {stage3_50[6],stage3_49[11],stage3_48[14],stage3_47[30],stage3_46[40]}
   );
   gpc615_5 gpc8991 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[37]},
      {stage2_48[42], stage2_48[43], stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47]},
      {stage3_50[7],stage3_49[12],stage3_48[15],stage3_47[31],stage3_46[41]}
   );
   gpc615_5 gpc8992 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[38]},
      {stage2_48[48], stage2_48[49], stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53]},
      {stage3_50[8],stage3_49[13],stage3_48[16],stage3_47[32],stage3_46[42]}
   );
   gpc615_5 gpc8993 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[39]},
      {stage2_48[54], stage2_48[55], stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59]},
      {stage3_50[9],stage3_49[14],stage3_48[17],stage3_47[33],stage3_46[43]}
   );
   gpc615_5 gpc8994 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[40]},
      {stage2_48[60], stage2_48[61], stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65]},
      {stage3_50[10],stage3_49[15],stage3_48[18],stage3_47[34],stage3_46[44]}
   );
   gpc615_5 gpc8995 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[41]},
      {stage2_48[66], stage2_48[67], stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71]},
      {stage3_50[11],stage3_49[16],stage3_48[19],stage3_47[35],stage3_46[45]}
   );
   gpc615_5 gpc8996 (
      {stage2_46[78], stage2_46[79], stage2_46[80], stage2_46[81], stage2_46[82]},
      {stage2_47[42]},
      {stage2_48[72], stage2_48[73], stage2_48[74], stage2_48[75], stage2_48[76], stage2_48[77]},
      {stage3_50[12],stage3_49[17],stage3_48[20],stage3_47[36],stage3_46[46]}
   );
   gpc615_5 gpc8997 (
      {stage2_46[83], stage2_46[84], stage2_46[85], stage2_46[86], stage2_46[87]},
      {stage2_47[43]},
      {stage2_48[78], stage2_48[79], stage2_48[80], stage2_48[81], stage2_48[82], stage2_48[83]},
      {stage3_50[13],stage3_49[18],stage3_48[21],stage3_47[37],stage3_46[47]}
   );
   gpc615_5 gpc8998 (
      {stage2_46[88], stage2_46[89], stage2_46[90], stage2_46[91], stage2_46[92]},
      {stage2_47[44]},
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage3_50[14],stage3_49[19],stage3_48[22],stage3_47[38],stage3_46[48]}
   );
   gpc1163_5 gpc8999 (
      {stage2_47[45], stage2_47[46], stage2_47[47]},
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_49[0]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[15],stage3_49[20],stage3_48[23],stage3_47[39]}
   );
   gpc1163_5 gpc9000 (
      {stage2_47[48], stage2_47[49], stage2_47[50]},
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_49[1]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[16],stage3_49[21],stage3_48[24],stage3_47[40]}
   );
   gpc1163_5 gpc9001 (
      {stage2_47[51], stage2_47[52], stage2_47[53]},
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_49[2]},
      {stage2_50[2]},
      {stage3_51[2],stage3_50[17],stage3_49[22],stage3_48[25],stage3_47[41]}
   );
   gpc1163_5 gpc9002 (
      {stage2_47[54], stage2_47[55], stage2_47[56]},
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_49[3]},
      {stage2_50[3]},
      {stage3_51[3],stage3_50[18],stage3_49[23],stage3_48[26],stage3_47[42]}
   );
   gpc1163_5 gpc9003 (
      {stage2_47[57], stage2_47[58], stage2_47[59]},
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_49[4]},
      {stage2_50[4]},
      {stage3_51[4],stage3_50[19],stage3_49[24],stage3_48[27],stage3_47[43]}
   );
   gpc1163_5 gpc9004 (
      {stage2_47[60], stage2_47[61], stage2_47[62]},
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_49[5]},
      {stage2_50[5]},
      {stage3_51[5],stage3_50[20],stage3_49[25],stage3_48[28],stage3_47[44]}
   );
   gpc615_5 gpc9005 (
      {stage2_47[63], stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67]},
      {stage2_48[126]},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[6],stage3_50[21],stage3_49[26],stage3_48[29],stage3_47[45]}
   );
   gpc615_5 gpc9006 (
      {stage2_47[68], stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72]},
      {stage2_48[127]},
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage3_51[7],stage3_50[22],stage3_49[27],stage3_48[30],stage3_47[46]}
   );
   gpc615_5 gpc9007 (
      {stage2_47[73], stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77]},
      {stage2_48[128]},
      {stage2_49[18], stage2_49[19], stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23]},
      {stage3_51[8],stage3_50[23],stage3_49[28],stage3_48[31],stage3_47[47]}
   );
   gpc615_5 gpc9008 (
      {stage2_47[78], stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82]},
      {stage2_48[129]},
      {stage2_49[24], stage2_49[25], stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29]},
      {stage3_51[9],stage3_50[24],stage3_49[29],stage3_48[32],stage3_47[48]}
   );
   gpc606_5 gpc9009 (
      {stage2_48[130], stage2_48[131], stage2_48[132], stage2_48[133], stage2_48[134], stage2_48[135]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[0],stage3_51[10],stage3_50[25],stage3_49[30],stage3_48[33]}
   );
   gpc606_5 gpc9010 (
      {stage2_48[136], stage2_48[137], stage2_48[138], stage2_48[139], stage2_48[140], stage2_48[141]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[1],stage3_51[11],stage3_50[26],stage3_49[31],stage3_48[34]}
   );
   gpc606_5 gpc9011 (
      {stage2_48[142], stage2_48[143], stage2_48[144], stage2_48[145], stage2_48[146], stage2_48[147]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[2],stage3_51[12],stage3_50[27],stage3_49[32],stage3_48[35]}
   );
   gpc606_5 gpc9012 (
      {stage2_48[148], stage2_48[149], stage2_48[150], stage2_48[151], stage2_48[152], stage2_48[153]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[3],stage3_51[13],stage3_50[28],stage3_49[33],stage3_48[36]}
   );
   gpc606_5 gpc9013 (
      {stage2_49[30], stage2_49[31], stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[4],stage3_51[14],stage3_50[29],stage3_49[34]}
   );
   gpc606_5 gpc9014 (
      {stage2_49[36], stage2_49[37], stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[5],stage3_51[15],stage3_50[30],stage3_49[35]}
   );
   gpc606_5 gpc9015 (
      {stage2_49[42], stage2_49[43], stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[6],stage3_51[16],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc9016 (
      {stage2_49[48], stage2_49[49], stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[7],stage3_51[17],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc9017 (
      {stage2_49[54], stage2_49[55], stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[8],stage3_51[18],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc9018 (
      {stage2_49[60], stage2_49[61], stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[9],stage3_51[19],stage3_50[34],stage3_49[39]}
   );
   gpc606_5 gpc9019 (
      {stage2_49[66], stage2_49[67], stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71]},
      {stage2_51[36], stage2_51[37], stage2_51[38], stage2_51[39], stage2_51[40], stage2_51[41]},
      {stage3_53[6],stage3_52[10],stage3_51[20],stage3_50[35],stage3_49[40]}
   );
   gpc606_5 gpc9020 (
      {stage2_49[72], stage2_49[73], stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77]},
      {stage2_51[42], stage2_51[43], stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47]},
      {stage3_53[7],stage3_52[11],stage3_51[21],stage3_50[36],stage3_49[41]}
   );
   gpc606_5 gpc9021 (
      {stage2_49[78], stage2_49[79], stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83]},
      {stage2_51[48], stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage3_53[8],stage3_52[12],stage3_51[22],stage3_50[37],stage3_49[42]}
   );
   gpc606_5 gpc9022 (
      {stage2_49[84], stage2_49[85], stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89]},
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58], stage2_51[59]},
      {stage3_53[9],stage3_52[13],stage3_51[23],stage3_50[38],stage3_49[43]}
   );
   gpc606_5 gpc9023 (
      {stage2_49[90], stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_51[60], stage2_51[61], stage2_51[62], stage2_51[63], stage2_51[64], stage2_51[65]},
      {stage3_53[10],stage3_52[14],stage3_51[24],stage3_50[39],stage3_49[44]}
   );
   gpc2135_5 gpc9024 (
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34]},
      {stage2_51[66], stage2_51[67], stage2_51[68]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[11],stage3_52[15],stage3_51[25],stage3_50[40]}
   );
   gpc1406_5 gpc9025 (
      {stage2_50[35], stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40]},
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4]},
      {stage2_53[2]},
      {stage3_54[1],stage3_53[12],stage3_52[16],stage3_51[26],stage3_50[41]}
   );
   gpc1406_5 gpc9026 (
      {stage2_50[41], stage2_50[42], stage2_50[43], stage2_50[44], stage2_50[45], stage2_50[46]},
      {stage2_52[5], stage2_52[6], stage2_52[7], stage2_52[8]},
      {stage2_53[3]},
      {stage3_54[2],stage3_53[13],stage3_52[17],stage3_51[27],stage3_50[42]}
   );
   gpc1406_5 gpc9027 (
      {stage2_50[47], stage2_50[48], stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52]},
      {stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12]},
      {stage2_53[4]},
      {stage3_54[3],stage3_53[14],stage3_52[18],stage3_51[28],stage3_50[43]}
   );
   gpc606_5 gpc9028 (
      {stage2_50[53], stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17], stage2_52[18]},
      {stage3_54[4],stage3_53[15],stage3_52[19],stage3_51[29],stage3_50[44]}
   );
   gpc606_5 gpc9029 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63], stage2_50[64]},
      {stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23], stage2_52[24]},
      {stage3_54[5],stage3_53[16],stage3_52[20],stage3_51[30],stage3_50[45]}
   );
   gpc606_5 gpc9030 (
      {stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68], stage2_50[69], stage2_50[70]},
      {stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29], stage2_52[30]},
      {stage3_54[6],stage3_53[17],stage3_52[21],stage3_51[31],stage3_50[46]}
   );
   gpc606_5 gpc9031 (
      {stage2_50[71], stage2_50[72], stage2_50[73], stage2_50[74], stage2_50[75], stage2_50[76]},
      {stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35], stage2_52[36]},
      {stage3_54[7],stage3_53[18],stage3_52[22],stage3_51[32],stage3_50[47]}
   );
   gpc606_5 gpc9032 (
      {stage2_50[77], stage2_50[78], stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82]},
      {stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41], stage2_52[42]},
      {stage3_54[8],stage3_53[19],stage3_52[23],stage3_51[33],stage3_50[48]}
   );
   gpc606_5 gpc9033 (
      {stage2_50[83], stage2_50[84], stage2_50[85], stage2_50[86], stage2_50[87], stage2_50[88]},
      {stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47], stage2_52[48]},
      {stage3_54[9],stage3_53[20],stage3_52[24],stage3_51[34],stage3_50[49]}
   );
   gpc606_5 gpc9034 (
      {stage2_50[89], stage2_50[90], stage2_50[91], stage2_50[92], stage2_50[93], stage2_50[94]},
      {stage2_52[49], stage2_52[50], stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54]},
      {stage3_54[10],stage3_53[21],stage3_52[25],stage3_51[35],stage3_50[50]}
   );
   gpc606_5 gpc9035 (
      {stage2_50[95], stage2_50[96], stage2_50[97], stage2_50[98], stage2_50[99], stage2_50[100]},
      {stage2_52[55], stage2_52[56], stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60]},
      {stage3_54[11],stage3_53[22],stage3_52[26],stage3_51[36],stage3_50[51]}
   );
   gpc606_5 gpc9036 (
      {stage2_50[101], stage2_50[102], stage2_50[103], stage2_50[104], stage2_50[105], stage2_50[106]},
      {stage2_52[61], stage2_52[62], stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66]},
      {stage3_54[12],stage3_53[23],stage3_52[27],stage3_51[37],stage3_50[52]}
   );
   gpc606_5 gpc9037 (
      {stage2_50[107], stage2_50[108], stage2_50[109], stage2_50[110], stage2_50[111], stage2_50[112]},
      {stage2_52[67], stage2_52[68], stage2_52[69], stage2_52[70], stage2_52[71], stage2_52[72]},
      {stage3_54[13],stage3_53[24],stage3_52[28],stage3_51[38],stage3_50[53]}
   );
   gpc606_5 gpc9038 (
      {stage2_50[113], stage2_50[114], stage2_50[115], stage2_50[116], stage2_50[117], stage2_50[118]},
      {stage2_52[73], stage2_52[74], stage2_52[75], stage2_52[76], stage2_52[77], stage2_52[78]},
      {stage3_54[14],stage3_53[25],stage3_52[29],stage3_51[39],stage3_50[54]}
   );
   gpc606_5 gpc9039 (
      {stage2_50[119], stage2_50[120], stage2_50[121], stage2_50[122], stage2_50[123], stage2_50[124]},
      {stage2_52[79], stage2_52[80], stage2_52[81], stage2_52[82], stage2_52[83], stage2_52[84]},
      {stage3_54[15],stage3_53[26],stage3_52[30],stage3_51[40],stage3_50[55]}
   );
   gpc606_5 gpc9040 (
      {stage2_50[125], stage2_50[126], stage2_50[127], stage2_50[128], stage2_50[129], stage2_50[130]},
      {stage2_52[85], stage2_52[86], stage2_52[87], stage2_52[88], stage2_52[89], stage2_52[90]},
      {stage3_54[16],stage3_53[27],stage3_52[31],stage3_51[41],stage3_50[56]}
   );
   gpc606_5 gpc9041 (
      {stage2_50[131], stage2_50[132], stage2_50[133], stage2_50[134], stage2_50[135], stage2_50[136]},
      {stage2_52[91], stage2_52[92], stage2_52[93], stage2_52[94], stage2_52[95], stage2_52[96]},
      {stage3_54[17],stage3_53[28],stage3_52[32],stage3_51[42],stage3_50[57]}
   );
   gpc606_5 gpc9042 (
      {stage2_50[137], stage2_50[138], stage2_50[139], stage2_50[140], stage2_50[141], stage2_50[142]},
      {stage2_52[97], stage2_52[98], stage2_52[99], stage2_52[100], stage2_52[101], stage2_52[102]},
      {stage3_54[18],stage3_53[29],stage3_52[33],stage3_51[43],stage3_50[58]}
   );
   gpc606_5 gpc9043 (
      {stage2_50[143], stage2_50[144], stage2_50[145], stage2_50[146], stage2_50[147], stage2_50[148]},
      {stage2_52[103], stage2_52[104], stage2_52[105], stage2_52[106], stage2_52[107], stage2_52[108]},
      {stage3_54[19],stage3_53[30],stage3_52[34],stage3_51[44],stage3_50[59]}
   );
   gpc606_5 gpc9044 (
      {stage2_51[69], stage2_51[70], stage2_51[71], stage2_51[72], stage2_51[73], stage2_51[74]},
      {stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10]},
      {stage3_55[0],stage3_54[20],stage3_53[31],stage3_52[35],stage3_51[45]}
   );
   gpc606_5 gpc9045 (
      {stage2_51[75], stage2_51[76], stage2_51[77], stage2_51[78], stage2_51[79], stage2_51[80]},
      {stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16]},
      {stage3_55[1],stage3_54[21],stage3_53[32],stage3_52[36],stage3_51[46]}
   );
   gpc606_5 gpc9046 (
      {stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[2],stage3_54[22],stage3_53[33]}
   );
   gpc606_5 gpc9047 (
      {stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[3],stage3_54[23],stage3_53[34]}
   );
   gpc606_5 gpc9048 (
      {stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[4],stage3_54[24],stage3_53[35]}
   );
   gpc606_5 gpc9049 (
      {stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[3],stage3_55[5],stage3_54[25],stage3_53[36]}
   );
   gpc606_5 gpc9050 (
      {stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[4],stage3_55[6],stage3_54[26],stage3_53[37]}
   );
   gpc606_5 gpc9051 (
      {stage2_53[47], stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[5],stage3_55[7],stage3_54[27],stage3_53[38]}
   );
   gpc606_5 gpc9052 (
      {stage2_53[53], stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[6],stage3_55[8],stage3_54[28],stage3_53[39]}
   );
   gpc606_5 gpc9053 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63], stage2_53[64]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[7],stage3_55[9],stage3_54[29],stage3_53[40]}
   );
   gpc606_5 gpc9054 (
      {stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68], stage2_53[69], stage2_53[70]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[8],stage3_55[10],stage3_54[30],stage3_53[41]}
   );
   gpc606_5 gpc9055 (
      {stage2_53[71], stage2_53[72], stage2_53[73], stage2_53[74], stage2_53[75], stage2_53[76]},
      {stage2_55[54], stage2_55[55], stage2_55[56], stage2_55[57], stage2_55[58], stage2_55[59]},
      {stage3_57[9],stage3_56[9],stage3_55[11],stage3_54[31],stage3_53[42]}
   );
   gpc606_5 gpc9056 (
      {stage2_53[77], stage2_53[78], stage2_53[79], stage2_53[80], stage2_53[81], stage2_53[82]},
      {stage2_55[60], stage2_55[61], stage2_55[62], stage2_55[63], stage2_55[64], stage2_55[65]},
      {stage3_57[10],stage3_56[10],stage3_55[12],stage3_54[32],stage3_53[43]}
   );
   gpc606_5 gpc9057 (
      {stage2_53[83], stage2_53[84], stage2_53[85], stage2_53[86], stage2_53[87], stage2_53[88]},
      {stage2_55[66], stage2_55[67], stage2_55[68], stage2_55[69], stage2_55[70], stage2_55[71]},
      {stage3_57[11],stage3_56[11],stage3_55[13],stage3_54[33],stage3_53[44]}
   );
   gpc606_5 gpc9058 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[12],stage3_56[12],stage3_55[14],stage3_54[34]}
   );
   gpc606_5 gpc9059 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[13],stage3_56[13],stage3_55[15],stage3_54[35]}
   );
   gpc606_5 gpc9060 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[14],stage3_56[14],stage3_55[16],stage3_54[36]}
   );
   gpc606_5 gpc9061 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22], stage2_54[23]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[15],stage3_56[15],stage3_55[17],stage3_54[37]}
   );
   gpc606_5 gpc9062 (
      {stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[16],stage3_56[16],stage3_55[18],stage3_54[38]}
   );
   gpc606_5 gpc9063 (
      {stage2_54[30], stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[17],stage3_56[17],stage3_55[19],stage3_54[39]}
   );
   gpc606_5 gpc9064 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40], stage2_54[41]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[18],stage3_56[18],stage3_55[20],stage3_54[40]}
   );
   gpc606_5 gpc9065 (
      {stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45], stage2_54[46], stage2_54[47]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[19],stage3_56[19],stage3_55[21],stage3_54[41]}
   );
   gpc606_5 gpc9066 (
      {stage2_54[48], stage2_54[49], stage2_54[50], stage2_54[51], stage2_54[52], stage2_54[53]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[20],stage3_56[20],stage3_55[22],stage3_54[42]}
   );
   gpc606_5 gpc9067 (
      {stage2_54[54], stage2_54[55], stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[21],stage3_56[21],stage3_55[23],stage3_54[43]}
   );
   gpc606_5 gpc9068 (
      {stage2_54[60], stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[22],stage3_56[22],stage3_55[24],stage3_54[44]}
   );
   gpc606_5 gpc9069 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70], stage2_54[71]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[23],stage3_56[23],stage3_55[25],stage3_54[45]}
   );
   gpc606_5 gpc9070 (
      {stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75], stage2_54[76], stage2_54[77]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[24],stage3_56[24],stage3_55[26],stage3_54[46]}
   );
   gpc606_5 gpc9071 (
      {stage2_54[78], stage2_54[79], stage2_54[80], stage2_54[81], stage2_54[82], stage2_54[83]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[25],stage3_56[25],stage3_55[27],stage3_54[47]}
   );
   gpc606_5 gpc9072 (
      {stage2_54[84], stage2_54[85], stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[26],stage3_56[26],stage3_55[28],stage3_54[48]}
   );
   gpc606_5 gpc9073 (
      {stage2_54[90], stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[27],stage3_56[27],stage3_55[29],stage3_54[49]}
   );
   gpc606_5 gpc9074 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], stage2_54[100], stage2_54[101]},
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100], stage2_56[101]},
      {stage3_58[16],stage3_57[28],stage3_56[28],stage3_55[30],stage3_54[50]}
   );
   gpc606_5 gpc9075 (
      {stage2_54[102], stage2_54[103], stage2_54[104], stage2_54[105], stage2_54[106], stage2_54[107]},
      {stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105], stage2_56[106], stage2_56[107]},
      {stage3_58[17],stage3_57[29],stage3_56[29],stage3_55[31],stage3_54[51]}
   );
   gpc606_5 gpc9076 (
      {stage2_54[108], stage2_54[109], stage2_54[110], stage2_54[111], stage2_54[112], stage2_54[113]},
      {stage2_56[108], stage2_56[109], stage2_56[110], stage2_56[111], stage2_56[112], stage2_56[113]},
      {stage3_58[18],stage3_57[30],stage3_56[30],stage3_55[32],stage3_54[52]}
   );
   gpc606_5 gpc9077 (
      {stage2_55[72], stage2_55[73], stage2_55[74], stage2_55[75], stage2_55[76], stage2_55[77]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[19],stage3_57[31],stage3_56[31],stage3_55[33]}
   );
   gpc606_5 gpc9078 (
      {stage2_55[78], stage2_55[79], stage2_55[80], stage2_55[81], stage2_55[82], stage2_55[83]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[20],stage3_57[32],stage3_56[32],stage3_55[34]}
   );
   gpc606_5 gpc9079 (
      {stage2_55[84], stage2_55[85], stage2_55[86], stage2_55[87], stage2_55[88], stage2_55[89]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[21],stage3_57[33],stage3_56[33],stage3_55[35]}
   );
   gpc606_5 gpc9080 (
      {stage2_55[90], stage2_55[91], stage2_55[92], stage2_55[93], stage2_55[94], stage2_55[95]},
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage3_59[3],stage3_58[22],stage3_57[34],stage3_56[34],stage3_55[36]}
   );
   gpc606_5 gpc9081 (
      {stage2_55[96], stage2_55[97], stage2_55[98], stage2_55[99], stage2_55[100], stage2_55[101]},
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage3_59[4],stage3_58[23],stage3_57[35],stage3_56[35],stage3_55[37]}
   );
   gpc606_5 gpc9082 (
      {stage2_56[114], stage2_56[115], stage2_56[116], stage2_56[117], stage2_56[118], stage2_56[119]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[5],stage3_58[24],stage3_57[36],stage3_56[36]}
   );
   gpc606_5 gpc9083 (
      {stage2_56[120], stage2_56[121], stage2_56[122], stage2_56[123], stage2_56[124], stage2_56[125]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[6],stage3_58[25],stage3_57[37],stage3_56[37]}
   );
   gpc606_5 gpc9084 (
      {stage2_56[126], stage2_56[127], stage2_56[128], stage2_56[129], stage2_56[130], stage2_56[131]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[7],stage3_58[26],stage3_57[38],stage3_56[38]}
   );
   gpc606_5 gpc9085 (
      {stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33], stage2_57[34], stage2_57[35]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[3],stage3_59[8],stage3_58[27],stage3_57[39]}
   );
   gpc606_5 gpc9086 (
      {stage2_57[36], stage2_57[37], stage2_57[38], stage2_57[39], stage2_57[40], stage2_57[41]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[4],stage3_59[9],stage3_58[28],stage3_57[40]}
   );
   gpc606_5 gpc9087 (
      {stage2_57[42], stage2_57[43], stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[5],stage3_59[10],stage3_58[29],stage3_57[41]}
   );
   gpc606_5 gpc9088 (
      {stage2_57[48], stage2_57[49], stage2_57[50], stage2_57[51], stage2_57[52], stage2_57[53]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[6],stage3_59[11],stage3_58[30],stage3_57[42]}
   );
   gpc606_5 gpc9089 (
      {stage2_57[54], stage2_57[55], stage2_57[56], stage2_57[57], stage2_57[58], stage2_57[59]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[7],stage3_59[12],stage3_58[31],stage3_57[43]}
   );
   gpc606_5 gpc9090 (
      {stage2_57[60], stage2_57[61], stage2_57[62], stage2_57[63], stage2_57[64], stage2_57[65]},
      {stage2_59[30], stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35]},
      {stage3_61[5],stage3_60[8],stage3_59[13],stage3_58[32],stage3_57[44]}
   );
   gpc606_5 gpc9091 (
      {stage2_57[66], stage2_57[67], stage2_57[68], stage2_57[69], stage2_57[70], stage2_57[71]},
      {stage2_59[36], stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41]},
      {stage3_61[6],stage3_60[9],stage3_59[14],stage3_58[33],stage3_57[45]}
   );
   gpc207_4 gpc9092 (
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23], stage2_58[24]},
      {stage2_60[0], stage2_60[1]},
      {stage3_61[7],stage3_60[10],stage3_59[15],stage3_58[34]}
   );
   gpc207_4 gpc9093 (
      {stage2_58[25], stage2_58[26], stage2_58[27], stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31]},
      {stage2_60[2], stage2_60[3]},
      {stage3_61[8],stage3_60[11],stage3_59[16],stage3_58[35]}
   );
   gpc207_4 gpc9094 (
      {stage2_58[32], stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37], stage2_58[38]},
      {stage2_60[4], stage2_60[5]},
      {stage3_61[9],stage3_60[12],stage3_59[17],stage3_58[36]}
   );
   gpc207_4 gpc9095 (
      {stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42], stage2_58[43], stage2_58[44], stage2_58[45]},
      {stage2_60[6], stage2_60[7]},
      {stage3_61[10],stage3_60[13],stage3_59[18],stage3_58[37]}
   );
   gpc207_4 gpc9096 (
      {stage2_58[46], stage2_58[47], stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_60[8], stage2_60[9]},
      {stage3_61[11],stage3_60[14],stage3_59[19],stage3_58[38]}
   );
   gpc207_4 gpc9097 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57], stage2_58[58], stage2_58[59]},
      {stage2_60[10], stage2_60[11]},
      {stage3_61[12],stage3_60[15],stage3_59[20],stage3_58[39]}
   );
   gpc207_4 gpc9098 (
      {stage2_58[60], stage2_58[61], stage2_58[62], stage2_58[63], stage2_58[64], stage2_58[65], stage2_58[66]},
      {stage2_60[12], stage2_60[13]},
      {stage3_61[13],stage3_60[16],stage3_59[21],stage3_58[40]}
   );
   gpc207_4 gpc9099 (
      {stage2_58[67], stage2_58[68], stage2_58[69], stage2_58[70], stage2_58[71], stage2_58[72], stage2_58[73]},
      {stage2_60[14], stage2_60[15]},
      {stage3_61[14],stage3_60[17],stage3_59[22],stage3_58[41]}
   );
   gpc615_5 gpc9100 (
      {stage2_58[74], stage2_58[75], stage2_58[76], stage2_58[77], stage2_58[78]},
      {stage2_59[42]},
      {stage2_60[16], stage2_60[17], stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21]},
      {stage3_62[0],stage3_61[15],stage3_60[18],stage3_59[23],stage3_58[42]}
   );
   gpc606_5 gpc9101 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[1],stage3_61[16],stage3_60[19],stage3_59[24]}
   );
   gpc606_5 gpc9102 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[2],stage3_61[17],stage3_60[20],stage3_59[25]}
   );
   gpc606_5 gpc9103 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59], stage2_59[60]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[3],stage3_61[18],stage3_60[21],stage3_59[26]}
   );
   gpc606_5 gpc9104 (
      {stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64], stage2_59[65], stage2_59[66]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[4],stage3_61[19],stage3_60[22],stage3_59[27]}
   );
   gpc606_5 gpc9105 (
      {stage2_59[67], stage2_59[68], stage2_59[69], stage2_59[70], stage2_59[71], stage2_59[72]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[5],stage3_61[20],stage3_60[23],stage3_59[28]}
   );
   gpc606_5 gpc9106 (
      {stage2_59[73], stage2_59[74], stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[6],stage3_61[21],stage3_60[24],stage3_59[29]}
   );
   gpc606_5 gpc9107 (
      {stage2_59[79], stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[7],stage3_61[22],stage3_60[25],stage3_59[30]}
   );
   gpc606_5 gpc9108 (
      {stage2_59[85], stage2_59[86], stage2_59[87], stage2_59[88], stage2_59[89], stage2_59[90]},
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage3_63[7],stage3_62[8],stage3_61[23],stage3_60[26],stage3_59[31]}
   );
   gpc606_5 gpc9109 (
      {stage2_59[91], stage2_59[92], stage2_59[93], stage2_59[94], stage2_59[95], stage2_59[96]},
      {stage2_61[48], stage2_61[49], stage2_61[50], stage2_61[51], stage2_61[52], stage2_61[53]},
      {stage3_63[8],stage3_62[9],stage3_61[24],stage3_60[27],stage3_59[32]}
   );
   gpc606_5 gpc9110 (
      {stage2_59[97], stage2_59[98], stage2_59[99], stage2_59[100], stage2_59[101], stage2_59[102]},
      {stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58], stage2_61[59]},
      {stage3_63[9],stage3_62[10],stage3_61[25],stage3_60[28],stage3_59[33]}
   );
   gpc606_5 gpc9111 (
      {stage2_59[103], stage2_59[104], stage2_59[105], stage2_59[106], stage2_59[107], stage2_59[108]},
      {stage2_61[60], stage2_61[61], stage2_61[62], stage2_61[63], stage2_61[64], stage2_61[65]},
      {stage3_63[10],stage3_62[11],stage3_61[26],stage3_60[29],stage3_59[34]}
   );
   gpc606_5 gpc9112 (
      {stage2_59[109], stage2_59[110], stage2_59[111], stage2_59[112], stage2_59[113], stage2_59[114]},
      {stage2_61[66], stage2_61[67], stage2_61[68], stage2_61[69], stage2_61[70], stage2_61[71]},
      {stage3_63[11],stage3_62[12],stage3_61[27],stage3_60[30],stage3_59[35]}
   );
   gpc606_5 gpc9113 (
      {stage2_59[115], stage2_59[116], stage2_59[117], stage2_59[118], stage2_59[119], stage2_59[120]},
      {stage2_61[72], stage2_61[73], stage2_61[74], stage2_61[75], stage2_61[76], stage2_61[77]},
      {stage3_63[12],stage3_62[13],stage3_61[28],stage3_60[31],stage3_59[36]}
   );
   gpc606_5 gpc9114 (
      {stage2_59[121], stage2_59[122], stage2_59[123], stage2_59[124], stage2_59[125], stage2_59[126]},
      {stage2_61[78], stage2_61[79], stage2_61[80], stage2_61[81], stage2_61[82], stage2_61[83]},
      {stage3_63[13],stage3_62[14],stage3_61[29],stage3_60[32],stage3_59[37]}
   );
   gpc606_5 gpc9115 (
      {stage2_59[127], stage2_59[128], stage2_59[129], stage2_59[130], stage2_59[131], stage2_59[132]},
      {stage2_61[84], stage2_61[85], stage2_61[86], stage2_61[87], stage2_61[88], stage2_61[89]},
      {stage3_63[14],stage3_62[15],stage3_61[30],stage3_60[33],stage3_59[38]}
   );
   gpc606_5 gpc9116 (
      {stage2_60[22], stage2_60[23], stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[15],stage3_62[16],stage3_61[31],stage3_60[34]}
   );
   gpc606_5 gpc9117 (
      {stage2_60[28], stage2_60[29], stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[16],stage3_62[17],stage3_61[32],stage3_60[35]}
   );
   gpc606_5 gpc9118 (
      {stage2_60[34], stage2_60[35], stage2_60[36], stage2_60[37], stage2_60[38], stage2_60[39]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[17],stage3_62[18],stage3_61[33],stage3_60[36]}
   );
   gpc606_5 gpc9119 (
      {stage2_60[40], stage2_60[41], stage2_60[42], stage2_60[43], stage2_60[44], stage2_60[45]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[18],stage3_62[19],stage3_61[34],stage3_60[37]}
   );
   gpc606_5 gpc9120 (
      {stage2_60[46], stage2_60[47], stage2_60[48], stage2_60[49], stage2_60[50], stage2_60[51]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[19],stage3_62[20],stage3_61[35],stage3_60[38]}
   );
   gpc606_5 gpc9121 (
      {stage2_60[52], stage2_60[53], stage2_60[54], stage2_60[55], stage2_60[56], stage2_60[57]},
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34], stage2_62[35]},
      {stage3_64[5],stage3_63[20],stage3_62[21],stage3_61[36],stage3_60[39]}
   );
   gpc606_5 gpc9122 (
      {stage2_60[58], stage2_60[59], stage2_60[60], stage2_60[61], stage2_60[62], stage2_60[63]},
      {stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39], stage2_62[40], stage2_62[41]},
      {stage3_64[6],stage3_63[21],stage3_62[22],stage3_61[37],stage3_60[40]}
   );
   gpc606_5 gpc9123 (
      {stage2_60[64], stage2_60[65], stage2_60[66], stage2_60[67], stage2_60[68], stage2_60[69]},
      {stage2_62[42], stage2_62[43], stage2_62[44], stage2_62[45], stage2_62[46], stage2_62[47]},
      {stage3_64[7],stage3_63[22],stage3_62[23],stage3_61[38],stage3_60[41]}
   );
   gpc606_5 gpc9124 (
      {stage2_60[70], stage2_60[71], stage2_60[72], stage2_60[73], stage2_60[74], stage2_60[75]},
      {stage2_62[48], stage2_62[49], stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53]},
      {stage3_64[8],stage3_63[23],stage3_62[24],stage3_61[39],stage3_60[42]}
   );
   gpc606_5 gpc9125 (
      {stage2_60[76], stage2_60[77], stage2_60[78], stage2_60[79], stage2_60[80], stage2_60[81]},
      {stage2_62[54], stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage3_64[9],stage3_63[24],stage3_62[25],stage3_61[40],stage3_60[43]}
   );
   gpc606_5 gpc9126 (
      {stage2_60[82], stage2_60[83], stage2_60[84], stage2_60[85], stage2_60[86], stage2_60[87]},
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64], stage2_62[65]},
      {stage3_64[10],stage3_63[25],stage3_62[26],stage3_61[41],stage3_60[44]}
   );
   gpc606_5 gpc9127 (
      {stage2_60[88], stage2_60[89], stage2_60[90], stage2_60[91], stage2_60[92], stage2_60[93]},
      {stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69], stage2_62[70], stage2_62[71]},
      {stage3_64[11],stage3_63[26],stage3_62[27],stage3_61[42],stage3_60[45]}
   );
   gpc606_5 gpc9128 (
      {stage2_60[94], stage2_60[95], stage2_60[96], stage2_60[97], stage2_60[98], stage2_60[99]},
      {stage2_62[72], stage2_62[73], stage2_62[74], stage2_62[75], stage2_62[76], stage2_62[77]},
      {stage3_64[12],stage3_63[27],stage3_62[28],stage3_61[43],stage3_60[46]}
   );
   gpc606_5 gpc9129 (
      {stage2_60[100], stage2_60[101], stage2_60[102], stage2_60[103], stage2_60[104], stage2_60[105]},
      {stage2_62[78], stage2_62[79], stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83]},
      {stage3_64[13],stage3_63[28],stage3_62[29],stage3_61[44],stage3_60[47]}
   );
   gpc606_5 gpc9130 (
      {stage2_62[84], stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[0],stage3_64[14],stage3_63[29],stage3_62[30]}
   );
   gpc606_5 gpc9131 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94], stage2_62[95]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[1],stage3_64[15],stage3_63[30],stage3_62[31]}
   );
   gpc606_5 gpc9132 (
      {stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99], stage2_62[100], stage2_62[101]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[2],stage3_64[16],stage3_63[31],stage3_62[32]}
   );
   gpc606_5 gpc9133 (
      {stage2_62[102], stage2_62[103], stage2_62[104], stage2_62[105], stage2_62[106], stage2_62[107]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[3],stage3_64[17],stage3_63[32],stage3_62[33]}
   );
   gpc606_5 gpc9134 (
      {stage2_62[108], stage2_62[109], stage2_62[110], stage2_62[111], stage2_62[112], stage2_62[113]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[4],stage3_64[18],stage3_63[33],stage3_62[34]}
   );
   gpc606_5 gpc9135 (
      {stage2_62[114], stage2_62[115], stage2_62[116], stage2_62[117], stage2_62[118], stage2_62[119]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[5],stage3_64[19],stage3_63[34],stage3_62[35]}
   );
   gpc606_5 gpc9136 (
      {stage2_62[120], stage2_62[121], stage2_62[122], stage2_62[123], stage2_62[124], stage2_62[125]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[6],stage3_64[20],stage3_63[35],stage3_62[36]}
   );
   gpc606_5 gpc9137 (
      {stage2_62[126], stage2_62[127], stage2_62[128], stage2_62[129], stage2_62[130], stage2_62[131]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[7],stage3_64[21],stage3_63[36],stage3_62[37]}
   );
   gpc606_5 gpc9138 (
      {stage2_62[132], stage2_62[133], stage2_62[134], stage2_62[135], stage2_62[136], stage2_62[137]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[8],stage3_64[22],stage3_63[37],stage3_62[38]}
   );
   gpc606_5 gpc9139 (
      {stage2_62[138], stage2_62[139], stage2_62[140], stage2_62[141], stage2_62[142], stage2_62[143]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[9],stage3_64[23],stage3_63[38],stage3_62[39]}
   );
   gpc117_4 gpc9140 (
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage2_64[60]},
      {stage2_65[0]},
      {stage3_66[10],stage3_65[10],stage3_64[24],stage3_63[39]}
   );
   gpc117_4 gpc9141 (
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12], stage2_63[13]},
      {stage2_64[61]},
      {stage2_65[1]},
      {stage3_66[11],stage3_65[11],stage3_64[25],stage3_63[40]}
   );
   gpc117_4 gpc9142 (
      {stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18], stage2_63[19], stage2_63[20]},
      {stage2_64[62]},
      {stage2_65[2]},
      {stage3_66[12],stage3_65[12],stage3_64[26],stage3_63[41]}
   );
   gpc117_4 gpc9143 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[63]},
      {stage2_65[3]},
      {stage3_66[13],stage3_65[13],stage3_64[27],stage3_63[42]}
   );
   gpc117_4 gpc9144 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[64]},
      {stage2_65[4]},
      {stage3_66[14],stage3_65[14],stage3_64[28],stage3_63[43]}
   );
   gpc606_5 gpc9145 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40]},
      {stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9], stage2_65[10]},
      {stage3_67[0],stage3_66[15],stage3_65[15],stage3_64[29],stage3_63[44]}
   );
   gpc606_5 gpc9146 (
      {stage2_63[41], stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46]},
      {stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14], stage2_65[15], stage2_65[16]},
      {stage3_67[1],stage3_66[16],stage3_65[16],stage3_64[30],stage3_63[45]}
   );
   gpc606_5 gpc9147 (
      {stage2_63[47], stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52]},
      {stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20], stage2_65[21], stage2_65[22]},
      {stage3_67[2],stage3_66[17],stage3_65[17],stage3_64[31],stage3_63[46]}
   );
   gpc606_5 gpc9148 (
      {stage2_63[53], stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58]},
      {stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26], stage2_65[27], stage2_65[28]},
      {stage3_67[3],stage3_66[18],stage3_65[18],stage3_64[32],stage3_63[47]}
   );
   gpc606_5 gpc9149 (
      {stage2_63[59], stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64]},
      {stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32], stage2_65[33], stage2_65[34]},
      {stage3_67[4],stage3_66[19],stage3_65[19],stage3_64[33],stage3_63[48]}
   );
   gpc606_5 gpc9150 (
      {stage2_63[65], stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70]},
      {stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38], stage2_65[39], stage2_65[40]},
      {stage3_67[5],stage3_66[20],stage3_65[20],stage3_64[34],stage3_63[49]}
   );
   gpc606_5 gpc9151 (
      {stage2_63[71], stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76]},
      {stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44], stage2_65[45], stage2_65[46]},
      {stage3_67[6],stage3_66[21],stage3_65[21],stage3_64[35],stage3_63[50]}
   );
   gpc606_5 gpc9152 (
      {stage2_63[77], stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82]},
      {stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50], stage2_65[51], stage2_65[52]},
      {stage3_67[7],stage3_66[22],stage3_65[22],stage3_64[36],stage3_63[51]}
   );
   gpc606_5 gpc9153 (
      {stage2_63[83], stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88]},
      {stage2_65[53], stage2_65[54], stage2_65[55], stage2_65[56], stage2_65[57], stage2_65[58]},
      {stage3_67[8],stage3_66[23],stage3_65[23],stage3_64[37],stage3_63[52]}
   );
   gpc606_5 gpc9154 (
      {stage2_63[89], stage2_63[90], stage2_63[91], stage2_63[92], stage2_63[93], stage2_63[94]},
      {stage2_65[59], stage2_65[60], stage2_65[61], stage2_65[62], stage2_65[63], stage2_65[64]},
      {stage3_67[9],stage3_66[24],stage3_65[24],stage3_64[38],stage3_63[53]}
   );
   gpc606_5 gpc9155 (
      {stage2_64[65], stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[10],stage3_66[25],stage3_65[25],stage3_64[39]}
   );
   gpc606_5 gpc9156 (
      {stage2_64[71], stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[11],stage3_66[26],stage3_65[26],stage3_64[40]}
   );
   gpc606_5 gpc9157 (
      {stage2_64[77], stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[12],stage3_66[27],stage3_65[27],stage3_64[41]}
   );
   gpc606_5 gpc9158 (
      {stage2_64[83], stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[13],stage3_66[28],stage3_65[28],stage3_64[42]}
   );
   gpc606_5 gpc9159 (
      {stage2_64[89], stage2_64[90], stage2_64[91], stage2_64[92], stage2_64[93], stage2_64[94]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[14],stage3_66[29],stage3_65[29],stage3_64[43]}
   );
   gpc1_1 gpc9160 (
      {stage2_0[29]},
      {stage3_0[6]}
   );
   gpc1_1 gpc9161 (
      {stage2_0[30]},
      {stage3_0[7]}
   );
   gpc1_1 gpc9162 (
      {stage2_0[31]},
      {stage3_0[8]}
   );
   gpc1_1 gpc9163 (
      {stage2_0[32]},
      {stage3_0[9]}
   );
   gpc1_1 gpc9164 (
      {stage2_0[33]},
      {stage3_0[10]}
   );
   gpc1_1 gpc9165 (
      {stage2_1[22]},
      {stage3_1[9]}
   );
   gpc1_1 gpc9166 (
      {stage2_1[23]},
      {stage3_1[10]}
   );
   gpc1_1 gpc9167 (
      {stage2_1[24]},
      {stage3_1[11]}
   );
   gpc1_1 gpc9168 (
      {stage2_1[25]},
      {stage3_1[12]}
   );
   gpc1_1 gpc9169 (
      {stage2_1[26]},
      {stage3_1[13]}
   );
   gpc1_1 gpc9170 (
      {stage2_1[27]},
      {stage3_1[14]}
   );
   gpc1_1 gpc9171 (
      {stage2_1[28]},
      {stage3_1[15]}
   );
   gpc1_1 gpc9172 (
      {stage2_1[29]},
      {stage3_1[16]}
   );
   gpc1_1 gpc9173 (
      {stage2_1[30]},
      {stage3_1[17]}
   );
   gpc1_1 gpc9174 (
      {stage2_1[31]},
      {stage3_1[18]}
   );
   gpc1_1 gpc9175 (
      {stage2_1[32]},
      {stage3_1[19]}
   );
   gpc1_1 gpc9176 (
      {stage2_1[33]},
      {stage3_1[20]}
   );
   gpc1_1 gpc9177 (
      {stage2_1[34]},
      {stage3_1[21]}
   );
   gpc1_1 gpc9178 (
      {stage2_1[35]},
      {stage3_1[22]}
   );
   gpc1_1 gpc9179 (
      {stage2_1[36]},
      {stage3_1[23]}
   );
   gpc1_1 gpc9180 (
      {stage2_1[37]},
      {stage3_1[24]}
   );
   gpc1_1 gpc9181 (
      {stage2_1[38]},
      {stage3_1[25]}
   );
   gpc1_1 gpc9182 (
      {stage2_7[85]},
      {stage3_7[43]}
   );
   gpc1_1 gpc9183 (
      {stage2_7[86]},
      {stage3_7[44]}
   );
   gpc1_1 gpc9184 (
      {stage2_7[87]},
      {stage3_7[45]}
   );
   gpc1_1 gpc9185 (
      {stage2_7[88]},
      {stage3_7[46]}
   );
   gpc1_1 gpc9186 (
      {stage2_7[89]},
      {stage3_7[47]}
   );
   gpc1_1 gpc9187 (
      {stage2_7[90]},
      {stage3_7[48]}
   );
   gpc1_1 gpc9188 (
      {stage2_7[91]},
      {stage3_7[49]}
   );
   gpc1_1 gpc9189 (
      {stage2_7[92]},
      {stage3_7[50]}
   );
   gpc1_1 gpc9190 (
      {stage2_7[93]},
      {stage3_7[51]}
   );
   gpc1_1 gpc9191 (
      {stage2_7[94]},
      {stage3_7[52]}
   );
   gpc1_1 gpc9192 (
      {stage2_7[95]},
      {stage3_7[53]}
   );
   gpc1_1 gpc9193 (
      {stage2_7[96]},
      {stage3_7[54]}
   );
   gpc1_1 gpc9194 (
      {stage2_10[125]},
      {stage3_10[59]}
   );
   gpc1_1 gpc9195 (
      {stage2_10[126]},
      {stage3_10[60]}
   );
   gpc1_1 gpc9196 (
      {stage2_10[127]},
      {stage3_10[61]}
   );
   gpc1_1 gpc9197 (
      {stage2_10[128]},
      {stage3_10[62]}
   );
   gpc1_1 gpc9198 (
      {stage2_10[129]},
      {stage3_10[63]}
   );
   gpc1_1 gpc9199 (
      {stage2_10[130]},
      {stage3_10[64]}
   );
   gpc1_1 gpc9200 (
      {stage2_10[131]},
      {stage3_10[65]}
   );
   gpc1_1 gpc9201 (
      {stage2_10[132]},
      {stage3_10[66]}
   );
   gpc1_1 gpc9202 (
      {stage2_10[133]},
      {stage3_10[67]}
   );
   gpc1_1 gpc9203 (
      {stage2_11[125]},
      {stage3_11[50]}
   );
   gpc1_1 gpc9204 (
      {stage2_11[126]},
      {stage3_11[51]}
   );
   gpc1_1 gpc9205 (
      {stage2_11[127]},
      {stage3_11[52]}
   );
   gpc1_1 gpc9206 (
      {stage2_11[128]},
      {stage3_11[53]}
   );
   gpc1_1 gpc9207 (
      {stage2_11[129]},
      {stage3_11[54]}
   );
   gpc1_1 gpc9208 (
      {stage2_11[130]},
      {stage3_11[55]}
   );
   gpc1_1 gpc9209 (
      {stage2_11[131]},
      {stage3_11[56]}
   );
   gpc1_1 gpc9210 (
      {stage2_11[132]},
      {stage3_11[57]}
   );
   gpc1_1 gpc9211 (
      {stage2_11[133]},
      {stage3_11[58]}
   );
   gpc1_1 gpc9212 (
      {stage2_11[134]},
      {stage3_11[59]}
   );
   gpc1_1 gpc9213 (
      {stage2_11[135]},
      {stage3_11[60]}
   );
   gpc1_1 gpc9214 (
      {stage2_12[98]},
      {stage3_12[51]}
   );
   gpc1_1 gpc9215 (
      {stage2_12[99]},
      {stage3_12[52]}
   );
   gpc1_1 gpc9216 (
      {stage2_12[100]},
      {stage3_12[53]}
   );
   gpc1_1 gpc9217 (
      {stage2_12[101]},
      {stage3_12[54]}
   );
   gpc1_1 gpc9218 (
      {stage2_12[102]},
      {stage3_12[55]}
   );
   gpc1_1 gpc9219 (
      {stage2_12[103]},
      {stage3_12[56]}
   );
   gpc1_1 gpc9220 (
      {stage2_12[104]},
      {stage3_12[57]}
   );
   gpc1_1 gpc9221 (
      {stage2_12[105]},
      {stage3_12[58]}
   );
   gpc1_1 gpc9222 (
      {stage2_12[106]},
      {stage3_12[59]}
   );
   gpc1_1 gpc9223 (
      {stage2_12[107]},
      {stage3_12[60]}
   );
   gpc1_1 gpc9224 (
      {stage2_12[108]},
      {stage3_12[61]}
   );
   gpc1_1 gpc9225 (
      {stage2_12[109]},
      {stage3_12[62]}
   );
   gpc1_1 gpc9226 (
      {stage2_12[110]},
      {stage3_12[63]}
   );
   gpc1_1 gpc9227 (
      {stage2_12[111]},
      {stage3_12[64]}
   );
   gpc1_1 gpc9228 (
      {stage2_12[112]},
      {stage3_12[65]}
   );
   gpc1_1 gpc9229 (
      {stage2_12[113]},
      {stage3_12[66]}
   );
   gpc1_1 gpc9230 (
      {stage2_12[114]},
      {stage3_12[67]}
   );
   gpc1_1 gpc9231 (
      {stage2_12[115]},
      {stage3_12[68]}
   );
   gpc1_1 gpc9232 (
      {stage2_12[116]},
      {stage3_12[69]}
   );
   gpc1_1 gpc9233 (
      {stage2_12[117]},
      {stage3_12[70]}
   );
   gpc1_1 gpc9234 (
      {stage2_12[118]},
      {stage3_12[71]}
   );
   gpc1_1 gpc9235 (
      {stage2_12[119]},
      {stage3_12[72]}
   );
   gpc1_1 gpc9236 (
      {stage2_12[120]},
      {stage3_12[73]}
   );
   gpc1_1 gpc9237 (
      {stage2_12[121]},
      {stage3_12[74]}
   );
   gpc1_1 gpc9238 (
      {stage2_12[122]},
      {stage3_12[75]}
   );
   gpc1_1 gpc9239 (
      {stage2_12[123]},
      {stage3_12[76]}
   );
   gpc1_1 gpc9240 (
      {stage2_12[124]},
      {stage3_12[77]}
   );
   gpc1_1 gpc9241 (
      {stage2_12[125]},
      {stage3_12[78]}
   );
   gpc1_1 gpc9242 (
      {stage2_12[126]},
      {stage3_12[79]}
   );
   gpc1_1 gpc9243 (
      {stage2_12[127]},
      {stage3_12[80]}
   );
   gpc1_1 gpc9244 (
      {stage2_13[70]},
      {stage3_13[45]}
   );
   gpc1_1 gpc9245 (
      {stage2_13[71]},
      {stage3_13[46]}
   );
   gpc1_1 gpc9246 (
      {stage2_15[108]},
      {stage3_15[44]}
   );
   gpc1_1 gpc9247 (
      {stage2_15[109]},
      {stage3_15[45]}
   );
   gpc1_1 gpc9248 (
      {stage2_15[110]},
      {stage3_15[46]}
   );
   gpc1_1 gpc9249 (
      {stage2_15[111]},
      {stage3_15[47]}
   );
   gpc1_1 gpc9250 (
      {stage2_15[112]},
      {stage3_15[48]}
   );
   gpc1_1 gpc9251 (
      {stage2_15[113]},
      {stage3_15[49]}
   );
   gpc1_1 gpc9252 (
      {stage2_15[114]},
      {stage3_15[50]}
   );
   gpc1_1 gpc9253 (
      {stage2_16[96]},
      {stage3_16[45]}
   );
   gpc1_1 gpc9254 (
      {stage2_16[97]},
      {stage3_16[46]}
   );
   gpc1_1 gpc9255 (
      {stage2_16[98]},
      {stage3_16[47]}
   );
   gpc1_1 gpc9256 (
      {stage2_16[99]},
      {stage3_16[48]}
   );
   gpc1_1 gpc9257 (
      {stage2_16[100]},
      {stage3_16[49]}
   );
   gpc1_1 gpc9258 (
      {stage2_16[101]},
      {stage3_16[50]}
   );
   gpc1_1 gpc9259 (
      {stage2_16[102]},
      {stage3_16[51]}
   );
   gpc1_1 gpc9260 (
      {stage2_16[103]},
      {stage3_16[52]}
   );
   gpc1_1 gpc9261 (
      {stage2_16[104]},
      {stage3_16[53]}
   );
   gpc1_1 gpc9262 (
      {stage2_16[105]},
      {stage3_16[54]}
   );
   gpc1_1 gpc9263 (
      {stage2_16[106]},
      {stage3_16[55]}
   );
   gpc1_1 gpc9264 (
      {stage2_16[107]},
      {stage3_16[56]}
   );
   gpc1_1 gpc9265 (
      {stage2_16[108]},
      {stage3_16[57]}
   );
   gpc1_1 gpc9266 (
      {stage2_16[109]},
      {stage3_16[58]}
   );
   gpc1_1 gpc9267 (
      {stage2_17[80]},
      {stage3_17[34]}
   );
   gpc1_1 gpc9268 (
      {stage2_17[81]},
      {stage3_17[35]}
   );
   gpc1_1 gpc9269 (
      {stage2_17[82]},
      {stage3_17[36]}
   );
   gpc1_1 gpc9270 (
      {stage2_17[83]},
      {stage3_17[37]}
   );
   gpc1_1 gpc9271 (
      {stage2_17[84]},
      {stage3_17[38]}
   );
   gpc1_1 gpc9272 (
      {stage2_17[85]},
      {stage3_17[39]}
   );
   gpc1_1 gpc9273 (
      {stage2_17[86]},
      {stage3_17[40]}
   );
   gpc1_1 gpc9274 (
      {stage2_17[87]},
      {stage3_17[41]}
   );
   gpc1_1 gpc9275 (
      {stage2_17[88]},
      {stage3_17[42]}
   );
   gpc1_1 gpc9276 (
      {stage2_17[89]},
      {stage3_17[43]}
   );
   gpc1_1 gpc9277 (
      {stage2_18[147]},
      {stage3_18[49]}
   );
   gpc1_1 gpc9278 (
      {stage2_18[148]},
      {stage3_18[50]}
   );
   gpc1_1 gpc9279 (
      {stage2_18[149]},
      {stage3_18[51]}
   );
   gpc1_1 gpc9280 (
      {stage2_18[150]},
      {stage3_18[52]}
   );
   gpc1_1 gpc9281 (
      {stage2_18[151]},
      {stage3_18[53]}
   );
   gpc1_1 gpc9282 (
      {stage2_18[152]},
      {stage3_18[54]}
   );
   gpc1_1 gpc9283 (
      {stage2_18[153]},
      {stage3_18[55]}
   );
   gpc1_1 gpc9284 (
      {stage2_18[154]},
      {stage3_18[56]}
   );
   gpc1_1 gpc9285 (
      {stage2_18[155]},
      {stage3_18[57]}
   );
   gpc1_1 gpc9286 (
      {stage2_18[156]},
      {stage3_18[58]}
   );
   gpc1_1 gpc9287 (
      {stage2_18[157]},
      {stage3_18[59]}
   );
   gpc1_1 gpc9288 (
      {stage2_18[158]},
      {stage3_18[60]}
   );
   gpc1_1 gpc9289 (
      {stage2_18[159]},
      {stage3_18[61]}
   );
   gpc1_1 gpc9290 (
      {stage2_18[160]},
      {stage3_18[62]}
   );
   gpc1_1 gpc9291 (
      {stage2_18[161]},
      {stage3_18[63]}
   );
   gpc1_1 gpc9292 (
      {stage2_20[72]},
      {stage3_20[42]}
   );
   gpc1_1 gpc9293 (
      {stage2_20[73]},
      {stage3_20[43]}
   );
   gpc1_1 gpc9294 (
      {stage2_20[74]},
      {stage3_20[44]}
   );
   gpc1_1 gpc9295 (
      {stage2_20[75]},
      {stage3_20[45]}
   );
   gpc1_1 gpc9296 (
      {stage2_20[76]},
      {stage3_20[46]}
   );
   gpc1_1 gpc9297 (
      {stage2_20[77]},
      {stage3_20[47]}
   );
   gpc1_1 gpc9298 (
      {stage2_20[78]},
      {stage3_20[48]}
   );
   gpc1_1 gpc9299 (
      {stage2_20[79]},
      {stage3_20[49]}
   );
   gpc1_1 gpc9300 (
      {stage2_20[80]},
      {stage3_20[50]}
   );
   gpc1_1 gpc9301 (
      {stage2_20[81]},
      {stage3_20[51]}
   );
   gpc1_1 gpc9302 (
      {stage2_20[82]},
      {stage3_20[52]}
   );
   gpc1_1 gpc9303 (
      {stage2_20[83]},
      {stage3_20[53]}
   );
   gpc1_1 gpc9304 (
      {stage2_20[84]},
      {stage3_20[54]}
   );
   gpc1_1 gpc9305 (
      {stage2_20[85]},
      {stage3_20[55]}
   );
   gpc1_1 gpc9306 (
      {stage2_20[86]},
      {stage3_20[56]}
   );
   gpc1_1 gpc9307 (
      {stage2_20[87]},
      {stage3_20[57]}
   );
   gpc1_1 gpc9308 (
      {stage2_21[86]},
      {stage3_21[37]}
   );
   gpc1_1 gpc9309 (
      {stage2_21[87]},
      {stage3_21[38]}
   );
   gpc1_1 gpc9310 (
      {stage2_21[88]},
      {stage3_21[39]}
   );
   gpc1_1 gpc9311 (
      {stage2_21[89]},
      {stage3_21[40]}
   );
   gpc1_1 gpc9312 (
      {stage2_21[90]},
      {stage3_21[41]}
   );
   gpc1_1 gpc9313 (
      {stage2_21[91]},
      {stage3_21[42]}
   );
   gpc1_1 gpc9314 (
      {stage2_21[92]},
      {stage3_21[43]}
   );
   gpc1_1 gpc9315 (
      {stage2_21[93]},
      {stage3_21[44]}
   );
   gpc1_1 gpc9316 (
      {stage2_21[94]},
      {stage3_21[45]}
   );
   gpc1_1 gpc9317 (
      {stage2_21[95]},
      {stage3_21[46]}
   );
   gpc1_1 gpc9318 (
      {stage2_21[96]},
      {stage3_21[47]}
   );
   gpc1_1 gpc9319 (
      {stage2_21[97]},
      {stage3_21[48]}
   );
   gpc1_1 gpc9320 (
      {stage2_21[98]},
      {stage3_21[49]}
   );
   gpc1_1 gpc9321 (
      {stage2_21[99]},
      {stage3_21[50]}
   );
   gpc1_1 gpc9322 (
      {stage2_21[100]},
      {stage3_21[51]}
   );
   gpc1_1 gpc9323 (
      {stage2_21[101]},
      {stage3_21[52]}
   );
   gpc1_1 gpc9324 (
      {stage2_21[102]},
      {stage3_21[53]}
   );
   gpc1_1 gpc9325 (
      {stage2_21[103]},
      {stage3_21[54]}
   );
   gpc1_1 gpc9326 (
      {stage2_21[104]},
      {stage3_21[55]}
   );
   gpc1_1 gpc9327 (
      {stage2_21[105]},
      {stage3_21[56]}
   );
   gpc1_1 gpc9328 (
      {stage2_21[106]},
      {stage3_21[57]}
   );
   gpc1_1 gpc9329 (
      {stage2_21[107]},
      {stage3_21[58]}
   );
   gpc1_1 gpc9330 (
      {stage2_21[108]},
      {stage3_21[59]}
   );
   gpc1_1 gpc9331 (
      {stage2_21[109]},
      {stage3_21[60]}
   );
   gpc1_1 gpc9332 (
      {stage2_21[110]},
      {stage3_21[61]}
   );
   gpc1_1 gpc9333 (
      {stage2_21[111]},
      {stage3_21[62]}
   );
   gpc1_1 gpc9334 (
      {stage2_22[108]},
      {stage3_22[48]}
   );
   gpc1_1 gpc9335 (
      {stage2_22[109]},
      {stage3_22[49]}
   );
   gpc1_1 gpc9336 (
      {stage2_23[89]},
      {stage3_23[40]}
   );
   gpc1_1 gpc9337 (
      {stage2_23[90]},
      {stage3_23[41]}
   );
   gpc1_1 gpc9338 (
      {stage2_23[91]},
      {stage3_23[42]}
   );
   gpc1_1 gpc9339 (
      {stage2_23[92]},
      {stage3_23[43]}
   );
   gpc1_1 gpc9340 (
      {stage2_23[93]},
      {stage3_23[44]}
   );
   gpc1_1 gpc9341 (
      {stage2_23[94]},
      {stage3_23[45]}
   );
   gpc1_1 gpc9342 (
      {stage2_23[95]},
      {stage3_23[46]}
   );
   gpc1_1 gpc9343 (
      {stage2_23[96]},
      {stage3_23[47]}
   );
   gpc1_1 gpc9344 (
      {stage2_23[97]},
      {stage3_23[48]}
   );
   gpc1_1 gpc9345 (
      {stage2_25[102]},
      {stage3_25[31]}
   );
   gpc1_1 gpc9346 (
      {stage2_25[103]},
      {stage3_25[32]}
   );
   gpc1_1 gpc9347 (
      {stage2_25[104]},
      {stage3_25[33]}
   );
   gpc1_1 gpc9348 (
      {stage2_25[105]},
      {stage3_25[34]}
   );
   gpc1_1 gpc9349 (
      {stage2_25[106]},
      {stage3_25[35]}
   );
   gpc1_1 gpc9350 (
      {stage2_25[107]},
      {stage3_25[36]}
   );
   gpc1_1 gpc9351 (
      {stage2_25[108]},
      {stage3_25[37]}
   );
   gpc1_1 gpc9352 (
      {stage2_25[109]},
      {stage3_25[38]}
   );
   gpc1_1 gpc9353 (
      {stage2_25[110]},
      {stage3_25[39]}
   );
   gpc1_1 gpc9354 (
      {stage2_25[111]},
      {stage3_25[40]}
   );
   gpc1_1 gpc9355 (
      {stage2_25[112]},
      {stage3_25[41]}
   );
   gpc1_1 gpc9356 (
      {stage2_25[113]},
      {stage3_25[42]}
   );
   gpc1_1 gpc9357 (
      {stage2_25[114]},
      {stage3_25[43]}
   );
   gpc1_1 gpc9358 (
      {stage2_25[115]},
      {stage3_25[44]}
   );
   gpc1_1 gpc9359 (
      {stage2_25[116]},
      {stage3_25[45]}
   );
   gpc1_1 gpc9360 (
      {stage2_25[117]},
      {stage3_25[46]}
   );
   gpc1_1 gpc9361 (
      {stage2_25[118]},
      {stage3_25[47]}
   );
   gpc1_1 gpc9362 (
      {stage2_25[119]},
      {stage3_25[48]}
   );
   gpc1_1 gpc9363 (
      {stage2_25[120]},
      {stage3_25[49]}
   );
   gpc1_1 gpc9364 (
      {stage2_25[121]},
      {stage3_25[50]}
   );
   gpc1_1 gpc9365 (
      {stage2_25[122]},
      {stage3_25[51]}
   );
   gpc1_1 gpc9366 (
      {stage2_26[126]},
      {stage3_26[47]}
   );
   gpc1_1 gpc9367 (
      {stage2_26[127]},
      {stage3_26[48]}
   );
   gpc1_1 gpc9368 (
      {stage2_26[128]},
      {stage3_26[49]}
   );
   gpc1_1 gpc9369 (
      {stage2_26[129]},
      {stage3_26[50]}
   );
   gpc1_1 gpc9370 (
      {stage2_26[130]},
      {stage3_26[51]}
   );
   gpc1_1 gpc9371 (
      {stage2_28[44]},
      {stage3_28[34]}
   );
   gpc1_1 gpc9372 (
      {stage2_28[45]},
      {stage3_28[35]}
   );
   gpc1_1 gpc9373 (
      {stage2_28[46]},
      {stage3_28[36]}
   );
   gpc1_1 gpc9374 (
      {stage2_28[47]},
      {stage3_28[37]}
   );
   gpc1_1 gpc9375 (
      {stage2_28[48]},
      {stage3_28[38]}
   );
   gpc1_1 gpc9376 (
      {stage2_28[49]},
      {stage3_28[39]}
   );
   gpc1_1 gpc9377 (
      {stage2_28[50]},
      {stage3_28[40]}
   );
   gpc1_1 gpc9378 (
      {stage2_28[51]},
      {stage3_28[41]}
   );
   gpc1_1 gpc9379 (
      {stage2_28[52]},
      {stage3_28[42]}
   );
   gpc1_1 gpc9380 (
      {stage2_28[53]},
      {stage3_28[43]}
   );
   gpc1_1 gpc9381 (
      {stage2_28[54]},
      {stage3_28[44]}
   );
   gpc1_1 gpc9382 (
      {stage2_28[55]},
      {stage3_28[45]}
   );
   gpc1_1 gpc9383 (
      {stage2_28[56]},
      {stage3_28[46]}
   );
   gpc1_1 gpc9384 (
      {stage2_28[57]},
      {stage3_28[47]}
   );
   gpc1_1 gpc9385 (
      {stage2_28[58]},
      {stage3_28[48]}
   );
   gpc1_1 gpc9386 (
      {stage2_28[59]},
      {stage3_28[49]}
   );
   gpc1_1 gpc9387 (
      {stage2_28[60]},
      {stage3_28[50]}
   );
   gpc1_1 gpc9388 (
      {stage2_28[61]},
      {stage3_28[51]}
   );
   gpc1_1 gpc9389 (
      {stage2_28[62]},
      {stage3_28[52]}
   );
   gpc1_1 gpc9390 (
      {stage2_28[63]},
      {stage3_28[53]}
   );
   gpc1_1 gpc9391 (
      {stage2_28[64]},
      {stage3_28[54]}
   );
   gpc1_1 gpc9392 (
      {stage2_28[65]},
      {stage3_28[55]}
   );
   gpc1_1 gpc9393 (
      {stage2_28[66]},
      {stage3_28[56]}
   );
   gpc1_1 gpc9394 (
      {stage2_28[67]},
      {stage3_28[57]}
   );
   gpc1_1 gpc9395 (
      {stage2_28[68]},
      {stage3_28[58]}
   );
   gpc1_1 gpc9396 (
      {stage2_28[69]},
      {stage3_28[59]}
   );
   gpc1_1 gpc9397 (
      {stage2_28[70]},
      {stage3_28[60]}
   );
   gpc1_1 gpc9398 (
      {stage2_28[71]},
      {stage3_28[61]}
   );
   gpc1_1 gpc9399 (
      {stage2_28[72]},
      {stage3_28[62]}
   );
   gpc1_1 gpc9400 (
      {stage2_28[73]},
      {stage3_28[63]}
   );
   gpc1_1 gpc9401 (
      {stage2_28[74]},
      {stage3_28[64]}
   );
   gpc1_1 gpc9402 (
      {stage2_28[75]},
      {stage3_28[65]}
   );
   gpc1_1 gpc9403 (
      {stage2_28[76]},
      {stage3_28[66]}
   );
   gpc1_1 gpc9404 (
      {stage2_28[77]},
      {stage3_28[67]}
   );
   gpc1_1 gpc9405 (
      {stage2_28[78]},
      {stage3_28[68]}
   );
   gpc1_1 gpc9406 (
      {stage2_28[79]},
      {stage3_28[69]}
   );
   gpc1_1 gpc9407 (
      {stage2_29[102]},
      {stage3_29[49]}
   );
   gpc1_1 gpc9408 (
      {stage2_29[103]},
      {stage3_29[50]}
   );
   gpc1_1 gpc9409 (
      {stage2_29[104]},
      {stage3_29[51]}
   );
   gpc1_1 gpc9410 (
      {stage2_29[105]},
      {stage3_29[52]}
   );
   gpc1_1 gpc9411 (
      {stage2_29[106]},
      {stage3_29[53]}
   );
   gpc1_1 gpc9412 (
      {stage2_29[107]},
      {stage3_29[54]}
   );
   gpc1_1 gpc9413 (
      {stage2_29[108]},
      {stage3_29[55]}
   );
   gpc1_1 gpc9414 (
      {stage2_29[109]},
      {stage3_29[56]}
   );
   gpc1_1 gpc9415 (
      {stage2_29[110]},
      {stage3_29[57]}
   );
   gpc1_1 gpc9416 (
      {stage2_29[111]},
      {stage3_29[58]}
   );
   gpc1_1 gpc9417 (
      {stage2_30[93]},
      {stage3_30[32]}
   );
   gpc1_1 gpc9418 (
      {stage2_30[94]},
      {stage3_30[33]}
   );
   gpc1_1 gpc9419 (
      {stage2_30[95]},
      {stage3_30[34]}
   );
   gpc1_1 gpc9420 (
      {stage2_30[96]},
      {stage3_30[35]}
   );
   gpc1_1 gpc9421 (
      {stage2_30[97]},
      {stage3_30[36]}
   );
   gpc1_1 gpc9422 (
      {stage2_30[98]},
      {stage3_30[37]}
   );
   gpc1_1 gpc9423 (
      {stage2_30[99]},
      {stage3_30[38]}
   );
   gpc1_1 gpc9424 (
      {stage2_31[124]},
      {stage3_31[38]}
   );
   gpc1_1 gpc9425 (
      {stage2_31[125]},
      {stage3_31[39]}
   );
   gpc1_1 gpc9426 (
      {stage2_31[126]},
      {stage3_31[40]}
   );
   gpc1_1 gpc9427 (
      {stage2_31[127]},
      {stage3_31[41]}
   );
   gpc1_1 gpc9428 (
      {stage2_32[112]},
      {stage3_32[50]}
   );
   gpc1_1 gpc9429 (
      {stage2_32[113]},
      {stage3_32[51]}
   );
   gpc1_1 gpc9430 (
      {stage2_32[114]},
      {stage3_32[52]}
   );
   gpc1_1 gpc9431 (
      {stage2_32[115]},
      {stage3_32[53]}
   );
   gpc1_1 gpc9432 (
      {stage2_32[116]},
      {stage3_32[54]}
   );
   gpc1_1 gpc9433 (
      {stage2_32[117]},
      {stage3_32[55]}
   );
   gpc1_1 gpc9434 (
      {stage2_33[91]},
      {stage3_33[45]}
   );
   gpc1_1 gpc9435 (
      {stage2_33[92]},
      {stage3_33[46]}
   );
   gpc1_1 gpc9436 (
      {stage2_33[93]},
      {stage3_33[47]}
   );
   gpc1_1 gpc9437 (
      {stage2_33[94]},
      {stage3_33[48]}
   );
   gpc1_1 gpc9438 (
      {stage2_33[95]},
      {stage3_33[49]}
   );
   gpc1_1 gpc9439 (
      {stage2_33[96]},
      {stage3_33[50]}
   );
   gpc1_1 gpc9440 (
      {stage2_33[97]},
      {stage3_33[51]}
   );
   gpc1_1 gpc9441 (
      {stage2_33[98]},
      {stage3_33[52]}
   );
   gpc1_1 gpc9442 (
      {stage2_33[99]},
      {stage3_33[53]}
   );
   gpc1_1 gpc9443 (
      {stage2_33[100]},
      {stage3_33[54]}
   );
   gpc1_1 gpc9444 (
      {stage2_33[101]},
      {stage3_33[55]}
   );
   gpc1_1 gpc9445 (
      {stage2_33[102]},
      {stage3_33[56]}
   );
   gpc1_1 gpc9446 (
      {stage2_33[103]},
      {stage3_33[57]}
   );
   gpc1_1 gpc9447 (
      {stage2_33[104]},
      {stage3_33[58]}
   );
   gpc1_1 gpc9448 (
      {stage2_33[105]},
      {stage3_33[59]}
   );
   gpc1_1 gpc9449 (
      {stage2_33[106]},
      {stage3_33[60]}
   );
   gpc1_1 gpc9450 (
      {stage2_33[107]},
      {stage3_33[61]}
   );
   gpc1_1 gpc9451 (
      {stage2_33[108]},
      {stage3_33[62]}
   );
   gpc1_1 gpc9452 (
      {stage2_36[114]},
      {stage3_36[50]}
   );
   gpc1_1 gpc9453 (
      {stage2_36[115]},
      {stage3_36[51]}
   );
   gpc1_1 gpc9454 (
      {stage2_36[116]},
      {stage3_36[52]}
   );
   gpc1_1 gpc9455 (
      {stage2_36[117]},
      {stage3_36[53]}
   );
   gpc1_1 gpc9456 (
      {stage2_36[118]},
      {stage3_36[54]}
   );
   gpc1_1 gpc9457 (
      {stage2_36[119]},
      {stage3_36[55]}
   );
   gpc1_1 gpc9458 (
      {stage2_38[81]},
      {stage3_38[50]}
   );
   gpc1_1 gpc9459 (
      {stage2_38[82]},
      {stage3_38[51]}
   );
   gpc1_1 gpc9460 (
      {stage2_38[83]},
      {stage3_38[52]}
   );
   gpc1_1 gpc9461 (
      {stage2_38[84]},
      {stage3_38[53]}
   );
   gpc1_1 gpc9462 (
      {stage2_38[85]},
      {stage3_38[54]}
   );
   gpc1_1 gpc9463 (
      {stage2_38[86]},
      {stage3_38[55]}
   );
   gpc1_1 gpc9464 (
      {stage2_38[87]},
      {stage3_38[56]}
   );
   gpc1_1 gpc9465 (
      {stage2_38[88]},
      {stage3_38[57]}
   );
   gpc1_1 gpc9466 (
      {stage2_38[89]},
      {stage3_38[58]}
   );
   gpc1_1 gpc9467 (
      {stage2_38[90]},
      {stage3_38[59]}
   );
   gpc1_1 gpc9468 (
      {stage2_38[91]},
      {stage3_38[60]}
   );
   gpc1_1 gpc9469 (
      {stage2_38[92]},
      {stage3_38[61]}
   );
   gpc1_1 gpc9470 (
      {stage2_38[93]},
      {stage3_38[62]}
   );
   gpc1_1 gpc9471 (
      {stage2_38[94]},
      {stage3_38[63]}
   );
   gpc1_1 gpc9472 (
      {stage2_38[95]},
      {stage3_38[64]}
   );
   gpc1_1 gpc9473 (
      {stage2_38[96]},
      {stage3_38[65]}
   );
   gpc1_1 gpc9474 (
      {stage2_38[97]},
      {stage3_38[66]}
   );
   gpc1_1 gpc9475 (
      {stage2_38[98]},
      {stage3_38[67]}
   );
   gpc1_1 gpc9476 (
      {stage2_38[99]},
      {stage3_38[68]}
   );
   gpc1_1 gpc9477 (
      {stage2_39[100]},
      {stage3_39[52]}
   );
   gpc1_1 gpc9478 (
      {stage2_39[101]},
      {stage3_39[53]}
   );
   gpc1_1 gpc9479 (
      {stage2_39[102]},
      {stage3_39[54]}
   );
   gpc1_1 gpc9480 (
      {stage2_39[103]},
      {stage3_39[55]}
   );
   gpc1_1 gpc9481 (
      {stage2_39[104]},
      {stage3_39[56]}
   );
   gpc1_1 gpc9482 (
      {stage2_39[105]},
      {stage3_39[57]}
   );
   gpc1_1 gpc9483 (
      {stage2_39[106]},
      {stage3_39[58]}
   );
   gpc1_1 gpc9484 (
      {stage2_39[107]},
      {stage3_39[59]}
   );
   gpc1_1 gpc9485 (
      {stage2_40[131]},
      {stage3_40[37]}
   );
   gpc1_1 gpc9486 (
      {stage2_40[132]},
      {stage3_40[38]}
   );
   gpc1_1 gpc9487 (
      {stage2_40[133]},
      {stage3_40[39]}
   );
   gpc1_1 gpc9488 (
      {stage2_40[134]},
      {stage3_40[40]}
   );
   gpc1_1 gpc9489 (
      {stage2_40[135]},
      {stage3_40[41]}
   );
   gpc1_1 gpc9490 (
      {stage2_40[136]},
      {stage3_40[42]}
   );
   gpc1_1 gpc9491 (
      {stage2_40[137]},
      {stage3_40[43]}
   );
   gpc1_1 gpc9492 (
      {stage2_40[138]},
      {stage3_40[44]}
   );
   gpc1_1 gpc9493 (
      {stage2_40[139]},
      {stage3_40[45]}
   );
   gpc1_1 gpc9494 (
      {stage2_41[102]},
      {stage3_41[36]}
   );
   gpc1_1 gpc9495 (
      {stage2_41[103]},
      {stage3_41[37]}
   );
   gpc1_1 gpc9496 (
      {stage2_41[104]},
      {stage3_41[38]}
   );
   gpc1_1 gpc9497 (
      {stage2_41[105]},
      {stage3_41[39]}
   );
   gpc1_1 gpc9498 (
      {stage2_41[106]},
      {stage3_41[40]}
   );
   gpc1_1 gpc9499 (
      {stage2_41[107]},
      {stage3_41[41]}
   );
   gpc1_1 gpc9500 (
      {stage2_41[108]},
      {stage3_41[42]}
   );
   gpc1_1 gpc9501 (
      {stage2_41[109]},
      {stage3_41[43]}
   );
   gpc1_1 gpc9502 (
      {stage2_41[110]},
      {stage3_41[44]}
   );
   gpc1_1 gpc9503 (
      {stage2_41[111]},
      {stage3_41[45]}
   );
   gpc1_1 gpc9504 (
      {stage2_41[112]},
      {stage3_41[46]}
   );
   gpc1_1 gpc9505 (
      {stage2_41[113]},
      {stage3_41[47]}
   );
   gpc1_1 gpc9506 (
      {stage2_41[114]},
      {stage3_41[48]}
   );
   gpc1_1 gpc9507 (
      {stage2_41[115]},
      {stage3_41[49]}
   );
   gpc1_1 gpc9508 (
      {stage2_41[116]},
      {stage3_41[50]}
   );
   gpc1_1 gpc9509 (
      {stage2_41[117]},
      {stage3_41[51]}
   );
   gpc1_1 gpc9510 (
      {stage2_41[118]},
      {stage3_41[52]}
   );
   gpc1_1 gpc9511 (
      {stage2_41[119]},
      {stage3_41[53]}
   );
   gpc1_1 gpc9512 (
      {stage2_41[120]},
      {stage3_41[54]}
   );
   gpc1_1 gpc9513 (
      {stage2_41[121]},
      {stage3_41[55]}
   );
   gpc1_1 gpc9514 (
      {stage2_41[122]},
      {stage3_41[56]}
   );
   gpc1_1 gpc9515 (
      {stage2_42[74]},
      {stage3_42[46]}
   );
   gpc1_1 gpc9516 (
      {stage2_42[75]},
      {stage3_42[47]}
   );
   gpc1_1 gpc9517 (
      {stage2_42[76]},
      {stage3_42[48]}
   );
   gpc1_1 gpc9518 (
      {stage2_42[77]},
      {stage3_42[49]}
   );
   gpc1_1 gpc9519 (
      {stage2_42[78]},
      {stage3_42[50]}
   );
   gpc1_1 gpc9520 (
      {stage2_42[79]},
      {stage3_42[51]}
   );
   gpc1_1 gpc9521 (
      {stage2_42[80]},
      {stage3_42[52]}
   );
   gpc1_1 gpc9522 (
      {stage2_42[81]},
      {stage3_42[53]}
   );
   gpc1_1 gpc9523 (
      {stage2_43[98]},
      {stage3_43[47]}
   );
   gpc1_1 gpc9524 (
      {stage2_43[99]},
      {stage3_43[48]}
   );
   gpc1_1 gpc9525 (
      {stage2_43[100]},
      {stage3_43[49]}
   );
   gpc1_1 gpc9526 (
      {stage2_43[101]},
      {stage3_43[50]}
   );
   gpc1_1 gpc9527 (
      {stage2_43[102]},
      {stage3_43[51]}
   );
   gpc1_1 gpc9528 (
      {stage2_43[103]},
      {stage3_43[52]}
   );
   gpc1_1 gpc9529 (
      {stage2_43[104]},
      {stage3_43[53]}
   );
   gpc1_1 gpc9530 (
      {stage2_43[105]},
      {stage3_43[54]}
   );
   gpc1_1 gpc9531 (
      {stage2_43[106]},
      {stage3_43[55]}
   );
   gpc1_1 gpc9532 (
      {stage2_43[107]},
      {stage3_43[56]}
   );
   gpc1_1 gpc9533 (
      {stage2_43[108]},
      {stage3_43[57]}
   );
   gpc1_1 gpc9534 (
      {stage2_43[109]},
      {stage3_43[58]}
   );
   gpc1_1 gpc9535 (
      {stage2_43[110]},
      {stage3_43[59]}
   );
   gpc1_1 gpc9536 (
      {stage2_44[86]},
      {stage3_44[33]}
   );
   gpc1_1 gpc9537 (
      {stage2_44[87]},
      {stage3_44[34]}
   );
   gpc1_1 gpc9538 (
      {stage2_44[88]},
      {stage3_44[35]}
   );
   gpc1_1 gpc9539 (
      {stage2_44[89]},
      {stage3_44[36]}
   );
   gpc1_1 gpc9540 (
      {stage2_44[90]},
      {stage3_44[37]}
   );
   gpc1_1 gpc9541 (
      {stage2_44[91]},
      {stage3_44[38]}
   );
   gpc1_1 gpc9542 (
      {stage2_44[92]},
      {stage3_44[39]}
   );
   gpc1_1 gpc9543 (
      {stage2_44[93]},
      {stage3_44[40]}
   );
   gpc1_1 gpc9544 (
      {stage2_44[94]},
      {stage3_44[41]}
   );
   gpc1_1 gpc9545 (
      {stage2_44[95]},
      {stage3_44[42]}
   );
   gpc1_1 gpc9546 (
      {stage2_44[96]},
      {stage3_44[43]}
   );
   gpc1_1 gpc9547 (
      {stage2_44[97]},
      {stage3_44[44]}
   );
   gpc1_1 gpc9548 (
      {stage2_44[98]},
      {stage3_44[45]}
   );
   gpc1_1 gpc9549 (
      {stage2_44[99]},
      {stage3_44[46]}
   );
   gpc1_1 gpc9550 (
      {stage2_44[100]},
      {stage3_44[47]}
   );
   gpc1_1 gpc9551 (
      {stage2_44[101]},
      {stage3_44[48]}
   );
   gpc1_1 gpc9552 (
      {stage2_44[102]},
      {stage3_44[49]}
   );
   gpc1_1 gpc9553 (
      {stage2_44[103]},
      {stage3_44[50]}
   );
   gpc1_1 gpc9554 (
      {stage2_44[104]},
      {stage3_44[51]}
   );
   gpc1_1 gpc9555 (
      {stage2_44[105]},
      {stage3_44[52]}
   );
   gpc1_1 gpc9556 (
      {stage2_44[106]},
      {stage3_44[53]}
   );
   gpc1_1 gpc9557 (
      {stage2_44[107]},
      {stage3_44[54]}
   );
   gpc1_1 gpc9558 (
      {stage2_44[108]},
      {stage3_44[55]}
   );
   gpc1_1 gpc9559 (
      {stage2_44[109]},
      {stage3_44[56]}
   );
   gpc1_1 gpc9560 (
      {stage2_44[110]},
      {stage3_44[57]}
   );
   gpc1_1 gpc9561 (
      {stage2_44[111]},
      {stage3_44[58]}
   );
   gpc1_1 gpc9562 (
      {stage2_44[112]},
      {stage3_44[59]}
   );
   gpc1_1 gpc9563 (
      {stage2_44[113]},
      {stage3_44[60]}
   );
   gpc1_1 gpc9564 (
      {stage2_44[114]},
      {stage3_44[61]}
   );
   gpc1_1 gpc9565 (
      {stage2_44[115]},
      {stage3_44[62]}
   );
   gpc1_1 gpc9566 (
      {stage2_44[116]},
      {stage3_44[63]}
   );
   gpc1_1 gpc9567 (
      {stage2_44[117]},
      {stage3_44[64]}
   );
   gpc1_1 gpc9568 (
      {stage2_44[118]},
      {stage3_44[65]}
   );
   gpc1_1 gpc9569 (
      {stage2_44[119]},
      {stage3_44[66]}
   );
   gpc1_1 gpc9570 (
      {stage2_44[120]},
      {stage3_44[67]}
   );
   gpc1_1 gpc9571 (
      {stage2_44[121]},
      {stage3_44[68]}
   );
   gpc1_1 gpc9572 (
      {stage2_44[122]},
      {stage3_44[69]}
   );
   gpc1_1 gpc9573 (
      {stage2_44[123]},
      {stage3_44[70]}
   );
   gpc1_1 gpc9574 (
      {stage2_44[124]},
      {stage3_44[71]}
   );
   gpc1_1 gpc9575 (
      {stage2_44[125]},
      {stage3_44[72]}
   );
   gpc1_1 gpc9576 (
      {stage2_44[126]},
      {stage3_44[73]}
   );
   gpc1_1 gpc9577 (
      {stage2_44[127]},
      {stage3_44[74]}
   );
   gpc1_1 gpc9578 (
      {stage2_44[128]},
      {stage3_44[75]}
   );
   gpc1_1 gpc9579 (
      {stage2_44[129]},
      {stage3_44[76]}
   );
   gpc1_1 gpc9580 (
      {stage2_44[130]},
      {stage3_44[77]}
   );
   gpc1_1 gpc9581 (
      {stage2_44[131]},
      {stage3_44[78]}
   );
   gpc1_1 gpc9582 (
      {stage2_44[132]},
      {stage3_44[79]}
   );
   gpc1_1 gpc9583 (
      {stage2_44[133]},
      {stage3_44[80]}
   );
   gpc1_1 gpc9584 (
      {stage2_44[134]},
      {stage3_44[81]}
   );
   gpc1_1 gpc9585 (
      {stage2_44[135]},
      {stage3_44[82]}
   );
   gpc1_1 gpc9586 (
      {stage2_44[136]},
      {stage3_44[83]}
   );
   gpc1_1 gpc9587 (
      {stage2_44[137]},
      {stage3_44[84]}
   );
   gpc1_1 gpc9588 (
      {stage2_45[126]},
      {stage3_45[34]}
   );
   gpc1_1 gpc9589 (
      {stage2_45[127]},
      {stage3_45[35]}
   );
   gpc1_1 gpc9590 (
      {stage2_45[128]},
      {stage3_45[36]}
   );
   gpc1_1 gpc9591 (
      {stage2_45[129]},
      {stage3_45[37]}
   );
   gpc1_1 gpc9592 (
      {stage2_45[130]},
      {stage3_45[38]}
   );
   gpc1_1 gpc9593 (
      {stage2_45[131]},
      {stage3_45[39]}
   );
   gpc1_1 gpc9594 (
      {stage2_47[83]},
      {stage3_47[49]}
   );
   gpc1_1 gpc9595 (
      {stage2_47[84]},
      {stage3_47[50]}
   );
   gpc1_1 gpc9596 (
      {stage2_47[85]},
      {stage3_47[51]}
   );
   gpc1_1 gpc9597 (
      {stage2_47[86]},
      {stage3_47[52]}
   );
   gpc1_1 gpc9598 (
      {stage2_47[87]},
      {stage3_47[53]}
   );
   gpc1_1 gpc9599 (
      {stage2_47[88]},
      {stage3_47[54]}
   );
   gpc1_1 gpc9600 (
      {stage2_47[89]},
      {stage3_47[55]}
   );
   gpc1_1 gpc9601 (
      {stage2_47[90]},
      {stage3_47[56]}
   );
   gpc1_1 gpc9602 (
      {stage2_47[91]},
      {stage3_47[57]}
   );
   gpc1_1 gpc9603 (
      {stage2_47[92]},
      {stage3_47[58]}
   );
   gpc1_1 gpc9604 (
      {stage2_47[93]},
      {stage3_47[59]}
   );
   gpc1_1 gpc9605 (
      {stage2_47[94]},
      {stage3_47[60]}
   );
   gpc1_1 gpc9606 (
      {stage2_47[95]},
      {stage3_47[61]}
   );
   gpc1_1 gpc9607 (
      {stage2_47[96]},
      {stage3_47[62]}
   );
   gpc1_1 gpc9608 (
      {stage2_47[97]},
      {stage3_47[63]}
   );
   gpc1_1 gpc9609 (
      {stage2_47[98]},
      {stage3_47[64]}
   );
   gpc1_1 gpc9610 (
      {stage2_47[99]},
      {stage3_47[65]}
   );
   gpc1_1 gpc9611 (
      {stage2_47[100]},
      {stage3_47[66]}
   );
   gpc1_1 gpc9612 (
      {stage2_47[101]},
      {stage3_47[67]}
   );
   gpc1_1 gpc9613 (
      {stage2_47[102]},
      {stage3_47[68]}
   );
   gpc1_1 gpc9614 (
      {stage2_47[103]},
      {stage3_47[69]}
   );
   gpc1_1 gpc9615 (
      {stage2_47[104]},
      {stage3_47[70]}
   );
   gpc1_1 gpc9616 (
      {stage2_47[105]},
      {stage3_47[71]}
   );
   gpc1_1 gpc9617 (
      {stage2_47[106]},
      {stage3_47[72]}
   );
   gpc1_1 gpc9618 (
      {stage2_47[107]},
      {stage3_47[73]}
   );
   gpc1_1 gpc9619 (
      {stage2_49[96]},
      {stage3_49[45]}
   );
   gpc1_1 gpc9620 (
      {stage2_49[97]},
      {stage3_49[46]}
   );
   gpc1_1 gpc9621 (
      {stage2_49[98]},
      {stage3_49[47]}
   );
   gpc1_1 gpc9622 (
      {stage2_49[99]},
      {stage3_49[48]}
   );
   gpc1_1 gpc9623 (
      {stage2_49[100]},
      {stage3_49[49]}
   );
   gpc1_1 gpc9624 (
      {stage2_49[101]},
      {stage3_49[50]}
   );
   gpc1_1 gpc9625 (
      {stage2_49[102]},
      {stage3_49[51]}
   );
   gpc1_1 gpc9626 (
      {stage2_49[103]},
      {stage3_49[52]}
   );
   gpc1_1 gpc9627 (
      {stage2_49[104]},
      {stage3_49[53]}
   );
   gpc1_1 gpc9628 (
      {stage2_49[105]},
      {stage3_49[54]}
   );
   gpc1_1 gpc9629 (
      {stage2_49[106]},
      {stage3_49[55]}
   );
   gpc1_1 gpc9630 (
      {stage2_49[107]},
      {stage3_49[56]}
   );
   gpc1_1 gpc9631 (
      {stage2_49[108]},
      {stage3_49[57]}
   );
   gpc1_1 gpc9632 (
      {stage2_49[109]},
      {stage3_49[58]}
   );
   gpc1_1 gpc9633 (
      {stage2_49[110]},
      {stage3_49[59]}
   );
   gpc1_1 gpc9634 (
      {stage2_49[111]},
      {stage3_49[60]}
   );
   gpc1_1 gpc9635 (
      {stage2_49[112]},
      {stage3_49[61]}
   );
   gpc1_1 gpc9636 (
      {stage2_49[113]},
      {stage3_49[62]}
   );
   gpc1_1 gpc9637 (
      {stage2_49[114]},
      {stage3_49[63]}
   );
   gpc1_1 gpc9638 (
      {stage2_49[115]},
      {stage3_49[64]}
   );
   gpc1_1 gpc9639 (
      {stage2_50[149]},
      {stage3_50[60]}
   );
   gpc1_1 gpc9640 (
      {stage2_50[150]},
      {stage3_50[61]}
   );
   gpc1_1 gpc9641 (
      {stage2_50[151]},
      {stage3_50[62]}
   );
   gpc1_1 gpc9642 (
      {stage2_50[152]},
      {stage3_50[63]}
   );
   gpc1_1 gpc9643 (
      {stage2_51[81]},
      {stage3_51[47]}
   );
   gpc1_1 gpc9644 (
      {stage2_51[82]},
      {stage3_51[48]}
   );
   gpc1_1 gpc9645 (
      {stage2_51[83]},
      {stage3_51[49]}
   );
   gpc1_1 gpc9646 (
      {stage2_51[84]},
      {stage3_51[50]}
   );
   gpc1_1 gpc9647 (
      {stage2_51[85]},
      {stage3_51[51]}
   );
   gpc1_1 gpc9648 (
      {stage2_51[86]},
      {stage3_51[52]}
   );
   gpc1_1 gpc9649 (
      {stage2_51[87]},
      {stage3_51[53]}
   );
   gpc1_1 gpc9650 (
      {stage2_52[109]},
      {stage3_52[37]}
   );
   gpc1_1 gpc9651 (
      {stage2_52[110]},
      {stage3_52[38]}
   );
   gpc1_1 gpc9652 (
      {stage2_52[111]},
      {stage3_52[39]}
   );
   gpc1_1 gpc9653 (
      {stage2_52[112]},
      {stage3_52[40]}
   );
   gpc1_1 gpc9654 (
      {stage2_52[113]},
      {stage3_52[41]}
   );
   gpc1_1 gpc9655 (
      {stage2_52[114]},
      {stage3_52[42]}
   );
   gpc1_1 gpc9656 (
      {stage2_52[115]},
      {stage3_52[43]}
   );
   gpc1_1 gpc9657 (
      {stage2_52[116]},
      {stage3_52[44]}
   );
   gpc1_1 gpc9658 (
      {stage2_52[117]},
      {stage3_52[45]}
   );
   gpc1_1 gpc9659 (
      {stage2_52[118]},
      {stage3_52[46]}
   );
   gpc1_1 gpc9660 (
      {stage2_52[119]},
      {stage3_52[47]}
   );
   gpc1_1 gpc9661 (
      {stage2_52[120]},
      {stage3_52[48]}
   );
   gpc1_1 gpc9662 (
      {stage2_52[121]},
      {stage3_52[49]}
   );
   gpc1_1 gpc9663 (
      {stage2_52[122]},
      {stage3_52[50]}
   );
   gpc1_1 gpc9664 (
      {stage2_52[123]},
      {stage3_52[51]}
   );
   gpc1_1 gpc9665 (
      {stage2_52[124]},
      {stage3_52[52]}
   );
   gpc1_1 gpc9666 (
      {stage2_52[125]},
      {stage3_52[53]}
   );
   gpc1_1 gpc9667 (
      {stage2_52[126]},
      {stage3_52[54]}
   );
   gpc1_1 gpc9668 (
      {stage2_52[127]},
      {stage3_52[55]}
   );
   gpc1_1 gpc9669 (
      {stage2_53[89]},
      {stage3_53[45]}
   );
   gpc1_1 gpc9670 (
      {stage2_53[90]},
      {stage3_53[46]}
   );
   gpc1_1 gpc9671 (
      {stage2_53[91]},
      {stage3_53[47]}
   );
   gpc1_1 gpc9672 (
      {stage2_53[92]},
      {stage3_53[48]}
   );
   gpc1_1 gpc9673 (
      {stage2_53[93]},
      {stage3_53[49]}
   );
   gpc1_1 gpc9674 (
      {stage2_53[94]},
      {stage3_53[50]}
   );
   gpc1_1 gpc9675 (
      {stage2_53[95]},
      {stage3_53[51]}
   );
   gpc1_1 gpc9676 (
      {stage2_53[96]},
      {stage3_53[52]}
   );
   gpc1_1 gpc9677 (
      {stage2_54[114]},
      {stage3_54[53]}
   );
   gpc1_1 gpc9678 (
      {stage2_54[115]},
      {stage3_54[54]}
   );
   gpc1_1 gpc9679 (
      {stage2_54[116]},
      {stage3_54[55]}
   );
   gpc1_1 gpc9680 (
      {stage2_54[117]},
      {stage3_54[56]}
   );
   gpc1_1 gpc9681 (
      {stage2_54[118]},
      {stage3_54[57]}
   );
   gpc1_1 gpc9682 (
      {stage2_54[119]},
      {stage3_54[58]}
   );
   gpc1_1 gpc9683 (
      {stage2_54[120]},
      {stage3_54[59]}
   );
   gpc1_1 gpc9684 (
      {stage2_54[121]},
      {stage3_54[60]}
   );
   gpc1_1 gpc9685 (
      {stage2_54[122]},
      {stage3_54[61]}
   );
   gpc1_1 gpc9686 (
      {stage2_54[123]},
      {stage3_54[62]}
   );
   gpc1_1 gpc9687 (
      {stage2_55[102]},
      {stage3_55[38]}
   );
   gpc1_1 gpc9688 (
      {stage2_55[103]},
      {stage3_55[39]}
   );
   gpc1_1 gpc9689 (
      {stage2_55[104]},
      {stage3_55[40]}
   );
   gpc1_1 gpc9690 (
      {stage2_55[105]},
      {stage3_55[41]}
   );
   gpc1_1 gpc9691 (
      {stage2_55[106]},
      {stage3_55[42]}
   );
   gpc1_1 gpc9692 (
      {stage2_55[107]},
      {stage3_55[43]}
   );
   gpc1_1 gpc9693 (
      {stage2_55[108]},
      {stage3_55[44]}
   );
   gpc1_1 gpc9694 (
      {stage2_55[109]},
      {stage3_55[45]}
   );
   gpc1_1 gpc9695 (
      {stage2_55[110]},
      {stage3_55[46]}
   );
   gpc1_1 gpc9696 (
      {stage2_57[72]},
      {stage3_57[46]}
   );
   gpc1_1 gpc9697 (
      {stage2_57[73]},
      {stage3_57[47]}
   );
   gpc1_1 gpc9698 (
      {stage2_57[74]},
      {stage3_57[48]}
   );
   gpc1_1 gpc9699 (
      {stage2_57[75]},
      {stage3_57[49]}
   );
   gpc1_1 gpc9700 (
      {stage2_57[76]},
      {stage3_57[50]}
   );
   gpc1_1 gpc9701 (
      {stage2_57[77]},
      {stage3_57[51]}
   );
   gpc1_1 gpc9702 (
      {stage2_57[78]},
      {stage3_57[52]}
   );
   gpc1_1 gpc9703 (
      {stage2_58[79]},
      {stage3_58[43]}
   );
   gpc1_1 gpc9704 (
      {stage2_58[80]},
      {stage3_58[44]}
   );
   gpc1_1 gpc9705 (
      {stage2_58[81]},
      {stage3_58[45]}
   );
   gpc1_1 gpc9706 (
      {stage2_58[82]},
      {stage3_58[46]}
   );
   gpc1_1 gpc9707 (
      {stage2_58[83]},
      {stage3_58[47]}
   );
   gpc1_1 gpc9708 (
      {stage2_58[84]},
      {stage3_58[48]}
   );
   gpc1_1 gpc9709 (
      {stage2_59[133]},
      {stage3_59[39]}
   );
   gpc1_1 gpc9710 (
      {stage2_59[134]},
      {stage3_59[40]}
   );
   gpc1_1 gpc9711 (
      {stage2_59[135]},
      {stage3_59[41]}
   );
   gpc1_1 gpc9712 (
      {stage2_59[136]},
      {stage3_59[42]}
   );
   gpc1_1 gpc9713 (
      {stage2_59[137]},
      {stage3_59[43]}
   );
   gpc1_1 gpc9714 (
      {stage2_59[138]},
      {stage3_59[44]}
   );
   gpc1_1 gpc9715 (
      {stage2_59[139]},
      {stage3_59[45]}
   );
   gpc1_1 gpc9716 (
      {stage2_60[106]},
      {stage3_60[48]}
   );
   gpc1_1 gpc9717 (
      {stage2_60[107]},
      {stage3_60[49]}
   );
   gpc1_1 gpc9718 (
      {stage2_60[108]},
      {stage3_60[50]}
   );
   gpc1_1 gpc9719 (
      {stage2_60[109]},
      {stage3_60[51]}
   );
   gpc1_1 gpc9720 (
      {stage2_60[110]},
      {stage3_60[52]}
   );
   gpc1_1 gpc9721 (
      {stage2_61[90]},
      {stage3_61[45]}
   );
   gpc1_1 gpc9722 (
      {stage2_61[91]},
      {stage3_61[46]}
   );
   gpc1_1 gpc9723 (
      {stage2_61[92]},
      {stage3_61[47]}
   );
   gpc1_1 gpc9724 (
      {stage2_61[93]},
      {stage3_61[48]}
   );
   gpc1_1 gpc9725 (
      {stage2_61[94]},
      {stage3_61[49]}
   );
   gpc1_1 gpc9726 (
      {stage2_61[95]},
      {stage3_61[50]}
   );
   gpc1_1 gpc9727 (
      {stage2_61[96]},
      {stage3_61[51]}
   );
   gpc1_1 gpc9728 (
      {stage2_61[97]},
      {stage3_61[52]}
   );
   gpc1_1 gpc9729 (
      {stage2_61[98]},
      {stage3_61[53]}
   );
   gpc1_1 gpc9730 (
      {stage2_61[99]},
      {stage3_61[54]}
   );
   gpc1_1 gpc9731 (
      {stage2_61[100]},
      {stage3_61[55]}
   );
   gpc1_1 gpc9732 (
      {stage2_61[101]},
      {stage3_61[56]}
   );
   gpc1_1 gpc9733 (
      {stage2_62[144]},
      {stage3_62[40]}
   );
   gpc1_1 gpc9734 (
      {stage2_63[95]},
      {stage3_63[54]}
   );
   gpc1_1 gpc9735 (
      {stage2_63[96]},
      {stage3_63[55]}
   );
   gpc1_1 gpc9736 (
      {stage2_63[97]},
      {stage3_63[56]}
   );
   gpc1_1 gpc9737 (
      {stage2_63[98]},
      {stage3_63[57]}
   );
   gpc1_1 gpc9738 (
      {stage2_63[99]},
      {stage3_63[58]}
   );
   gpc1_1 gpc9739 (
      {stage2_63[100]},
      {stage3_63[59]}
   );
   gpc1_1 gpc9740 (
      {stage2_63[101]},
      {stage3_63[60]}
   );
   gpc1_1 gpc9741 (
      {stage2_63[102]},
      {stage3_63[61]}
   );
   gpc1_1 gpc9742 (
      {stage2_63[103]},
      {stage3_63[62]}
   );
   gpc1_1 gpc9743 (
      {stage2_63[104]},
      {stage3_63[63]}
   );
   gpc1_1 gpc9744 (
      {stage2_63[105]},
      {stage3_63[64]}
   );
   gpc1_1 gpc9745 (
      {stage2_63[106]},
      {stage3_63[65]}
   );
   gpc1_1 gpc9746 (
      {stage2_63[107]},
      {stage3_63[66]}
   );
   gpc1_1 gpc9747 (
      {stage2_63[108]},
      {stage3_63[67]}
   );
   gpc1_1 gpc9748 (
      {stage2_63[109]},
      {stage3_63[68]}
   );
   gpc1_1 gpc9749 (
      {stage2_63[110]},
      {stage3_63[69]}
   );
   gpc1_1 gpc9750 (
      {stage2_63[111]},
      {stage3_63[70]}
   );
   gpc1_1 gpc9751 (
      {stage2_63[112]},
      {stage3_63[71]}
   );
   gpc1_1 gpc9752 (
      {stage2_64[95]},
      {stage3_64[44]}
   );
   gpc1_1 gpc9753 (
      {stage2_64[96]},
      {stage3_64[45]}
   );
   gpc1_1 gpc9754 (
      {stage2_64[97]},
      {stage3_64[46]}
   );
   gpc1_1 gpc9755 (
      {stage2_64[98]},
      {stage3_64[47]}
   );
   gpc1_1 gpc9756 (
      {stage2_64[99]},
      {stage3_64[48]}
   );
   gpc1_1 gpc9757 (
      {stage2_64[100]},
      {stage3_64[49]}
   );
   gpc1_1 gpc9758 (
      {stage2_64[101]},
      {stage3_64[50]}
   );
   gpc1_1 gpc9759 (
      {stage2_65[65]},
      {stage3_65[30]}
   );
   gpc1_1 gpc9760 (
      {stage2_65[66]},
      {stage3_65[31]}
   );
   gpc1_1 gpc9761 (
      {stage2_65[67]},
      {stage3_65[32]}
   );
   gpc1_1 gpc9762 (
      {stage2_66[30]},
      {stage3_66[30]}
   );
   gpc1_1 gpc9763 (
      {stage2_66[31]},
      {stage3_66[31]}
   );
   gpc1_1 gpc9764 (
      {stage2_66[32]},
      {stage3_66[32]}
   );
   gpc1_1 gpc9765 (
      {stage2_66[33]},
      {stage3_66[33]}
   );
   gpc1_1 gpc9766 (
      {stage2_66[34]},
      {stage3_66[34]}
   );
   gpc1_1 gpc9767 (
      {stage2_66[35]},
      {stage3_66[35]}
   );
   gpc1_1 gpc9768 (
      {stage2_66[36]},
      {stage3_66[36]}
   );
   gpc1_1 gpc9769 (
      {stage2_66[37]},
      {stage3_66[37]}
   );
   gpc1_1 gpc9770 (
      {stage2_66[38]},
      {stage3_66[38]}
   );
   gpc1_1 gpc9771 (
      {stage2_66[39]},
      {stage3_66[39]}
   );
   gpc1_1 gpc9772 (
      {stage2_66[40]},
      {stage3_66[40]}
   );
   gpc1_1 gpc9773 (
      {stage2_66[41]},
      {stage3_66[41]}
   );
   gpc1_1 gpc9774 (
      {stage2_66[42]},
      {stage3_66[42]}
   );
   gpc1_1 gpc9775 (
      {stage2_66[43]},
      {stage3_66[43]}
   );
   gpc1_1 gpc9776 (
      {stage2_66[44]},
      {stage3_66[44]}
   );
   gpc1_1 gpc9777 (
      {stage2_66[45]},
      {stage3_66[45]}
   );
   gpc1_1 gpc9778 (
      {stage2_66[46]},
      {stage3_66[46]}
   );
   gpc1_1 gpc9779 (
      {stage2_66[47]},
      {stage3_66[47]}
   );
   gpc1_1 gpc9780 (
      {stage2_66[48]},
      {stage3_66[48]}
   );
   gpc1_1 gpc9781 (
      {stage2_66[49]},
      {stage3_66[49]}
   );
   gpc1_1 gpc9782 (
      {stage2_66[50]},
      {stage3_66[50]}
   );
   gpc1_1 gpc9783 (
      {stage2_66[51]},
      {stage3_66[51]}
   );
   gpc1_1 gpc9784 (
      {stage2_66[52]},
      {stage3_66[52]}
   );
   gpc1_1 gpc9785 (
      {stage2_66[53]},
      {stage3_66[53]}
   );
   gpc606_5 gpc9786 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc9787 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc9788 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc9789 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc9790 (
      {stage3_1[18], stage3_1[19], stage3_1[20], stage3_1[21], stage3_1[22], stage3_1[23]},
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc9791 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc9792 (
      {stage3_3[24], stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc9793 (
      {stage3_3[29], stage3_3[30], stage3_3[31], stage3_3[32], stage3_3[33]},
      {stage3_4[7]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc9794 (
      {stage3_3[34], stage3_3[35], stage3_3[36], stage3_3[37], stage3_3[38]},
      {stage3_4[8]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[3],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc9795 (
      {stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[4],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc9796 (
      {stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[5],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc9797 (
      {stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[5],stage4_6[6],stage4_5[10],stage4_4[11]}
   );
   gpc606_5 gpc9798 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[3],stage4_7[6],stage4_6[7],stage4_5[11],stage4_4[12]}
   );
   gpc606_5 gpc9799 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[4],stage4_7[7],stage4_6[8],stage4_5[12],stage4_4[13]}
   );
   gpc606_5 gpc9800 (
      {stage3_4[39], stage3_4[40], stage3_4[41], stage3_4[42], stage3_4[43], stage3_4[44]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[5],stage4_7[8],stage4_6[9],stage4_5[13],stage4_4[14]}
   );
   gpc606_5 gpc9801 (
      {stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48], stage3_4[49], stage3_4[50]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[6],stage4_7[9],stage4_6[10],stage4_5[14],stage4_4[15]}
   );
   gpc606_5 gpc9802 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[7],stage4_7[10],stage4_6[11],stage4_5[15]}
   );
   gpc615_5 gpc9803 (
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[8],stage4_7[11],stage4_6[12]}
   );
   gpc615_5 gpc9804 (
      {stage3_6[47], stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[9],stage4_7[12],stage4_6[13]}
   );
   gpc615_5 gpc9805 (
      {stage3_6[52], stage3_6[53], stage3_6[54], stage3_6[55], stage3_6[56]},
      {stage3_7[8]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[10],stage4_7[13],stage4_6[14]}
   );
   gpc615_5 gpc9806 (
      {stage3_6[57], stage3_6[58], stage3_6[59], stage3_6[60], stage3_6[61]},
      {stage3_7[9]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[4],stage4_8[11],stage4_7[14],stage4_6[15]}
   );
   gpc615_5 gpc9807 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[24]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[4],stage4_9[5],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc9808 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[25]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[5],stage4_9[6],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc9809 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[26]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[6],stage4_9[7],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc9810 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[27]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[7],stage4_9[8],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc9811 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[28]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[8],stage4_9[9],stage4_8[16],stage4_7[19]}
   );
   gpc606_5 gpc9812 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[5],stage4_10[9],stage4_9[10]}
   );
   gpc606_5 gpc9813 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[6],stage4_10[10],stage4_9[11]}
   );
   gpc606_5 gpc9814 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[7],stage4_10[11],stage4_9[12]}
   );
   gpc606_5 gpc9815 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], 1'b0},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[8],stage4_10[12],stage4_9[13]}
   );
   gpc615_5 gpc9816 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[24]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[4],stage4_12[4],stage4_11[9],stage4_10[13]}
   );
   gpc615_5 gpc9817 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[25]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[5],stage4_12[5],stage4_11[10],stage4_10[14]}
   );
   gpc615_5 gpc9818 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[26]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[6],stage4_12[6],stage4_11[11],stage4_10[15]}
   );
   gpc615_5 gpc9819 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[27]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[7],stage4_12[7],stage4_11[12],stage4_10[16]}
   );
   gpc615_5 gpc9820 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24]},
      {stage3_11[28]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[8],stage4_12[8],stage4_11[13],stage4_10[17]}
   );
   gpc615_5 gpc9821 (
      {stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29]},
      {stage3_11[29]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[9],stage4_12[9],stage4_11[14],stage4_10[18]}
   );
   gpc615_5 gpc9822 (
      {stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33], stage3_10[34]},
      {stage3_11[30]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[10],stage4_12[10],stage4_11[15],stage4_10[19]}
   );
   gpc615_5 gpc9823 (
      {stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38], stage3_10[39]},
      {stage3_11[31]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[11],stage4_12[11],stage4_11[16],stage4_10[20]}
   );
   gpc615_5 gpc9824 (
      {stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43], stage3_10[44]},
      {stage3_11[32]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[12],stage4_12[12],stage4_11[17],stage4_10[21]}
   );
   gpc615_5 gpc9825 (
      {stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48], stage3_10[49]},
      {stage3_11[33]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[13],stage4_12[13],stage4_11[18],stage4_10[22]}
   );
   gpc615_5 gpc9826 (
      {stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53], stage3_10[54]},
      {stage3_11[34]},
      {stage3_12[60], stage3_12[61], stage3_12[62], stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage4_14[10],stage4_13[14],stage4_12[14],stage4_11[19],stage4_10[23]}
   );
   gpc615_5 gpc9827 (
      {stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58], stage3_10[59]},
      {stage3_11[35]},
      {stage3_12[66], stage3_12[67], stage3_12[68], stage3_12[69], stage3_12[70], stage3_12[71]},
      {stage4_14[11],stage4_13[15],stage4_12[15],stage4_11[20],stage4_10[24]}
   );
   gpc615_5 gpc9828 (
      {stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63], stage3_10[64]},
      {stage3_11[36]},
      {stage3_12[72], stage3_12[73], stage3_12[74], stage3_12[75], stage3_12[76], stage3_12[77]},
      {stage4_14[12],stage4_13[16],stage4_12[16],stage4_11[21],stage4_10[25]}
   );
   gpc615_5 gpc9829 (
      {stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[78]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[13],stage4_13[17],stage4_12[17],stage4_11[22]}
   );
   gpc615_5 gpc9830 (
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46]},
      {stage3_12[79]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[14],stage4_13[18],stage4_12[18],stage4_11[23]}
   );
   gpc615_5 gpc9831 (
      {stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51]},
      {stage3_12[80]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[15],stage4_13[19],stage4_12[19],stage4_11[24]}
   );
   gpc117_4 gpc9832 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[3],stage4_14[16],stage4_13[20]}
   );
   gpc606_5 gpc9833 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6]},
      {stage4_17[0],stage4_16[1],stage4_15[4],stage4_14[17],stage4_13[21]}
   );
   gpc606_5 gpc9834 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage4_17[1],stage4_16[2],stage4_15[5],stage4_14[18],stage4_13[22]}
   );
   gpc606_5 gpc9835 (
      {stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42]},
      {stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18]},
      {stage4_17[2],stage4_16[3],stage4_15[6],stage4_14[19],stage4_13[23]}
   );
   gpc615_5 gpc9836 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_15[19]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[3],stage4_16[4],stage4_15[7],stage4_14[20]}
   );
   gpc615_5 gpc9837 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[20]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[4],stage4_16[5],stage4_15[8],stage4_14[21]}
   );
   gpc615_5 gpc9838 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[21]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[5],stage4_16[6],stage4_15[9],stage4_14[22]}
   );
   gpc615_5 gpc9839 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[22]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[6],stage4_16[7],stage4_15[10],stage4_14[23]}
   );
   gpc615_5 gpc9840 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[23]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[7],stage4_16[8],stage4_15[11],stage4_14[24]}
   );
   gpc615_5 gpc9841 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[24]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[8],stage4_16[9],stage4_15[12],stage4_14[25]}
   );
   gpc615_5 gpc9842 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[9],stage4_16[10],stage4_15[13]}
   );
   gpc615_5 gpc9843 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[37]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[7],stage4_17[10],stage4_16[11],stage4_15[14]}
   );
   gpc615_5 gpc9844 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[38]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[8],stage4_17[11],stage4_16[12],stage4_15[15]}
   );
   gpc615_5 gpc9845 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[39]},
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage4_19[3],stage4_18[9],stage4_17[12],stage4_16[13],stage4_15[16]}
   );
   gpc606_5 gpc9846 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[4],stage4_18[10],stage4_17[13]}
   );
   gpc606_5 gpc9847 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[5],stage4_18[11],stage4_17[14]}
   );
   gpc207_4 gpc9848 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[2],stage4_20[2],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc9849 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[3],stage4_20[3],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc9850 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[4],stage4_20[4],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc9851 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[5],stage4_20[5],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc9852 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[6],stage4_20[6],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc9853 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[7],stage4_20[7],stage4_19[11],stage4_18[17]}
   );
   gpc615_5 gpc9854 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46]},
      {stage3_19[12]},
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage4_22[0],stage4_21[8],stage4_20[8],stage4_19[12],stage4_18[18]}
   );
   gpc615_5 gpc9855 (
      {stage3_18[47], stage3_18[48], stage3_18[49], stage3_18[50], stage3_18[51]},
      {stage3_19[13]},
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage4_22[1],stage4_21[9],stage4_20[9],stage4_19[13],stage4_18[19]}
   );
   gpc606_5 gpc9856 (
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[2],stage4_21[10],stage4_20[10],stage4_19[14]}
   );
   gpc606_5 gpc9857 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[3],stage4_21[11],stage4_20[11],stage4_19[15]}
   );
   gpc615_5 gpc9858 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[24]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[4],stage4_21[12],stage4_20[12],stage4_19[16]}
   );
   gpc615_5 gpc9859 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35]},
      {stage3_20[25]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[5],stage4_21[13],stage4_20[13],stage4_19[17]}
   );
   gpc615_5 gpc9860 (
      {stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40]},
      {stage3_20[26]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[6],stage4_21[14],stage4_20[14],stage4_19[18]}
   );
   gpc615_5 gpc9861 (
      {stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45]},
      {stage3_20[27]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[7],stage4_21[15],stage4_20[15],stage4_19[19]}
   );
   gpc606_5 gpc9862 (
      {stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31], stage3_20[32], stage3_20[33]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[6],stage4_22[8],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc9863 (
      {stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37], stage3_20[38], stage3_20[39]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[7],stage4_22[9],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc9864 (
      {stage3_20[40], stage3_20[41], stage3_20[42], stage3_20[43], stage3_20[44], stage3_20[45]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[8],stage4_22[10],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc9865 (
      {stage3_20[46], stage3_20[47], stage3_20[48], stage3_20[49], stage3_20[50], stage3_20[51]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[9],stage4_22[11],stage4_21[19],stage4_20[19]}
   );
   gpc615_5 gpc9866 (
      {stage3_20[52], stage3_20[53], stage3_20[54], stage3_20[55], stage3_20[56]},
      {stage3_21[36]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[10],stage4_22[12],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc9867 (
      {stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[5],stage4_23[11],stage4_22[13],stage4_21[21]}
   );
   gpc606_5 gpc9868 (
      {stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[6],stage4_23[12],stage4_22[14],stage4_21[22]}
   );
   gpc606_5 gpc9869 (
      {stage3_21[49], stage3_21[50], stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[7],stage4_23[13],stage4_22[15],stage4_21[23]}
   );
   gpc606_5 gpc9870 (
      {stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59], stage3_21[60]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[8],stage4_23[14],stage4_22[16],stage4_21[24]}
   );
   gpc615_5 gpc9871 (
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[9],stage4_23[15],stage4_22[17]}
   );
   gpc615_5 gpc9872 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[10],stage4_23[16],stage4_22[18]}
   );
   gpc615_5 gpc9873 (
      {stage3_22[40], stage3_22[41], stage3_22[42], stage3_22[43], stage3_22[44]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[11],stage4_23[17],stage4_22[19]}
   );
   gpc615_5 gpc9874 (
      {stage3_22[45], stage3_22[46], stage3_22[47], stage3_22[48], stage3_22[49]},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[12],stage4_23[18],stage4_22[20]}
   );
   gpc615_5 gpc9875 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[13],stage4_23[19]}
   );
   gpc615_5 gpc9876 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[14],stage4_23[20]}
   );
   gpc615_5 gpc9877 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[15],stage4_23[21]}
   );
   gpc615_5 gpc9878 (
      {stage3_23[43], stage3_23[44], stage3_23[45], stage3_23[46], stage3_23[47]},
      {stage3_24[27]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[7],stage4_25[11],stage4_24[16],stage4_23[22]}
   );
   gpc615_5 gpc9879 (
      {stage3_23[48], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_24[28]},
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage4_27[4],stage4_26[8],stage4_25[12],stage4_24[17],stage4_23[23]}
   );
   gpc606_5 gpc9880 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[5],stage4_26[9],stage4_25[13]}
   );
   gpc606_5 gpc9881 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[6],stage4_26[10],stage4_25[14]}
   );
   gpc606_5 gpc9882 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46], stage3_25[47]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[7],stage4_26[11],stage4_25[15]}
   );
   gpc606_5 gpc9883 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[3],stage4_28[3],stage4_27[8],stage4_26[12]}
   );
   gpc606_5 gpc9884 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[4],stage4_28[4],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc9885 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[5],stage4_28[5],stage4_27[10],stage4_26[14]}
   );
   gpc606_5 gpc9886 (
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[6],stage4_28[6],stage4_27[11],stage4_26[15]}
   );
   gpc606_5 gpc9887 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage4_30[4],stage4_29[7],stage4_28[7],stage4_27[12],stage4_26[16]}
   );
   gpc606_5 gpc9888 (
      {stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage4_30[5],stage4_29[8],stage4_28[8],stage4_27[13],stage4_26[17]}
   );
   gpc606_5 gpc9889 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40], stage3_26[41]},
      {stage3_28[36], stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41]},
      {stage4_30[6],stage4_29[9],stage4_28[9],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc9890 (
      {stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47]},
      {stage3_28[42], stage3_28[43], stage3_28[44], stage3_28[45], stage3_28[46], stage3_28[47]},
      {stage4_30[7],stage4_29[10],stage4_28[10],stage4_27[15],stage4_26[19]}
   );
   gpc606_5 gpc9891 (
      {stage3_26[48], stage3_26[49], stage3_26[50], stage3_26[51], 1'b0, 1'b0},
      {stage3_28[48], stage3_28[49], stage3_28[50], stage3_28[51], stage3_28[52], stage3_28[53]},
      {stage4_30[8],stage4_29[11],stage4_28[11],stage4_27[16],stage4_26[20]}
   );
   gpc606_5 gpc9892 (
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[9],stage4_29[12],stage4_28[12],stage4_27[17]}
   );
   gpc606_5 gpc9893 (
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[10],stage4_29[13],stage4_28[13],stage4_27[18]}
   );
   gpc606_5 gpc9894 (
      {stage3_27[30], stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[11],stage4_29[14],stage4_28[14],stage4_27[19]}
   );
   gpc606_5 gpc9895 (
      {stage3_27[36], stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[12],stage4_29[15],stage4_28[15],stage4_27[20]}
   );
   gpc1163_5 gpc9896 (
      {stage3_29[24], stage3_29[25], stage3_29[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[4],stage4_30[13],stage4_29[16]}
   );
   gpc1163_5 gpc9897 (
      {stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[5],stage4_30[14],stage4_29[17]}
   );
   gpc1163_5 gpc9898 (
      {stage3_29[30], stage3_29[31], stage3_29[32]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[6],stage4_30[15],stage4_29[18]}
   );
   gpc1163_5 gpc9899 (
      {stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[7],stage4_30[16],stage4_29[19]}
   );
   gpc606_5 gpc9900 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[4],stage4_32[4],stage4_31[8],stage4_30[17],stage4_29[20]}
   );
   gpc606_5 gpc9901 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15]},
      {stage4_33[5],stage4_32[5],stage4_31[9],stage4_30[18],stage4_29[21]}
   );
   gpc606_5 gpc9902 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52], stage3_29[53]},
      {stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21]},
      {stage4_33[6],stage4_32[6],stage4_31[10],stage4_30[19],stage4_29[22]}
   );
   gpc606_5 gpc9903 (
      {stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57], stage3_29[58], 1'b0},
      {stage3_31[22], stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage4_33[7],stage4_32[7],stage4_31[11],stage4_30[20],stage4_29[23]}
   );
   gpc606_5 gpc9904 (
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_32[4], stage3_32[5], stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9]},
      {stage4_34[0],stage4_33[8],stage4_32[8],stage4_31[12],stage4_30[21]}
   );
   gpc606_5 gpc9905 (
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage4_34[1],stage4_33[9],stage4_32[9],stage4_31[13],stage4_30[22]}
   );
   gpc615_5 gpc9906 (
      {stage3_31[28], stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32]},
      {stage3_32[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[10],stage4_32[10],stage4_31[14]}
   );
   gpc615_5 gpc9907 (
      {stage3_31[33], stage3_31[34], stage3_31[35], stage3_31[36], stage3_31[37]},
      {stage3_32[17]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[11],stage4_32[11],stage4_31[15]}
   );
   gpc615_5 gpc9908 (
      {stage3_31[38], stage3_31[39], stage3_31[40], stage3_31[41], 1'b0},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[12],stage4_32[12],stage4_31[16]}
   );
   gpc2116_5 gpc9909 (
      {stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24]},
      {stage3_33[18]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[13],stage4_32[13]}
   );
   gpc2116_5 gpc9910 (
      {stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[19]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc9911 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[20]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc9912 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[21]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[16],stage4_32[16]}
   );
   gpc615_5 gpc9913 (
      {stage3_32[41], stage3_32[42], stage3_32[43], stage3_32[44], stage3_32[45]},
      {stage3_33[22]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[17],stage4_32[17]}
   );
   gpc615_5 gpc9914 (
      {stage3_32[46], stage3_32[47], stage3_32[48], stage3_32[49], stage3_32[50]},
      {stage3_33[23]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[8],stage4_34[10],stage4_33[18],stage4_32[18]}
   );
   gpc215_4 gpc9915 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28]},
      {stage3_34[26]},
      {stage3_35[4], stage3_35[5]},
      {stage4_36[6],stage4_35[9],stage4_34[11],stage4_33[19]}
   );
   gpc606_5 gpc9916 (
      {stage3_33[29], stage3_33[30], stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[7],stage4_35[10],stage4_34[12],stage4_33[20]}
   );
   gpc606_5 gpc9917 (
      {stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38], stage3_33[39], stage3_33[40]},
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage4_37[1],stage4_36[8],stage4_35[11],stage4_34[13],stage4_33[21]}
   );
   gpc606_5 gpc9918 (
      {stage3_33[41], stage3_33[42], stage3_33[43], stage3_33[44], stage3_33[45], stage3_33[46]},
      {stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage4_37[2],stage4_36[9],stage4_35[12],stage4_34[14],stage4_33[22]}
   );
   gpc606_5 gpc9919 (
      {stage3_33[47], stage3_33[48], stage3_33[49], stage3_33[50], stage3_33[51], stage3_33[52]},
      {stage3_35[24], stage3_35[25], stage3_35[26], stage3_35[27], stage3_35[28], stage3_35[29]},
      {stage4_37[3],stage4_36[10],stage4_35[13],stage4_34[15],stage4_33[23]}
   );
   gpc615_5 gpc9920 (
      {stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage3_35[30]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage4_38[0],stage4_37[4],stage4_36[11],stage4_35[14],stage4_34[16]}
   );
   gpc606_5 gpc9921 (
      {stage3_35[31], stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[1],stage4_37[5],stage4_36[12],stage4_35[15]}
   );
   gpc615_5 gpc9922 (
      {stage3_35[37], stage3_35[38], stage3_35[39], stage3_35[40], stage3_35[41]},
      {stage3_36[6]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[2],stage4_37[6],stage4_36[13],stage4_35[16]}
   );
   gpc615_5 gpc9923 (
      {stage3_35[42], stage3_35[43], stage3_35[44], stage3_35[45], stage3_35[46]},
      {stage3_36[7]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[3],stage4_37[7],stage4_36[14],stage4_35[17]}
   );
   gpc615_5 gpc9924 (
      {stage3_35[47], stage3_35[48], stage3_35[49], stage3_35[50], stage3_35[51]},
      {stage3_36[8]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[4],stage4_37[8],stage4_36[15],stage4_35[18]}
   );
   gpc606_5 gpc9925 (
      {stage3_36[9], stage3_36[10], stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[4],stage4_38[5],stage4_37[9],stage4_36[16]}
   );
   gpc606_5 gpc9926 (
      {stage3_36[15], stage3_36[16], stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[5],stage4_38[6],stage4_37[10],stage4_36[17]}
   );
   gpc606_5 gpc9927 (
      {stage3_36[21], stage3_36[22], stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[6],stage4_38[7],stage4_37[11],stage4_36[18]}
   );
   gpc606_5 gpc9928 (
      {stage3_36[27], stage3_36[28], stage3_36[29], stage3_36[30], stage3_36[31], stage3_36[32]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[7],stage4_38[8],stage4_37[12],stage4_36[19]}
   );
   gpc606_5 gpc9929 (
      {stage3_36[33], stage3_36[34], stage3_36[35], stage3_36[36], stage3_36[37], stage3_36[38]},
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28], stage3_38[29]},
      {stage4_40[4],stage4_39[8],stage4_38[9],stage4_37[13],stage4_36[20]}
   );
   gpc606_5 gpc9930 (
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[5],stage4_39[9],stage4_38[10],stage4_37[14]}
   );
   gpc606_5 gpc9931 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], 1'b0},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[6],stage4_39[10],stage4_38[11],stage4_37[15]}
   );
   gpc615_5 gpc9932 (
      {stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33], stage3_38[34]},
      {stage3_39[12]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[2],stage4_40[7],stage4_39[11],stage4_38[12]}
   );
   gpc615_5 gpc9933 (
      {stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38], stage3_38[39]},
      {stage3_39[13]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[3],stage4_40[8],stage4_39[12],stage4_38[13]}
   );
   gpc615_5 gpc9934 (
      {stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43], stage3_38[44]},
      {stage3_39[14]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[4],stage4_40[9],stage4_39[13],stage4_38[14]}
   );
   gpc615_5 gpc9935 (
      {stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48], stage3_38[49]},
      {stage3_39[15]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[5],stage4_40[10],stage4_39[14],stage4_38[15]}
   );
   gpc615_5 gpc9936 (
      {stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53], stage3_38[54]},
      {stage3_39[16]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[6],stage4_40[11],stage4_39[15],stage4_38[16]}
   );
   gpc615_5 gpc9937 (
      {stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58], stage3_38[59]},
      {stage3_39[17]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[7],stage4_40[12],stage4_39[16],stage4_38[17]}
   );
   gpc207_4 gpc9938 (
      {stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22], stage3_39[23], stage3_39[24]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[6],stage4_41[8],stage4_40[13],stage4_39[17]}
   );
   gpc207_4 gpc9939 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[7],stage4_41[9],stage4_40[14],stage4_39[18]}
   );
   gpc207_4 gpc9940 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[8],stage4_41[10],stage4_40[15],stage4_39[19]}
   );
   gpc207_4 gpc9941 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[9],stage4_41[11],stage4_40[16],stage4_39[20]}
   );
   gpc207_4 gpc9942 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[8], stage3_41[9]},
      {stage4_42[10],stage4_41[12],stage4_40[17],stage4_39[21]}
   );
   gpc207_4 gpc9943 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57], stage3_39[58], stage3_39[59]},
      {stage3_41[10], stage3_41[11]},
      {stage4_42[11],stage4_41[13],stage4_40[18],stage4_39[22]}
   );
   gpc606_5 gpc9944 (
      {stage3_41[12], stage3_41[13], stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[12],stage4_41[14]}
   );
   gpc606_5 gpc9945 (
      {stage3_41[18], stage3_41[19], stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[13],stage4_41[15]}
   );
   gpc606_5 gpc9946 (
      {stage3_41[24], stage3_41[25], stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[14],stage4_41[16]}
   );
   gpc606_5 gpc9947 (
      {stage3_41[30], stage3_41[31], stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[15],stage4_41[17]}
   );
   gpc606_5 gpc9948 (
      {stage3_41[36], stage3_41[37], stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41]},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[16],stage4_41[18]}
   );
   gpc606_5 gpc9949 (
      {stage3_41[42], stage3_41[43], stage3_41[44], stage3_41[45], stage3_41[46], stage3_41[47]},
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[17],stage4_41[19]}
   );
   gpc606_5 gpc9950 (
      {stage3_41[48], stage3_41[49], stage3_41[50], stage3_41[51], stage3_41[52], stage3_41[53]},
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage4_45[6],stage4_44[6],stage4_43[6],stage4_42[18],stage4_41[20]}
   );
   gpc207_4 gpc9951 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[7],stage4_44[7],stage4_43[7],stage4_42[19]}
   );
   gpc207_4 gpc9952 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[8],stage4_44[8],stage4_43[8],stage4_42[20]}
   );
   gpc615_5 gpc9953 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18]},
      {stage3_43[42]},
      {stage3_44[4], stage3_44[5], stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[9],stage4_42[21]}
   );
   gpc615_5 gpc9954 (
      {stage3_42[19], stage3_42[20], stage3_42[21], stage3_42[22], stage3_42[23]},
      {stage3_43[43]},
      {stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[10],stage4_42[22]}
   );
   gpc615_5 gpc9955 (
      {stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27], stage3_42[28]},
      {stage3_43[44]},
      {stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21]},
      {stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[11],stage4_42[23]}
   );
   gpc615_5 gpc9956 (
      {stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_43[45]},
      {stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26], stage3_44[27]},
      {stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[12],stage4_42[24]}
   );
   gpc615_5 gpc9957 (
      {stage3_42[34], stage3_42[35], stage3_42[36], stage3_42[37], stage3_42[38]},
      {stage3_43[46]},
      {stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31], stage3_44[32], stage3_44[33]},
      {stage4_46[4],stage4_45[13],stage4_44[13],stage4_43[13],stage4_42[25]}
   );
   gpc615_5 gpc9958 (
      {stage3_42[39], stage3_42[40], stage3_42[41], stage3_42[42], stage3_42[43]},
      {stage3_43[47]},
      {stage3_44[34], stage3_44[35], stage3_44[36], stage3_44[37], stage3_44[38], stage3_44[39]},
      {stage4_46[5],stage4_45[14],stage4_44[14],stage4_43[14],stage4_42[26]}
   );
   gpc615_5 gpc9959 (
      {stage3_42[44], stage3_42[45], stage3_42[46], stage3_42[47], stage3_42[48]},
      {stage3_43[48]},
      {stage3_44[40], stage3_44[41], stage3_44[42], stage3_44[43], stage3_44[44], stage3_44[45]},
      {stage4_46[6],stage4_45[15],stage4_44[15],stage4_43[15],stage4_42[27]}
   );
   gpc615_5 gpc9960 (
      {stage3_42[49], stage3_42[50], stage3_42[51], stage3_42[52], stage3_42[53]},
      {stage3_43[49]},
      {stage3_44[46], stage3_44[47], stage3_44[48], stage3_44[49], stage3_44[50], stage3_44[51]},
      {stage4_46[7],stage4_45[16],stage4_44[16],stage4_43[16],stage4_42[28]}
   );
   gpc615_5 gpc9961 (
      {stage3_43[50], stage3_43[51], stage3_43[52], stage3_43[53], stage3_43[54]},
      {stage3_44[52]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[8],stage4_45[17],stage4_44[17],stage4_43[17]}
   );
   gpc1343_5 gpc9962 (
      {stage3_44[53], stage3_44[54], stage3_44[55]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[1],stage4_46[9],stage4_45[18],stage4_44[18]}
   );
   gpc1343_5 gpc9963 (
      {stage3_44[56], stage3_44[57], stage3_44[58]},
      {stage3_45[10], stage3_45[11], stage3_45[12], stage3_45[13]},
      {stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[1]},
      {stage4_48[1],stage4_47[2],stage4_46[10],stage4_45[19],stage4_44[19]}
   );
   gpc1343_5 gpc9964 (
      {stage3_44[59], stage3_44[60], stage3_44[61]},
      {stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_46[6], stage3_46[7], stage3_46[8]},
      {stage3_47[2]},
      {stage4_48[2],stage4_47[3],stage4_46[11],stage4_45[20],stage4_44[20]}
   );
   gpc623_5 gpc9965 (
      {stage3_44[62], stage3_44[63], stage3_44[64]},
      {stage3_45[18], stage3_45[19]},
      {stage3_46[9], stage3_46[10], stage3_46[11], stage3_46[12], stage3_46[13], stage3_46[14]},
      {stage4_48[3],stage4_47[4],stage4_46[12],stage4_45[21],stage4_44[21]}
   );
   gpc623_5 gpc9966 (
      {stage3_44[65], stage3_44[66], stage3_44[67]},
      {stage3_45[20], stage3_45[21]},
      {stage3_46[15], stage3_46[16], stage3_46[17], stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage4_48[4],stage4_47[5],stage4_46[13],stage4_45[22],stage4_44[22]}
   );
   gpc606_5 gpc9967 (
      {stage3_45[22], stage3_45[23], stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27]},
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8]},
      {stage4_49[0],stage4_48[5],stage4_47[6],stage4_46[14],stage4_45[23]}
   );
   gpc606_5 gpc9968 (
      {stage3_45[28], stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage4_49[1],stage4_48[6],stage4_47[7],stage4_46[15],stage4_45[24]}
   );
   gpc606_5 gpc9969 (
      {stage3_45[34], stage3_45[35], stage3_45[36], stage3_45[37], stage3_45[38], stage3_45[39]},
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage4_49[2],stage4_48[7],stage4_47[8],stage4_46[16],stage4_45[25]}
   );
   gpc615_5 gpc9970 (
      {stage3_46[21], stage3_46[22], stage3_46[23], stage3_46[24], stage3_46[25]},
      {stage3_47[21]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[3],stage4_48[8],stage4_47[9],stage4_46[17]}
   );
   gpc615_5 gpc9971 (
      {stage3_46[26], stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30]},
      {stage3_47[22]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[4],stage4_48[9],stage4_47[10],stage4_46[18]}
   );
   gpc615_5 gpc9972 (
      {stage3_46[31], stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35]},
      {stage3_47[23]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[5],stage4_48[10],stage4_47[11],stage4_46[19]}
   );
   gpc615_5 gpc9973 (
      {stage3_46[36], stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40]},
      {stage3_47[24]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[6],stage4_48[11],stage4_47[12],stage4_46[20]}
   );
   gpc615_5 gpc9974 (
      {stage3_46[41], stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45]},
      {stage3_47[25]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[7],stage4_48[12],stage4_47[13],stage4_46[21]}
   );
   gpc615_5 gpc9975 (
      {stage3_47[26], stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30]},
      {stage3_48[30]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[5],stage4_49[8],stage4_48[13],stage4_47[14]}
   );
   gpc615_5 gpc9976 (
      {stage3_47[31], stage3_47[32], stage3_47[33], stage3_47[34], stage3_47[35]},
      {stage3_48[31]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[6],stage4_49[9],stage4_48[14],stage4_47[15]}
   );
   gpc615_5 gpc9977 (
      {stage3_47[36], stage3_47[37], stage3_47[38], stage3_47[39], stage3_47[40]},
      {stage3_48[32]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[7],stage4_49[10],stage4_48[15],stage4_47[16]}
   );
   gpc615_5 gpc9978 (
      {stage3_47[41], stage3_47[42], stage3_47[43], stage3_47[44], stage3_47[45]},
      {stage3_48[33]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[8],stage4_49[11],stage4_48[16],stage4_47[17]}
   );
   gpc615_5 gpc9979 (
      {stage3_47[46], stage3_47[47], stage3_47[48], stage3_47[49], stage3_47[50]},
      {stage3_48[34]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[9],stage4_49[12],stage4_48[17],stage4_47[18]}
   );
   gpc615_5 gpc9980 (
      {stage3_47[51], stage3_47[52], stage3_47[53], stage3_47[54], stage3_47[55]},
      {stage3_48[35]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[10],stage4_49[13],stage4_48[18],stage4_47[19]}
   );
   gpc615_5 gpc9981 (
      {stage3_47[56], stage3_47[57], stage3_47[58], stage3_47[59], stage3_47[60]},
      {stage3_48[36]},
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage4_51[6],stage4_50[11],stage4_49[14],stage4_48[19],stage4_47[20]}
   );
   gpc615_5 gpc9982 (
      {stage3_47[61], stage3_47[62], stage3_47[63], stage3_47[64], stage3_47[65]},
      {1'b0},
      {stage3_49[42], stage3_49[43], stage3_49[44], stage3_49[45], stage3_49[46], stage3_49[47]},
      {stage4_51[7],stage4_50[12],stage4_49[15],stage4_48[20],stage4_47[21]}
   );
   gpc615_5 gpc9983 (
      {stage3_47[66], stage3_47[67], stage3_47[68], stage3_47[69], stage3_47[70]},
      {1'b0},
      {stage3_49[48], stage3_49[49], stage3_49[50], stage3_49[51], stage3_49[52], stage3_49[53]},
      {stage4_51[8],stage4_50[13],stage4_49[16],stage4_48[21],stage4_47[22]}
   );
   gpc117_4 gpc9984 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[0]},
      {stage3_52[0]},
      {stage4_53[0],stage4_52[0],stage4_51[9],stage4_50[14]}
   );
   gpc117_4 gpc9985 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[1]},
      {stage3_52[1]},
      {stage4_53[1],stage4_52[1],stage4_51[10],stage4_50[15]}
   );
   gpc117_4 gpc9986 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18], stage3_50[19], stage3_50[20]},
      {stage3_51[2]},
      {stage3_52[2]},
      {stage4_53[2],stage4_52[2],stage4_51[11],stage4_50[16]}
   );
   gpc117_4 gpc9987 (
      {stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27]},
      {stage3_51[3]},
      {stage3_52[3]},
      {stage4_53[3],stage4_52[3],stage4_51[12],stage4_50[17]}
   );
   gpc117_4 gpc9988 (
      {stage3_50[28], stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33], stage3_50[34]},
      {stage3_51[4]},
      {stage3_52[4]},
      {stage4_53[4],stage4_52[4],stage4_51[13],stage4_50[18]}
   );
   gpc117_4 gpc9989 (
      {stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38], stage3_50[39], stage3_50[40], stage3_50[41]},
      {stage3_51[5]},
      {stage3_52[5]},
      {stage4_53[5],stage4_52[5],stage4_51[14],stage4_50[19]}
   );
   gpc117_4 gpc9990 (
      {stage3_50[42], stage3_50[43], stage3_50[44], stage3_50[45], stage3_50[46], stage3_50[47], stage3_50[48]},
      {stage3_51[6]},
      {stage3_52[6]},
      {stage4_53[6],stage4_52[6],stage4_51[15],stage4_50[20]}
   );
   gpc117_4 gpc9991 (
      {stage3_50[49], stage3_50[50], stage3_50[51], stage3_50[52], stage3_50[53], stage3_50[54], stage3_50[55]},
      {stage3_51[7]},
      {stage3_52[7]},
      {stage4_53[7],stage4_52[7],stage4_51[16],stage4_50[21]}
   );
   gpc117_4 gpc9992 (
      {stage3_50[56], stage3_50[57], stage3_50[58], stage3_50[59], stage3_50[60], stage3_50[61], stage3_50[62]},
      {stage3_51[8]},
      {stage3_52[8]},
      {stage4_53[8],stage4_52[8],stage4_51[17],stage4_50[22]}
   );
   gpc2135_5 gpc9993 (
      {stage3_51[9], stage3_51[10], stage3_51[11], stage3_51[12], stage3_51[13]},
      {stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[0],stage4_53[9],stage4_52[9],stage4_51[18]}
   );
   gpc2135_5 gpc9994 (
      {stage3_51[14], stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18]},
      {stage3_52[12], stage3_52[13], stage3_52[14]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[1],stage4_53[10],stage4_52[10],stage4_51[19]}
   );
   gpc2135_5 gpc9995 (
      {stage3_51[19], stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23]},
      {stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[2],stage4_53[11],stage4_52[11],stage4_51[20]}
   );
   gpc2135_5 gpc9996 (
      {stage3_51[24], stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28]},
      {stage3_52[18], stage3_52[19], stage3_52[20]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[3],stage4_53[12],stage4_52[12],stage4_51[21]}
   );
   gpc2135_5 gpc9997 (
      {stage3_51[29], stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33]},
      {stage3_52[21], stage3_52[22], stage3_52[23]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[4],stage4_53[13],stage4_52[13],stage4_51[22]}
   );
   gpc2135_5 gpc9998 (
      {stage3_51[34], stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38]},
      {stage3_52[24], stage3_52[25], stage3_52[26]},
      {stage3_53[5]},
      {stage3_54[10], stage3_54[11]},
      {stage4_55[5],stage4_54[5],stage4_53[14],stage4_52[14],stage4_51[23]}
   );
   gpc2135_5 gpc9999 (
      {stage3_51[39], stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43]},
      {stage3_52[27], stage3_52[28], stage3_52[29]},
      {stage3_53[6]},
      {stage3_54[12], stage3_54[13]},
      {stage4_55[6],stage4_54[6],stage4_53[15],stage4_52[15],stage4_51[24]}
   );
   gpc2135_5 gpc10000 (
      {stage3_51[44], stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48]},
      {stage3_52[30], stage3_52[31], stage3_52[32]},
      {stage3_53[7]},
      {stage3_54[14], stage3_54[15]},
      {stage4_55[7],stage4_54[7],stage4_53[16],stage4_52[16],stage4_51[25]}
   );
   gpc2135_5 gpc10001 (
      {stage3_51[49], stage3_51[50], stage3_51[51], stage3_51[52], stage3_51[53]},
      {stage3_52[33], stage3_52[34], stage3_52[35]},
      {stage3_53[8]},
      {stage3_54[16], stage3_54[17]},
      {stage4_55[8],stage4_54[8],stage4_53[17],stage4_52[17],stage4_51[26]}
   );
   gpc606_5 gpc10002 (
      {stage3_52[36], stage3_52[37], stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41]},
      {stage3_54[18], stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage4_56[0],stage4_55[9],stage4_54[9],stage4_53[18],stage4_52[18]}
   );
   gpc606_5 gpc10003 (
      {stage3_52[42], stage3_52[43], stage3_52[44], stage3_52[45], stage3_52[46], stage3_52[47]},
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28], stage3_54[29]},
      {stage4_56[1],stage4_55[10],stage4_54[10],stage4_53[19],stage4_52[19]}
   );
   gpc606_5 gpc10004 (
      {stage3_52[48], stage3_52[49], stage3_52[50], stage3_52[51], stage3_52[52], stage3_52[53]},
      {stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33], stage3_54[34], stage3_54[35]},
      {stage4_56[2],stage4_55[11],stage4_54[11],stage4_53[20],stage4_52[20]}
   );
   gpc1415_5 gpc10005 (
      {stage3_53[9], stage3_53[10], stage3_53[11], stage3_53[12], stage3_53[13]},
      {stage3_54[36]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[3],stage4_55[12],stage4_54[12],stage4_53[21]}
   );
   gpc1415_5 gpc10006 (
      {stage3_53[14], stage3_53[15], stage3_53[16], stage3_53[17], stage3_53[18]},
      {stage3_54[37]},
      {stage3_55[4], stage3_55[5], stage3_55[6], stage3_55[7]},
      {stage3_56[1]},
      {stage4_57[1],stage4_56[4],stage4_55[13],stage4_54[13],stage4_53[22]}
   );
   gpc1415_5 gpc10007 (
      {stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22], stage3_53[23]},
      {stage3_54[38]},
      {stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage3_56[2]},
      {stage4_57[2],stage4_56[5],stage4_55[14],stage4_54[14],stage4_53[23]}
   );
   gpc1415_5 gpc10008 (
      {stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_54[39]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15]},
      {stage3_56[3]},
      {stage4_57[3],stage4_56[6],stage4_55[15],stage4_54[15],stage4_53[24]}
   );
   gpc606_5 gpc10009 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[16], stage3_55[17], stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21]},
      {stage4_57[4],stage4_56[7],stage4_55[16],stage4_54[16],stage4_53[25]}
   );
   gpc606_5 gpc10010 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39], stage3_53[40]},
      {stage3_55[22], stage3_55[23], stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27]},
      {stage4_57[5],stage4_56[8],stage4_55[17],stage4_54[17],stage4_53[26]}
   );
   gpc606_5 gpc10011 (
      {stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44], stage3_53[45], stage3_53[46]},
      {stage3_55[28], stage3_55[29], stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33]},
      {stage4_57[6],stage4_56[9],stage4_55[18],stage4_54[18],stage4_53[27]}
   );
   gpc606_5 gpc10012 (
      {stage3_53[47], stage3_53[48], stage3_53[49], stage3_53[50], stage3_53[51], stage3_53[52]},
      {stage3_55[34], stage3_55[35], stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39]},
      {stage4_57[7],stage4_56[10],stage4_55[19],stage4_54[19],stage4_53[28]}
   );
   gpc207_4 gpc10013 (
      {stage3_54[40], stage3_54[41], stage3_54[42], stage3_54[43], stage3_54[44], stage3_54[45], stage3_54[46]},
      {stage3_56[4], stage3_56[5]},
      {stage4_57[8],stage4_56[11],stage4_55[20],stage4_54[20]}
   );
   gpc207_4 gpc10014 (
      {stage3_54[47], stage3_54[48], stage3_54[49], stage3_54[50], stage3_54[51], stage3_54[52], stage3_54[53]},
      {stage3_56[6], stage3_56[7]},
      {stage4_57[9],stage4_56[12],stage4_55[21],stage4_54[21]}
   );
   gpc606_5 gpc10015 (
      {stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12], stage3_56[13]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[0],stage4_58[0],stage4_57[10],stage4_56[13]}
   );
   gpc606_5 gpc10016 (
      {stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18], stage3_56[19]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[1],stage4_58[1],stage4_57[11],stage4_56[14]}
   );
   gpc606_5 gpc10017 (
      {stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23], stage3_56[24], stage3_56[25]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[2],stage4_58[2],stage4_57[12],stage4_56[15]}
   );
   gpc1163_5 gpc10018 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[3],stage4_59[3],stage4_58[3],stage4_57[13]}
   );
   gpc1163_5 gpc10019 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[4],stage4_59[4],stage4_58[4],stage4_57[14]}
   );
   gpc1163_5 gpc10020 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[5],stage4_59[5],stage4_58[5],stage4_57[15]}
   );
   gpc606_5 gpc10021 (
      {stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7], stage3_59[8]},
      {stage4_61[3],stage4_60[6],stage4_59[6],stage4_58[6],stage4_57[16]}
   );
   gpc606_5 gpc10022 (
      {stage3_57[15], stage3_57[16], stage3_57[17], stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[4],stage4_60[7],stage4_59[7],stage4_58[7],stage4_57[17]}
   );
   gpc606_5 gpc10023 (
      {stage3_57[21], stage3_57[22], stage3_57[23], stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[5],stage4_60[8],stage4_59[8],stage4_58[8],stage4_57[18]}
   );
   gpc606_5 gpc10024 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[6],stage4_60[9],stage4_59[9],stage4_58[9],stage4_57[19]}
   );
   gpc606_5 gpc10025 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[7],stage4_60[10],stage4_59[10],stage4_58[10],stage4_57[20]}
   );
   gpc606_5 gpc10026 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43], stage3_57[44]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[8],stage4_60[11],stage4_59[11],stage4_58[11],stage4_57[21]}
   );
   gpc606_5 gpc10027 (
      {stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48], stage3_57[49], stage3_57[50]},
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43], stage3_59[44]},
      {stage4_61[9],stage4_60[12],stage4_59[12],stage4_58[12],stage4_57[22]}
   );
   gpc1406_5 gpc10028 (
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_60[3], stage3_60[4], stage3_60[5], stage3_60[6]},
      {stage3_61[0]},
      {stage4_62[0],stage4_61[10],stage4_60[13],stage4_59[13],stage4_58[13]}
   );
   gpc606_5 gpc10029 (
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10], stage3_60[11], stage3_60[12]},
      {stage4_62[1],stage4_61[11],stage4_60[14],stage4_59[14],stage4_58[14]}
   );
   gpc1406_5 gpc10030 (
      {stage3_60[13], stage3_60[14], stage3_60[15], stage3_60[16], stage3_60[17], stage3_60[18]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0]},
      {stage4_64[0],stage4_63[0],stage4_62[2],stage4_61[12],stage4_60[15]}
   );
   gpc606_5 gpc10031 (
      {stage3_60[19], stage3_60[20], stage3_60[21], stage3_60[22], stage3_60[23], stage3_60[24]},
      {stage3_62[4], stage3_62[5], stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9]},
      {stage4_64[1],stage4_63[1],stage4_62[3],stage4_61[13],stage4_60[16]}
   );
   gpc606_5 gpc10032 (
      {stage3_60[25], stage3_60[26], stage3_60[27], stage3_60[28], stage3_60[29], stage3_60[30]},
      {stage3_62[10], stage3_62[11], stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15]},
      {stage4_64[2],stage4_63[2],stage4_62[4],stage4_61[14],stage4_60[17]}
   );
   gpc606_5 gpc10033 (
      {stage3_60[31], stage3_60[32], stage3_60[33], stage3_60[34], stage3_60[35], stage3_60[36]},
      {stage3_62[16], stage3_62[17], stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21]},
      {stage4_64[3],stage4_63[3],stage4_62[5],stage4_61[15],stage4_60[18]}
   );
   gpc606_5 gpc10034 (
      {stage3_60[37], stage3_60[38], stage3_60[39], stage3_60[40], stage3_60[41], stage3_60[42]},
      {stage3_62[22], stage3_62[23], stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27]},
      {stage4_64[4],stage4_63[4],stage4_62[6],stage4_61[16],stage4_60[19]}
   );
   gpc606_5 gpc10035 (
      {stage3_60[43], stage3_60[44], stage3_60[45], stage3_60[46], stage3_60[47], stage3_60[48]},
      {stage3_62[28], stage3_62[29], stage3_62[30], stage3_62[31], stage3_62[32], stage3_62[33]},
      {stage4_64[5],stage4_63[5],stage4_62[7],stage4_61[17],stage4_60[20]}
   );
   gpc606_5 gpc10036 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5], stage3_61[6]},
      {stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6]},
      {stage4_65[0],stage4_64[6],stage4_63[6],stage4_62[8],stage4_61[18]}
   );
   gpc606_5 gpc10037 (
      {stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11], stage3_61[12]},
      {stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11], stage3_63[12]},
      {stage4_65[1],stage4_64[7],stage4_63[7],stage4_62[9],stage4_61[19]}
   );
   gpc606_5 gpc10038 (
      {stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17], stage3_61[18]},
      {stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17], stage3_63[18]},
      {stage4_65[2],stage4_64[8],stage4_63[8],stage4_62[10],stage4_61[20]}
   );
   gpc606_5 gpc10039 (
      {stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23], stage3_61[24]},
      {stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23], stage3_63[24]},
      {stage4_65[3],stage4_64[9],stage4_63[9],stage4_62[11],stage4_61[21]}
   );
   gpc606_5 gpc10040 (
      {stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29], stage3_61[30]},
      {stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29], stage3_63[30]},
      {stage4_65[4],stage4_64[10],stage4_63[10],stage4_62[12],stage4_61[22]}
   );
   gpc606_5 gpc10041 (
      {stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35], stage3_61[36]},
      {stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35], stage3_63[36]},
      {stage4_65[5],stage4_64[11],stage4_63[11],stage4_62[13],stage4_61[23]}
   );
   gpc606_5 gpc10042 (
      {stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41], stage3_61[42]},
      {stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41], stage3_63[42]},
      {stage4_65[6],stage4_64[12],stage4_63[12],stage4_62[14],stage4_61[24]}
   );
   gpc606_5 gpc10043 (
      {stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47], stage3_61[48]},
      {stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47], stage3_63[48]},
      {stage4_65[7],stage4_64[13],stage4_63[13],stage4_62[15],stage4_61[25]}
   );
   gpc606_5 gpc10044 (
      {stage3_61[49], stage3_61[50], stage3_61[51], stage3_61[52], stage3_61[53], stage3_61[54]},
      {stage3_63[49], stage3_63[50], stage3_63[51], stage3_63[52], stage3_63[53], stage3_63[54]},
      {stage4_65[8],stage4_64[14],stage4_63[14],stage4_62[16],stage4_61[26]}
   );
   gpc606_5 gpc10045 (
      {stage3_63[55], stage3_63[56], stage3_63[57], stage3_63[58], stage3_63[59], stage3_63[60]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[9],stage4_64[15],stage4_63[15]}
   );
   gpc606_5 gpc10046 (
      {stage3_63[61], stage3_63[62], stage3_63[63], stage3_63[64], stage3_63[65], stage3_63[66]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[1],stage4_65[10],stage4_64[16],stage4_63[16]}
   );
   gpc606_5 gpc10047 (
      {stage3_63[67], stage3_63[68], stage3_63[69], stage3_63[70], stage3_63[71], 1'b0},
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage4_67[2],stage4_66[2],stage4_65[11],stage4_64[17],stage4_63[17]}
   );
   gpc1163_5 gpc10048 (
      {stage3_64[0], stage3_64[1], stage3_64[2]},
      {stage3_65[18], stage3_65[19], stage3_65[20], stage3_65[21], stage3_65[22], stage3_65[23]},
      {stage3_66[0]},
      {stage3_67[0]},
      {stage4_68[0],stage4_67[3],stage4_66[3],stage4_65[12],stage4_64[18]}
   );
   gpc606_5 gpc10049 (
      {stage3_64[3], stage3_64[4], stage3_64[5], stage3_64[6], stage3_64[7], stage3_64[8]},
      {stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5], stage3_66[6]},
      {stage4_68[1],stage4_67[4],stage4_66[4],stage4_65[13],stage4_64[19]}
   );
   gpc606_5 gpc10050 (
      {stage3_64[9], stage3_64[10], stage3_64[11], stage3_64[12], stage3_64[13], stage3_64[14]},
      {stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11], stage3_66[12]},
      {stage4_68[2],stage4_67[5],stage4_66[5],stage4_65[14],stage4_64[20]}
   );
   gpc606_5 gpc10051 (
      {stage3_64[15], stage3_64[16], stage3_64[17], stage3_64[18], stage3_64[19], stage3_64[20]},
      {stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17], stage3_66[18]},
      {stage4_68[3],stage4_67[6],stage4_66[6],stage4_65[15],stage4_64[21]}
   );
   gpc606_5 gpc10052 (
      {stage3_64[21], stage3_64[22], stage3_64[23], stage3_64[24], stage3_64[25], stage3_64[26]},
      {stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23], stage3_66[24]},
      {stage4_68[4],stage4_67[7],stage4_66[7],stage4_65[16],stage4_64[22]}
   );
   gpc606_5 gpc10053 (
      {stage3_64[27], stage3_64[28], stage3_64[29], stage3_64[30], stage3_64[31], stage3_64[32]},
      {stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29], stage3_66[30]},
      {stage4_68[5],stage4_67[8],stage4_66[8],stage4_65[17],stage4_64[23]}
   );
   gpc606_5 gpc10054 (
      {stage3_64[33], stage3_64[34], stage3_64[35], stage3_64[36], stage3_64[37], stage3_64[38]},
      {stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35], stage3_66[36]},
      {stage4_68[6],stage4_67[9],stage4_66[9],stage4_65[18],stage4_64[24]}
   );
   gpc606_5 gpc10055 (
      {stage3_64[39], stage3_64[40], stage3_64[41], stage3_64[42], stage3_64[43], stage3_64[44]},
      {stage3_66[37], stage3_66[38], stage3_66[39], stage3_66[40], stage3_66[41], stage3_66[42]},
      {stage4_68[7],stage4_67[10],stage4_66[10],stage4_65[19],stage4_64[25]}
   );
   gpc606_5 gpc10056 (
      {stage3_64[45], stage3_64[46], stage3_64[47], stage3_64[48], stage3_64[49], stage3_64[50]},
      {stage3_66[43], stage3_66[44], stage3_66[45], stage3_66[46], stage3_66[47], stage3_66[48]},
      {stage4_68[8],stage4_67[11],stage4_66[11],stage4_65[20],stage4_64[26]}
   );
   gpc606_5 gpc10057 (
      {stage3_65[24], stage3_65[25], stage3_65[26], stage3_65[27], stage3_65[28], stage3_65[29]},
      {stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5], stage3_67[6]},
      {stage4_69[0],stage4_68[9],stage4_67[12],stage4_66[12],stage4_65[21]}
   );
   gpc606_5 gpc10058 (
      {stage3_65[30], stage3_65[31], stage3_65[32], 1'b0, 1'b0, 1'b0},
      {stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11], stage3_67[12]},
      {stage4_69[1],stage4_68[10],stage4_67[13],stage4_66[13],stage4_65[22]}
   );
   gpc606_5 gpc10059 (
      {stage3_66[49], stage3_66[50], stage3_66[51], stage3_66[52], stage3_66[53], 1'b0},
      {stage3_68[0], stage3_68[1], stage3_68[2], stage3_68[3], stage3_68[4], 1'b0},
      {stage4_70[0],stage4_69[2],stage4_68[11],stage4_67[14],stage4_66[14]}
   );
   gpc1_1 gpc10060 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc10061 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc10062 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc10063 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc10064 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc10065 (
      {stage3_1[24]},
      {stage4_1[5]}
   );
   gpc1_1 gpc10066 (
      {stage3_1[25]},
      {stage4_1[6]}
   );
   gpc1_1 gpc10067 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc10068 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc10069 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc10070 (
      {stage3_3[39]},
      {stage4_3[9]}
   );
   gpc1_1 gpc10071 (
      {stage3_3[40]},
      {stage4_3[10]}
   );
   gpc1_1 gpc10072 (
      {stage3_3[41]},
      {stage4_3[11]}
   );
   gpc1_1 gpc10073 (
      {stage3_3[42]},
      {stage4_3[12]}
   );
   gpc1_1 gpc10074 (
      {stage3_3[43]},
      {stage4_3[13]}
   );
   gpc1_1 gpc10075 (
      {stage3_3[44]},
      {stage4_3[14]}
   );
   gpc1_1 gpc10076 (
      {stage3_3[45]},
      {stage4_3[15]}
   );
   gpc1_1 gpc10077 (
      {stage3_3[46]},
      {stage4_3[16]}
   );
   gpc1_1 gpc10078 (
      {stage3_3[47]},
      {stage4_3[17]}
   );
   gpc1_1 gpc10079 (
      {stage3_3[48]},
      {stage4_3[18]}
   );
   gpc1_1 gpc10080 (
      {stage3_3[49]},
      {stage4_3[19]}
   );
   gpc1_1 gpc10081 (
      {stage3_3[50]},
      {stage4_3[20]}
   );
   gpc1_1 gpc10082 (
      {stage3_3[51]},
      {stage4_3[21]}
   );
   gpc1_1 gpc10083 (
      {stage3_4[51]},
      {stage4_4[16]}
   );
   gpc1_1 gpc10084 (
      {stage3_4[52]},
      {stage4_4[17]}
   );
   gpc1_1 gpc10085 (
      {stage3_4[53]},
      {stage4_4[18]}
   );
   gpc1_1 gpc10086 (
      {stage3_4[54]},
      {stage4_4[19]}
   );
   gpc1_1 gpc10087 (
      {stage3_4[55]},
      {stage4_4[20]}
   );
   gpc1_1 gpc10088 (
      {stage3_4[56]},
      {stage4_4[21]}
   );
   gpc1_1 gpc10089 (
      {stage3_4[57]},
      {stage4_4[22]}
   );
   gpc1_1 gpc10090 (
      {stage3_4[58]},
      {stage4_4[23]}
   );
   gpc1_1 gpc10091 (
      {stage3_4[59]},
      {stage4_4[24]}
   );
   gpc1_1 gpc10092 (
      {stage3_5[24]},
      {stage4_5[16]}
   );
   gpc1_1 gpc10093 (
      {stage3_5[25]},
      {stage4_5[17]}
   );
   gpc1_1 gpc10094 (
      {stage3_5[26]},
      {stage4_5[18]}
   );
   gpc1_1 gpc10095 (
      {stage3_5[27]},
      {stage4_5[19]}
   );
   gpc1_1 gpc10096 (
      {stage3_5[28]},
      {stage4_5[20]}
   );
   gpc1_1 gpc10097 (
      {stage3_5[29]},
      {stage4_5[21]}
   );
   gpc1_1 gpc10098 (
      {stage3_5[30]},
      {stage4_5[22]}
   );
   gpc1_1 gpc10099 (
      {stage3_5[31]},
      {stage4_5[23]}
   );
   gpc1_1 gpc10100 (
      {stage3_5[32]},
      {stage4_5[24]}
   );
   gpc1_1 gpc10101 (
      {stage3_5[33]},
      {stage4_5[25]}
   );
   gpc1_1 gpc10102 (
      {stage3_5[34]},
      {stage4_5[26]}
   );
   gpc1_1 gpc10103 (
      {stage3_5[35]},
      {stage4_5[27]}
   );
   gpc1_1 gpc10104 (
      {stage3_5[36]},
      {stage4_5[28]}
   );
   gpc1_1 gpc10105 (
      {stage3_5[37]},
      {stage4_5[29]}
   );
   gpc1_1 gpc10106 (
      {stage3_5[38]},
      {stage4_5[30]}
   );
   gpc1_1 gpc10107 (
      {stage3_5[39]},
      {stage4_5[31]}
   );
   gpc1_1 gpc10108 (
      {stage3_5[40]},
      {stage4_5[32]}
   );
   gpc1_1 gpc10109 (
      {stage3_5[41]},
      {stage4_5[33]}
   );
   gpc1_1 gpc10110 (
      {stage3_5[42]},
      {stage4_5[34]}
   );
   gpc1_1 gpc10111 (
      {stage3_5[43]},
      {stage4_5[35]}
   );
   gpc1_1 gpc10112 (
      {stage3_5[44]},
      {stage4_5[36]}
   );
   gpc1_1 gpc10113 (
      {stage3_5[45]},
      {stage4_5[37]}
   );
   gpc1_1 gpc10114 (
      {stage3_5[46]},
      {stage4_5[38]}
   );
   gpc1_1 gpc10115 (
      {stage3_5[47]},
      {stage4_5[39]}
   );
   gpc1_1 gpc10116 (
      {stage3_5[48]},
      {stage4_5[40]}
   );
   gpc1_1 gpc10117 (
      {stage3_5[49]},
      {stage4_5[41]}
   );
   gpc1_1 gpc10118 (
      {stage3_5[50]},
      {stage4_5[42]}
   );
   gpc1_1 gpc10119 (
      {stage3_5[51]},
      {stage4_5[43]}
   );
   gpc1_1 gpc10120 (
      {stage3_5[52]},
      {stage4_5[44]}
   );
   gpc1_1 gpc10121 (
      {stage3_5[53]},
      {stage4_5[45]}
   );
   gpc1_1 gpc10122 (
      {stage3_5[54]},
      {stage4_5[46]}
   );
   gpc1_1 gpc10123 (
      {stage3_6[62]},
      {stage4_6[16]}
   );
   gpc1_1 gpc10124 (
      {stage3_6[63]},
      {stage4_6[17]}
   );
   gpc1_1 gpc10125 (
      {stage3_6[64]},
      {stage4_6[18]}
   );
   gpc1_1 gpc10126 (
      {stage3_6[65]},
      {stage4_6[19]}
   );
   gpc1_1 gpc10127 (
      {stage3_6[66]},
      {stage4_6[20]}
   );
   gpc1_1 gpc10128 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc10129 (
      {stage3_7[36]},
      {stage4_7[21]}
   );
   gpc1_1 gpc10130 (
      {stage3_7[37]},
      {stage4_7[22]}
   );
   gpc1_1 gpc10131 (
      {stage3_7[38]},
      {stage4_7[23]}
   );
   gpc1_1 gpc10132 (
      {stage3_7[39]},
      {stage4_7[24]}
   );
   gpc1_1 gpc10133 (
      {stage3_7[40]},
      {stage4_7[25]}
   );
   gpc1_1 gpc10134 (
      {stage3_7[41]},
      {stage4_7[26]}
   );
   gpc1_1 gpc10135 (
      {stage3_7[42]},
      {stage4_7[27]}
   );
   gpc1_1 gpc10136 (
      {stage3_7[43]},
      {stage4_7[28]}
   );
   gpc1_1 gpc10137 (
      {stage3_7[44]},
      {stage4_7[29]}
   );
   gpc1_1 gpc10138 (
      {stage3_7[45]},
      {stage4_7[30]}
   );
   gpc1_1 gpc10139 (
      {stage3_7[46]},
      {stage4_7[31]}
   );
   gpc1_1 gpc10140 (
      {stage3_7[47]},
      {stage4_7[32]}
   );
   gpc1_1 gpc10141 (
      {stage3_7[48]},
      {stage4_7[33]}
   );
   gpc1_1 gpc10142 (
      {stage3_7[49]},
      {stage4_7[34]}
   );
   gpc1_1 gpc10143 (
      {stage3_7[50]},
      {stage4_7[35]}
   );
   gpc1_1 gpc10144 (
      {stage3_7[51]},
      {stage4_7[36]}
   );
   gpc1_1 gpc10145 (
      {stage3_7[52]},
      {stage4_7[37]}
   );
   gpc1_1 gpc10146 (
      {stage3_7[53]},
      {stage4_7[38]}
   );
   gpc1_1 gpc10147 (
      {stage3_7[54]},
      {stage4_7[39]}
   );
   gpc1_1 gpc10148 (
      {stage3_8[29]},
      {stage4_8[17]}
   );
   gpc1_1 gpc10149 (
      {stage3_8[30]},
      {stage4_8[18]}
   );
   gpc1_1 gpc10150 (
      {stage3_8[31]},
      {stage4_8[19]}
   );
   gpc1_1 gpc10151 (
      {stage3_8[32]},
      {stage4_8[20]}
   );
   gpc1_1 gpc10152 (
      {stage3_8[33]},
      {stage4_8[21]}
   );
   gpc1_1 gpc10153 (
      {stage3_8[34]},
      {stage4_8[22]}
   );
   gpc1_1 gpc10154 (
      {stage3_8[35]},
      {stage4_8[23]}
   );
   gpc1_1 gpc10155 (
      {stage3_8[36]},
      {stage4_8[24]}
   );
   gpc1_1 gpc10156 (
      {stage3_8[37]},
      {stage4_8[25]}
   );
   gpc1_1 gpc10157 (
      {stage3_8[38]},
      {stage4_8[26]}
   );
   gpc1_1 gpc10158 (
      {stage3_8[39]},
      {stage4_8[27]}
   );
   gpc1_1 gpc10159 (
      {stage3_8[40]},
      {stage4_8[28]}
   );
   gpc1_1 gpc10160 (
      {stage3_8[41]},
      {stage4_8[29]}
   );
   gpc1_1 gpc10161 (
      {stage3_8[42]},
      {stage4_8[30]}
   );
   gpc1_1 gpc10162 (
      {stage3_8[43]},
      {stage4_8[31]}
   );
   gpc1_1 gpc10163 (
      {stage3_8[44]},
      {stage4_8[32]}
   );
   gpc1_1 gpc10164 (
      {stage3_8[45]},
      {stage4_8[33]}
   );
   gpc1_1 gpc10165 (
      {stage3_8[46]},
      {stage4_8[34]}
   );
   gpc1_1 gpc10166 (
      {stage3_10[65]},
      {stage4_10[26]}
   );
   gpc1_1 gpc10167 (
      {stage3_10[66]},
      {stage4_10[27]}
   );
   gpc1_1 gpc10168 (
      {stage3_10[67]},
      {stage4_10[28]}
   );
   gpc1_1 gpc10169 (
      {stage3_11[52]},
      {stage4_11[25]}
   );
   gpc1_1 gpc10170 (
      {stage3_11[53]},
      {stage4_11[26]}
   );
   gpc1_1 gpc10171 (
      {stage3_11[54]},
      {stage4_11[27]}
   );
   gpc1_1 gpc10172 (
      {stage3_11[55]},
      {stage4_11[28]}
   );
   gpc1_1 gpc10173 (
      {stage3_11[56]},
      {stage4_11[29]}
   );
   gpc1_1 gpc10174 (
      {stage3_11[57]},
      {stage4_11[30]}
   );
   gpc1_1 gpc10175 (
      {stage3_11[58]},
      {stage4_11[31]}
   );
   gpc1_1 gpc10176 (
      {stage3_11[59]},
      {stage4_11[32]}
   );
   gpc1_1 gpc10177 (
      {stage3_11[60]},
      {stage4_11[33]}
   );
   gpc1_1 gpc10178 (
      {stage3_13[43]},
      {stage4_13[24]}
   );
   gpc1_1 gpc10179 (
      {stage3_13[44]},
      {stage4_13[25]}
   );
   gpc1_1 gpc10180 (
      {stage3_13[45]},
      {stage4_13[26]}
   );
   gpc1_1 gpc10181 (
      {stage3_13[46]},
      {stage4_13[27]}
   );
   gpc1_1 gpc10182 (
      {stage3_14[31]},
      {stage4_14[26]}
   );
   gpc1_1 gpc10183 (
      {stage3_14[32]},
      {stage4_14[27]}
   );
   gpc1_1 gpc10184 (
      {stage3_14[33]},
      {stage4_14[28]}
   );
   gpc1_1 gpc10185 (
      {stage3_14[34]},
      {stage4_14[29]}
   );
   gpc1_1 gpc10186 (
      {stage3_15[45]},
      {stage4_15[17]}
   );
   gpc1_1 gpc10187 (
      {stage3_15[46]},
      {stage4_15[18]}
   );
   gpc1_1 gpc10188 (
      {stage3_15[47]},
      {stage4_15[19]}
   );
   gpc1_1 gpc10189 (
      {stage3_15[48]},
      {stage4_15[20]}
   );
   gpc1_1 gpc10190 (
      {stage3_15[49]},
      {stage4_15[21]}
   );
   gpc1_1 gpc10191 (
      {stage3_15[50]},
      {stage4_15[22]}
   );
   gpc1_1 gpc10192 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc10193 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc10194 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc10195 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc10196 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc10197 (
      {stage3_16[45]},
      {stage4_16[19]}
   );
   gpc1_1 gpc10198 (
      {stage3_16[46]},
      {stage4_16[20]}
   );
   gpc1_1 gpc10199 (
      {stage3_16[47]},
      {stage4_16[21]}
   );
   gpc1_1 gpc10200 (
      {stage3_16[48]},
      {stage4_16[22]}
   );
   gpc1_1 gpc10201 (
      {stage3_16[49]},
      {stage4_16[23]}
   );
   gpc1_1 gpc10202 (
      {stage3_16[50]},
      {stage4_16[24]}
   );
   gpc1_1 gpc10203 (
      {stage3_16[51]},
      {stage4_16[25]}
   );
   gpc1_1 gpc10204 (
      {stage3_16[52]},
      {stage4_16[26]}
   );
   gpc1_1 gpc10205 (
      {stage3_16[53]},
      {stage4_16[27]}
   );
   gpc1_1 gpc10206 (
      {stage3_16[54]},
      {stage4_16[28]}
   );
   gpc1_1 gpc10207 (
      {stage3_16[55]},
      {stage4_16[29]}
   );
   gpc1_1 gpc10208 (
      {stage3_16[56]},
      {stage4_16[30]}
   );
   gpc1_1 gpc10209 (
      {stage3_16[57]},
      {stage4_16[31]}
   );
   gpc1_1 gpc10210 (
      {stage3_16[58]},
      {stage4_16[32]}
   );
   gpc1_1 gpc10211 (
      {stage3_17[36]},
      {stage4_17[15]}
   );
   gpc1_1 gpc10212 (
      {stage3_17[37]},
      {stage4_17[16]}
   );
   gpc1_1 gpc10213 (
      {stage3_17[38]},
      {stage4_17[17]}
   );
   gpc1_1 gpc10214 (
      {stage3_17[39]},
      {stage4_17[18]}
   );
   gpc1_1 gpc10215 (
      {stage3_17[40]},
      {stage4_17[19]}
   );
   gpc1_1 gpc10216 (
      {stage3_17[41]},
      {stage4_17[20]}
   );
   gpc1_1 gpc10217 (
      {stage3_17[42]},
      {stage4_17[21]}
   );
   gpc1_1 gpc10218 (
      {stage3_17[43]},
      {stage4_17[22]}
   );
   gpc1_1 gpc10219 (
      {stage3_18[52]},
      {stage4_18[20]}
   );
   gpc1_1 gpc10220 (
      {stage3_18[53]},
      {stage4_18[21]}
   );
   gpc1_1 gpc10221 (
      {stage3_18[54]},
      {stage4_18[22]}
   );
   gpc1_1 gpc10222 (
      {stage3_18[55]},
      {stage4_18[23]}
   );
   gpc1_1 gpc10223 (
      {stage3_18[56]},
      {stage4_18[24]}
   );
   gpc1_1 gpc10224 (
      {stage3_18[57]},
      {stage4_18[25]}
   );
   gpc1_1 gpc10225 (
      {stage3_18[58]},
      {stage4_18[26]}
   );
   gpc1_1 gpc10226 (
      {stage3_18[59]},
      {stage4_18[27]}
   );
   gpc1_1 gpc10227 (
      {stage3_18[60]},
      {stage4_18[28]}
   );
   gpc1_1 gpc10228 (
      {stage3_18[61]},
      {stage4_18[29]}
   );
   gpc1_1 gpc10229 (
      {stage3_18[62]},
      {stage4_18[30]}
   );
   gpc1_1 gpc10230 (
      {stage3_18[63]},
      {stage4_18[31]}
   );
   gpc1_1 gpc10231 (
      {stage3_20[57]},
      {stage4_20[21]}
   );
   gpc1_1 gpc10232 (
      {stage3_21[61]},
      {stage4_21[25]}
   );
   gpc1_1 gpc10233 (
      {stage3_21[62]},
      {stage4_21[26]}
   );
   gpc1_1 gpc10234 (
      {stage3_24[29]},
      {stage4_24[18]}
   );
   gpc1_1 gpc10235 (
      {stage3_24[30]},
      {stage4_24[19]}
   );
   gpc1_1 gpc10236 (
      {stage3_24[31]},
      {stage4_24[20]}
   );
   gpc1_1 gpc10237 (
      {stage3_24[32]},
      {stage4_24[21]}
   );
   gpc1_1 gpc10238 (
      {stage3_24[33]},
      {stage4_24[22]}
   );
   gpc1_1 gpc10239 (
      {stage3_24[34]},
      {stage4_24[23]}
   );
   gpc1_1 gpc10240 (
      {stage3_25[48]},
      {stage4_25[16]}
   );
   gpc1_1 gpc10241 (
      {stage3_25[49]},
      {stage4_25[17]}
   );
   gpc1_1 gpc10242 (
      {stage3_25[50]},
      {stage4_25[18]}
   );
   gpc1_1 gpc10243 (
      {stage3_25[51]},
      {stage4_25[19]}
   );
   gpc1_1 gpc10244 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc10245 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc10246 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc10247 (
      {stage3_28[57]},
      {stage4_28[19]}
   );
   gpc1_1 gpc10248 (
      {stage3_28[58]},
      {stage4_28[20]}
   );
   gpc1_1 gpc10249 (
      {stage3_28[59]},
      {stage4_28[21]}
   );
   gpc1_1 gpc10250 (
      {stage3_28[60]},
      {stage4_28[22]}
   );
   gpc1_1 gpc10251 (
      {stage3_28[61]},
      {stage4_28[23]}
   );
   gpc1_1 gpc10252 (
      {stage3_28[62]},
      {stage4_28[24]}
   );
   gpc1_1 gpc10253 (
      {stage3_28[63]},
      {stage4_28[25]}
   );
   gpc1_1 gpc10254 (
      {stage3_28[64]},
      {stage4_28[26]}
   );
   gpc1_1 gpc10255 (
      {stage3_28[65]},
      {stage4_28[27]}
   );
   gpc1_1 gpc10256 (
      {stage3_28[66]},
      {stage4_28[28]}
   );
   gpc1_1 gpc10257 (
      {stage3_28[67]},
      {stage4_28[29]}
   );
   gpc1_1 gpc10258 (
      {stage3_28[68]},
      {stage4_28[30]}
   );
   gpc1_1 gpc10259 (
      {stage3_28[69]},
      {stage4_28[31]}
   );
   gpc1_1 gpc10260 (
      {stage3_30[36]},
      {stage4_30[23]}
   );
   gpc1_1 gpc10261 (
      {stage3_30[37]},
      {stage4_30[24]}
   );
   gpc1_1 gpc10262 (
      {stage3_30[38]},
      {stage4_30[25]}
   );
   gpc1_1 gpc10263 (
      {stage3_32[51]},
      {stage4_32[19]}
   );
   gpc1_1 gpc10264 (
      {stage3_32[52]},
      {stage4_32[20]}
   );
   gpc1_1 gpc10265 (
      {stage3_32[53]},
      {stage4_32[21]}
   );
   gpc1_1 gpc10266 (
      {stage3_32[54]},
      {stage4_32[22]}
   );
   gpc1_1 gpc10267 (
      {stage3_32[55]},
      {stage4_32[23]}
   );
   gpc1_1 gpc10268 (
      {stage3_33[53]},
      {stage4_33[24]}
   );
   gpc1_1 gpc10269 (
      {stage3_33[54]},
      {stage4_33[25]}
   );
   gpc1_1 gpc10270 (
      {stage3_33[55]},
      {stage4_33[26]}
   );
   gpc1_1 gpc10271 (
      {stage3_33[56]},
      {stage4_33[27]}
   );
   gpc1_1 gpc10272 (
      {stage3_33[57]},
      {stage4_33[28]}
   );
   gpc1_1 gpc10273 (
      {stage3_33[58]},
      {stage4_33[29]}
   );
   gpc1_1 gpc10274 (
      {stage3_33[59]},
      {stage4_33[30]}
   );
   gpc1_1 gpc10275 (
      {stage3_33[60]},
      {stage4_33[31]}
   );
   gpc1_1 gpc10276 (
      {stage3_33[61]},
      {stage4_33[32]}
   );
   gpc1_1 gpc10277 (
      {stage3_33[62]},
      {stage4_33[33]}
   );
   gpc1_1 gpc10278 (
      {stage3_34[32]},
      {stage4_34[17]}
   );
   gpc1_1 gpc10279 (
      {stage3_34[33]},
      {stage4_34[18]}
   );
   gpc1_1 gpc10280 (
      {stage3_34[34]},
      {stage4_34[19]}
   );
   gpc1_1 gpc10281 (
      {stage3_34[35]},
      {stage4_34[20]}
   );
   gpc1_1 gpc10282 (
      {stage3_34[36]},
      {stage4_34[21]}
   );
   gpc1_1 gpc10283 (
      {stage3_34[37]},
      {stage4_34[22]}
   );
   gpc1_1 gpc10284 (
      {stage3_34[38]},
      {stage4_34[23]}
   );
   gpc1_1 gpc10285 (
      {stage3_34[39]},
      {stage4_34[24]}
   );
   gpc1_1 gpc10286 (
      {stage3_34[40]},
      {stage4_34[25]}
   );
   gpc1_1 gpc10287 (
      {stage3_34[41]},
      {stage4_34[26]}
   );
   gpc1_1 gpc10288 (
      {stage3_34[42]},
      {stage4_34[27]}
   );
   gpc1_1 gpc10289 (
      {stage3_34[43]},
      {stage4_34[28]}
   );
   gpc1_1 gpc10290 (
      {stage3_34[44]},
      {stage4_34[29]}
   );
   gpc1_1 gpc10291 (
      {stage3_35[52]},
      {stage4_35[19]}
   );
   gpc1_1 gpc10292 (
      {stage3_35[53]},
      {stage4_35[20]}
   );
   gpc1_1 gpc10293 (
      {stage3_35[54]},
      {stage4_35[21]}
   );
   gpc1_1 gpc10294 (
      {stage3_35[55]},
      {stage4_35[22]}
   );
   gpc1_1 gpc10295 (
      {stage3_35[56]},
      {stage4_35[23]}
   );
   gpc1_1 gpc10296 (
      {stage3_36[39]},
      {stage4_36[21]}
   );
   gpc1_1 gpc10297 (
      {stage3_36[40]},
      {stage4_36[22]}
   );
   gpc1_1 gpc10298 (
      {stage3_36[41]},
      {stage4_36[23]}
   );
   gpc1_1 gpc10299 (
      {stage3_36[42]},
      {stage4_36[24]}
   );
   gpc1_1 gpc10300 (
      {stage3_36[43]},
      {stage4_36[25]}
   );
   gpc1_1 gpc10301 (
      {stage3_36[44]},
      {stage4_36[26]}
   );
   gpc1_1 gpc10302 (
      {stage3_36[45]},
      {stage4_36[27]}
   );
   gpc1_1 gpc10303 (
      {stage3_36[46]},
      {stage4_36[28]}
   );
   gpc1_1 gpc10304 (
      {stage3_36[47]},
      {stage4_36[29]}
   );
   gpc1_1 gpc10305 (
      {stage3_36[48]},
      {stage4_36[30]}
   );
   gpc1_1 gpc10306 (
      {stage3_36[49]},
      {stage4_36[31]}
   );
   gpc1_1 gpc10307 (
      {stage3_36[50]},
      {stage4_36[32]}
   );
   gpc1_1 gpc10308 (
      {stage3_36[51]},
      {stage4_36[33]}
   );
   gpc1_1 gpc10309 (
      {stage3_36[52]},
      {stage4_36[34]}
   );
   gpc1_1 gpc10310 (
      {stage3_36[53]},
      {stage4_36[35]}
   );
   gpc1_1 gpc10311 (
      {stage3_36[54]},
      {stage4_36[36]}
   );
   gpc1_1 gpc10312 (
      {stage3_36[55]},
      {stage4_36[37]}
   );
   gpc1_1 gpc10313 (
      {stage3_38[60]},
      {stage4_38[18]}
   );
   gpc1_1 gpc10314 (
      {stage3_38[61]},
      {stage4_38[19]}
   );
   gpc1_1 gpc10315 (
      {stage3_38[62]},
      {stage4_38[20]}
   );
   gpc1_1 gpc10316 (
      {stage3_38[63]},
      {stage4_38[21]}
   );
   gpc1_1 gpc10317 (
      {stage3_38[64]},
      {stage4_38[22]}
   );
   gpc1_1 gpc10318 (
      {stage3_38[65]},
      {stage4_38[23]}
   );
   gpc1_1 gpc10319 (
      {stage3_38[66]},
      {stage4_38[24]}
   );
   gpc1_1 gpc10320 (
      {stage3_38[67]},
      {stage4_38[25]}
   );
   gpc1_1 gpc10321 (
      {stage3_38[68]},
      {stage4_38[26]}
   );
   gpc1_1 gpc10322 (
      {stage3_40[36]},
      {stage4_40[19]}
   );
   gpc1_1 gpc10323 (
      {stage3_40[37]},
      {stage4_40[20]}
   );
   gpc1_1 gpc10324 (
      {stage3_40[38]},
      {stage4_40[21]}
   );
   gpc1_1 gpc10325 (
      {stage3_40[39]},
      {stage4_40[22]}
   );
   gpc1_1 gpc10326 (
      {stage3_40[40]},
      {stage4_40[23]}
   );
   gpc1_1 gpc10327 (
      {stage3_40[41]},
      {stage4_40[24]}
   );
   gpc1_1 gpc10328 (
      {stage3_40[42]},
      {stage4_40[25]}
   );
   gpc1_1 gpc10329 (
      {stage3_40[43]},
      {stage4_40[26]}
   );
   gpc1_1 gpc10330 (
      {stage3_40[44]},
      {stage4_40[27]}
   );
   gpc1_1 gpc10331 (
      {stage3_40[45]},
      {stage4_40[28]}
   );
   gpc1_1 gpc10332 (
      {stage3_41[54]},
      {stage4_41[21]}
   );
   gpc1_1 gpc10333 (
      {stage3_41[55]},
      {stage4_41[22]}
   );
   gpc1_1 gpc10334 (
      {stage3_41[56]},
      {stage4_41[23]}
   );
   gpc1_1 gpc10335 (
      {stage3_43[55]},
      {stage4_43[18]}
   );
   gpc1_1 gpc10336 (
      {stage3_43[56]},
      {stage4_43[19]}
   );
   gpc1_1 gpc10337 (
      {stage3_43[57]},
      {stage4_43[20]}
   );
   gpc1_1 gpc10338 (
      {stage3_43[58]},
      {stage4_43[21]}
   );
   gpc1_1 gpc10339 (
      {stage3_43[59]},
      {stage4_43[22]}
   );
   gpc1_1 gpc10340 (
      {stage3_44[68]},
      {stage4_44[23]}
   );
   gpc1_1 gpc10341 (
      {stage3_44[69]},
      {stage4_44[24]}
   );
   gpc1_1 gpc10342 (
      {stage3_44[70]},
      {stage4_44[25]}
   );
   gpc1_1 gpc10343 (
      {stage3_44[71]},
      {stage4_44[26]}
   );
   gpc1_1 gpc10344 (
      {stage3_44[72]},
      {stage4_44[27]}
   );
   gpc1_1 gpc10345 (
      {stage3_44[73]},
      {stage4_44[28]}
   );
   gpc1_1 gpc10346 (
      {stage3_44[74]},
      {stage4_44[29]}
   );
   gpc1_1 gpc10347 (
      {stage3_44[75]},
      {stage4_44[30]}
   );
   gpc1_1 gpc10348 (
      {stage3_44[76]},
      {stage4_44[31]}
   );
   gpc1_1 gpc10349 (
      {stage3_44[77]},
      {stage4_44[32]}
   );
   gpc1_1 gpc10350 (
      {stage3_44[78]},
      {stage4_44[33]}
   );
   gpc1_1 gpc10351 (
      {stage3_44[79]},
      {stage4_44[34]}
   );
   gpc1_1 gpc10352 (
      {stage3_44[80]},
      {stage4_44[35]}
   );
   gpc1_1 gpc10353 (
      {stage3_44[81]},
      {stage4_44[36]}
   );
   gpc1_1 gpc10354 (
      {stage3_44[82]},
      {stage4_44[37]}
   );
   gpc1_1 gpc10355 (
      {stage3_44[83]},
      {stage4_44[38]}
   );
   gpc1_1 gpc10356 (
      {stage3_44[84]},
      {stage4_44[39]}
   );
   gpc1_1 gpc10357 (
      {stage3_46[46]},
      {stage4_46[22]}
   );
   gpc1_1 gpc10358 (
      {stage3_46[47]},
      {stage4_46[23]}
   );
   gpc1_1 gpc10359 (
      {stage3_46[48]},
      {stage4_46[24]}
   );
   gpc1_1 gpc10360 (
      {stage3_47[71]},
      {stage4_47[23]}
   );
   gpc1_1 gpc10361 (
      {stage3_47[72]},
      {stage4_47[24]}
   );
   gpc1_1 gpc10362 (
      {stage3_47[73]},
      {stage4_47[25]}
   );
   gpc1_1 gpc10363 (
      {stage3_49[54]},
      {stage4_49[17]}
   );
   gpc1_1 gpc10364 (
      {stage3_49[55]},
      {stage4_49[18]}
   );
   gpc1_1 gpc10365 (
      {stage3_49[56]},
      {stage4_49[19]}
   );
   gpc1_1 gpc10366 (
      {stage3_49[57]},
      {stage4_49[20]}
   );
   gpc1_1 gpc10367 (
      {stage3_49[58]},
      {stage4_49[21]}
   );
   gpc1_1 gpc10368 (
      {stage3_49[59]},
      {stage4_49[22]}
   );
   gpc1_1 gpc10369 (
      {stage3_49[60]},
      {stage4_49[23]}
   );
   gpc1_1 gpc10370 (
      {stage3_49[61]},
      {stage4_49[24]}
   );
   gpc1_1 gpc10371 (
      {stage3_49[62]},
      {stage4_49[25]}
   );
   gpc1_1 gpc10372 (
      {stage3_49[63]},
      {stage4_49[26]}
   );
   gpc1_1 gpc10373 (
      {stage3_49[64]},
      {stage4_49[27]}
   );
   gpc1_1 gpc10374 (
      {stage3_50[63]},
      {stage4_50[23]}
   );
   gpc1_1 gpc10375 (
      {stage3_52[54]},
      {stage4_52[21]}
   );
   gpc1_1 gpc10376 (
      {stage3_52[55]},
      {stage4_52[22]}
   );
   gpc1_1 gpc10377 (
      {stage3_54[54]},
      {stage4_54[22]}
   );
   gpc1_1 gpc10378 (
      {stage3_54[55]},
      {stage4_54[23]}
   );
   gpc1_1 gpc10379 (
      {stage3_54[56]},
      {stage4_54[24]}
   );
   gpc1_1 gpc10380 (
      {stage3_54[57]},
      {stage4_54[25]}
   );
   gpc1_1 gpc10381 (
      {stage3_54[58]},
      {stage4_54[26]}
   );
   gpc1_1 gpc10382 (
      {stage3_54[59]},
      {stage4_54[27]}
   );
   gpc1_1 gpc10383 (
      {stage3_54[60]},
      {stage4_54[28]}
   );
   gpc1_1 gpc10384 (
      {stage3_54[61]},
      {stage4_54[29]}
   );
   gpc1_1 gpc10385 (
      {stage3_54[62]},
      {stage4_54[30]}
   );
   gpc1_1 gpc10386 (
      {stage3_55[40]},
      {stage4_55[22]}
   );
   gpc1_1 gpc10387 (
      {stage3_55[41]},
      {stage4_55[23]}
   );
   gpc1_1 gpc10388 (
      {stage3_55[42]},
      {stage4_55[24]}
   );
   gpc1_1 gpc10389 (
      {stage3_55[43]},
      {stage4_55[25]}
   );
   gpc1_1 gpc10390 (
      {stage3_55[44]},
      {stage4_55[26]}
   );
   gpc1_1 gpc10391 (
      {stage3_55[45]},
      {stage4_55[27]}
   );
   gpc1_1 gpc10392 (
      {stage3_55[46]},
      {stage4_55[28]}
   );
   gpc1_1 gpc10393 (
      {stage3_56[26]},
      {stage4_56[16]}
   );
   gpc1_1 gpc10394 (
      {stage3_56[27]},
      {stage4_56[17]}
   );
   gpc1_1 gpc10395 (
      {stage3_56[28]},
      {stage4_56[18]}
   );
   gpc1_1 gpc10396 (
      {stage3_56[29]},
      {stage4_56[19]}
   );
   gpc1_1 gpc10397 (
      {stage3_56[30]},
      {stage4_56[20]}
   );
   gpc1_1 gpc10398 (
      {stage3_56[31]},
      {stage4_56[21]}
   );
   gpc1_1 gpc10399 (
      {stage3_56[32]},
      {stage4_56[22]}
   );
   gpc1_1 gpc10400 (
      {stage3_56[33]},
      {stage4_56[23]}
   );
   gpc1_1 gpc10401 (
      {stage3_56[34]},
      {stage4_56[24]}
   );
   gpc1_1 gpc10402 (
      {stage3_56[35]},
      {stage4_56[25]}
   );
   gpc1_1 gpc10403 (
      {stage3_56[36]},
      {stage4_56[26]}
   );
   gpc1_1 gpc10404 (
      {stage3_56[37]},
      {stage4_56[27]}
   );
   gpc1_1 gpc10405 (
      {stage3_56[38]},
      {stage4_56[28]}
   );
   gpc1_1 gpc10406 (
      {stage3_57[51]},
      {stage4_57[23]}
   );
   gpc1_1 gpc10407 (
      {stage3_57[52]},
      {stage4_57[24]}
   );
   gpc1_1 gpc10408 (
      {stage3_58[48]},
      {stage4_58[15]}
   );
   gpc1_1 gpc10409 (
      {stage3_59[45]},
      {stage4_59[15]}
   );
   gpc1_1 gpc10410 (
      {stage3_60[49]},
      {stage4_60[21]}
   );
   gpc1_1 gpc10411 (
      {stage3_60[50]},
      {stage4_60[22]}
   );
   gpc1_1 gpc10412 (
      {stage3_60[51]},
      {stage4_60[23]}
   );
   gpc1_1 gpc10413 (
      {stage3_60[52]},
      {stage4_60[24]}
   );
   gpc1_1 gpc10414 (
      {stage3_61[55]},
      {stage4_61[27]}
   );
   gpc1_1 gpc10415 (
      {stage3_61[56]},
      {stage4_61[28]}
   );
   gpc1_1 gpc10416 (
      {stage3_62[34]},
      {stage4_62[17]}
   );
   gpc1_1 gpc10417 (
      {stage3_62[35]},
      {stage4_62[18]}
   );
   gpc1_1 gpc10418 (
      {stage3_62[36]},
      {stage4_62[19]}
   );
   gpc1_1 gpc10419 (
      {stage3_62[37]},
      {stage4_62[20]}
   );
   gpc1_1 gpc10420 (
      {stage3_62[38]},
      {stage4_62[21]}
   );
   gpc1_1 gpc10421 (
      {stage3_62[39]},
      {stage4_62[22]}
   );
   gpc1_1 gpc10422 (
      {stage3_62[40]},
      {stage4_62[23]}
   );
   gpc1_1 gpc10423 (
      {stage3_67[13]},
      {stage4_67[15]}
   );
   gpc1_1 gpc10424 (
      {stage3_67[14]},
      {stage4_67[16]}
   );
   gpc606_5 gpc10425 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1406_5 gpc10426 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc1163_5 gpc10427 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[4]},
      {stage4_5[1]},
      {stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc606_5 gpc10428 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16], stage4_3[17]},
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage5_7[0],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc606_5 gpc10429 (
      {stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[1],stage5_6[3],stage5_5[4],stage5_4[4]}
   );
   gpc606_5 gpc10430 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[2],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc10431 (
      {stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21], stage4_4[22]},
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17]},
      {stage5_8[2],stage5_7[3],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc606_5 gpc10432 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc10433 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc10434 (
      {stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24], stage4_5[25]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[5],stage5_7[6],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc10435 (
      {stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage4_7[18], stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23]},
      {stage5_9[3],stage5_8[6],stage5_7[7],stage5_6[9],stage5_5[10]}
   );
   gpc606_5 gpc10436 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37]},
      {stage4_7[24], stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29]},
      {stage5_9[4],stage5_8[7],stage5_7[8],stage5_6[10],stage5_5[11]}
   );
   gpc615_5 gpc10437 (
      {stage4_7[30], stage4_7[31], stage4_7[32], stage4_7[33], stage4_7[34]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[5],stage5_8[8],stage5_7[9]}
   );
   gpc615_5 gpc10438 (
      {stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38], stage4_7[39]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[6],stage5_8[9],stage5_7[10]}
   );
   gpc1406_5 gpc10439 (
      {stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[7],stage5_8[10]}
   );
   gpc215_4 gpc10440 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage5_11[3],stage5_10[3],stage5_9[8],stage5_8[11]}
   );
   gpc215_4 gpc10441 (
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[13]},
      {stage4_10[6], stage4_10[7]},
      {stage5_11[4],stage5_10[4],stage5_9[9],stage5_8[12]}
   );
   gpc207_4 gpc10442 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24]},
      {stage4_10[8], stage4_10[9]},
      {stage5_11[5],stage5_10[5],stage5_9[10],stage5_8[13]}
   );
   gpc606_5 gpc10443 (
      {stage4_8[25], stage4_8[26], stage4_8[27], stage4_8[28], stage4_8[29], stage4_8[30]},
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15]},
      {stage5_12[1],stage5_11[6],stage5_10[6],stage5_9[11],stage5_8[14]}
   );
   gpc606_5 gpc10444 (
      {stage4_8[31], stage4_8[32], stage4_8[33], stage4_8[34], 1'b0, 1'b0},
      {stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19], stage4_10[20], stage4_10[21]},
      {stage5_12[2],stage5_11[7],stage5_10[7],stage5_9[12],stage5_8[15]}
   );
   gpc1163_5 gpc10445 (
      {stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[0]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[3],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc10446 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], 1'b0},
      {stage4_11[7]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[1],stage5_12[4],stage5_11[9],stage5_10[9]}
   );
   gpc615_5 gpc10447 (
      {stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12]},
      {stage4_12[7]},
      {stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[5],stage5_11[10]}
   );
   gpc615_5 gpc10448 (
      {stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage4_12[8]},
      {stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[6],stage5_11[11]}
   );
   gpc615_5 gpc10449 (
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22]},
      {stage4_12[9]},
      {stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[7],stage5_11[12]}
   );
   gpc615_5 gpc10450 (
      {stage4_11[23], stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27]},
      {stage4_12[10]},
      {stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[8],stage5_11[13]}
   );
   gpc615_5 gpc10451 (
      {stage4_12[11], stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15]},
      {stage4_13[25]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[9]}
   );
   gpc615_5 gpc10452 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc10453 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc10454 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc10455 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[10]}
   );
   gpc615_5 gpc10456 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc10457 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc10458 (
      {stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc606_5 gpc10459 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7],stage5_17[7]}
   );
   gpc2116_5 gpc10460 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[6]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc2116_5 gpc10461 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[1]},
      {stage4_21[2], stage4_21[3]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc2116_5 gpc10462 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[8]},
      {stage4_20[2]},
      {stage4_21[4], stage4_21[5]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc10463 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[9]},
      {stage4_20[3], stage4_20[4], stage4_20[5], stage4_20[6], stage4_20[7], stage4_20[8]},
      {stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[7],stage5_18[11]}
   );
   gpc615_5 gpc10464 (
      {stage4_18[23], stage4_18[24], stage4_18[25], stage4_18[26], stage4_18[27]},
      {stage4_19[10]},
      {stage4_20[9], stage4_20[10], stage4_20[11], stage4_20[12], stage4_20[13], stage4_20[14]},
      {stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[8],stage5_18[12]}
   );
   gpc615_5 gpc10465 (
      {stage4_18[28], stage4_18[29], stage4_18[30], stage4_18[31], 1'b0},
      {stage4_19[11]},
      {stage4_20[15], stage4_20[16], stage4_20[17], stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[9],stage5_18[13]}
   );
   gpc615_5 gpc10466 (
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16]},
      {stage4_20[21]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[0],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc7_3 gpc10467 (
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[1],stage5_22[7],stage5_21[8]}
   );
   gpc7_3 gpc10468 (
      {stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23], stage4_21[24], stage4_21[25]},
      {stage5_23[2],stage5_22[8],stage5_21[9]}
   );
   gpc1163_5 gpc10469 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[3],stage5_22[9]}
   );
   gpc1163_5 gpc10470 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage4_24[1]},
      {stage4_25[1]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[4],stage5_22[10]}
   );
   gpc1163_5 gpc10471 (
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[2]},
      {stage4_25[2]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[5],stage5_22[11]}
   );
   gpc615_5 gpc10472 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[18]},
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[6],stage5_22[12]}
   );
   gpc615_5 gpc10473 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[19]},
      {stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12], stage4_24[13], stage4_24[14]},
      {stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[7],stage5_22[13]}
   );
   gpc615_5 gpc10474 (
      {stage4_22[19], stage4_22[20], 1'b0, 1'b0, 1'b0},
      {stage4_23[20]},
      {stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18], stage4_24[19], stage4_24[20]},
      {stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[8],stage5_22[14]}
   );
   gpc606_5 gpc10475 (
      {stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[6],stage5_25[6]}
   );
   gpc606_5 gpc10476 (
      {stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12], stage4_25[13], stage4_25[14]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[7],stage5_25[7]}
   );
   gpc207_4 gpc10477 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[8]}
   );
   gpc207_4 gpc10478 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {stage4_28[2], stage4_28[3]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[9]}
   );
   gpc615_5 gpc10479 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_28[4]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4]}
   );
   gpc606_5 gpc10480 (
      {stage4_28[5], stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[5],stage5_28[5]}
   );
   gpc606_5 gpc10481 (
      {stage4_28[11], stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[6],stage5_28[6]}
   );
   gpc606_5 gpc10482 (
      {stage4_28[17], stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[3],stage5_30[3],stage5_29[7],stage5_28[7]}
   );
   gpc606_5 gpc10483 (
      {stage4_28[23], stage4_28[24], stage4_28[25], stage4_28[26], stage4_28[27], stage4_28[28]},
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23]},
      {stage5_32[3],stage5_31[4],stage5_30[4],stage5_29[8],stage5_28[8]}
   );
   gpc207_4 gpc10484 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[4],stage5_31[5],stage5_30[5],stage5_29[9]}
   );
   gpc207_4 gpc10485 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17], stage4_29[18], stage4_29[19]},
      {stage4_31[2], stage4_31[3]},
      {stage5_32[5],stage5_31[6],stage5_30[6],stage5_29[10]}
   );
   gpc615_5 gpc10486 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[0]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[6],stage5_31[7]}
   );
   gpc615_5 gpc10487 (
      {stage4_31[9], stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13]},
      {stage4_32[1]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[1],stage5_33[1],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc10488 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[2],stage5_34[2],stage5_33[2],stage5_32[8]}
   );
   gpc606_5 gpc10489 (
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage5_36[1],stage5_35[3],stage5_34[3],stage5_33[3],stage5_32[9]}
   );
   gpc606_5 gpc10490 (
      {stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17], stage4_32[18], stage4_32[19]},
      {stage4_34[12], stage4_34[13], stage4_34[14], stage4_34[15], stage4_34[16], stage4_34[17]},
      {stage5_36[2],stage5_35[4],stage5_34[4],stage5_33[4],stage5_32[10]}
   );
   gpc606_5 gpc10491 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[3],stage5_35[5],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc10492 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[4],stage5_35[6],stage5_34[6],stage5_33[6]}
   );
   gpc606_5 gpc10493 (
      {stage4_33[24], stage4_33[25], stage4_33[26], stage4_33[27], stage4_33[28], stage4_33[29]},
      {stage4_35[12], stage4_35[13], stage4_35[14], stage4_35[15], stage4_35[16], stage4_35[17]},
      {stage5_37[2],stage5_36[5],stage5_35[7],stage5_34[7],stage5_33[7]}
   );
   gpc606_5 gpc10494 (
      {stage4_33[30], stage4_33[31], stage4_33[32], stage4_33[33], 1'b0, 1'b0},
      {stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21], stage4_35[22], stage4_35[23]},
      {stage5_37[3],stage5_36[6],stage5_35[8],stage5_34[8],stage5_33[8]}
   );
   gpc1163_5 gpc10495 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[4],stage5_36[7]}
   );
   gpc1163_5 gpc10496 (
      {stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage4_38[1]},
      {stage4_39[1]},
      {stage5_40[1],stage5_39[1],stage5_38[1],stage5_37[5],stage5_36[8]}
   );
   gpc1163_5 gpc10497 (
      {stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], 1'b0, 1'b0},
      {stage4_38[2]},
      {stage4_39[2]},
      {stage5_40[2],stage5_39[2],stage5_38[2],stage5_37[6],stage5_36[9]}
   );
   gpc606_5 gpc10498 (
      {stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12], stage4_36[13], stage4_36[14]},
      {stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6], stage4_38[7], stage4_38[8]},
      {stage5_40[3],stage5_39[3],stage5_38[3],stage5_37[7],stage5_36[10]}
   );
   gpc606_5 gpc10499 (
      {stage4_36[15], stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20]},
      {stage4_38[9], stage4_38[10], stage4_38[11], stage4_38[12], stage4_38[13], stage4_38[14]},
      {stage5_40[4],stage5_39[4],stage5_38[4],stage5_37[8],stage5_36[11]}
   );
   gpc606_5 gpc10500 (
      {stage4_36[21], stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26]},
      {stage4_38[15], stage4_38[16], stage4_38[17], stage4_38[18], stage4_38[19], stage4_38[20]},
      {stage5_40[5],stage5_39[5],stage5_38[5],stage5_37[9],stage5_36[12]}
   );
   gpc606_5 gpc10501 (
      {stage4_36[27], stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32]},
      {stage4_38[21], stage4_38[22], stage4_38[23], stage4_38[24], stage4_38[25], stage4_38[26]},
      {stage5_40[6],stage5_39[6],stage5_38[6],stage5_37[10],stage5_36[13]}
   );
   gpc135_4 gpc10502 (
      {stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6], stage4_39[7]},
      {stage4_40[0], stage4_40[1], stage4_40[2]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[7],stage5_39[7]}
   );
   gpc135_4 gpc10503 (
      {stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12]},
      {stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[8],stage5_39[8]}
   );
   gpc135_4 gpc10504 (
      {stage4_39[13], stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17]},
      {stage4_40[6], stage4_40[7], stage4_40[8]},
      {stage4_41[2]},
      {stage5_42[2],stage5_41[2],stage5_40[9],stage5_39[9]}
   );
   gpc615_5 gpc10505 (
      {stage4_39[18], stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22]},
      {stage4_40[9]},
      {stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7], stage4_41[8]},
      {stage5_43[0],stage5_42[3],stage5_41[3],stage5_40[10],stage5_39[10]}
   );
   gpc606_5 gpc10506 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[4],stage5_41[4],stage5_40[11]}
   );
   gpc606_5 gpc10507 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[2],stage5_42[5],stage5_41[5],stage5_40[12]}
   );
   gpc606_5 gpc10508 (
      {stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13], stage4_41[14]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[3],stage5_42[6],stage5_41[6]}
   );
   gpc606_5 gpc10509 (
      {stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19], stage4_41[20]},
      {stage4_43[6], stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage5_45[1],stage5_44[3],stage5_43[4],stage5_42[7],stage5_41[7]}
   );
   gpc606_5 gpc10510 (
      {stage4_41[21], stage4_41[22], stage4_41[23], 1'b0, 1'b0, 1'b0},
      {stage4_43[12], stage4_43[13], stage4_43[14], stage4_43[15], stage4_43[16], stage4_43[17]},
      {stage5_45[2],stage5_44[4],stage5_43[5],stage5_42[8],stage5_41[8]}
   );
   gpc7_3 gpc10511 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17], stage4_42[18]},
      {stage5_44[5],stage5_43[6],stage5_42[9]}
   );
   gpc615_5 gpc10512 (
      {stage4_43[18], stage4_43[19], stage4_43[20], stage4_43[21], stage4_43[22]},
      {stage4_44[0]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[3],stage5_44[6],stage5_43[7]}
   );
   gpc135_4 gpc10513 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[1],stage5_45[4],stage5_44[7]}
   );
   gpc135_4 gpc10514 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[2],stage5_45[5],stage5_44[8]}
   );
   gpc135_4 gpc10515 (
      {stage4_44[11], stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[3],stage5_45[6],stage5_44[9]}
   );
   gpc135_4 gpc10516 (
      {stage4_44[16], stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20]},
      {stage4_45[15], stage4_45[16], stage4_45[17]},
      {stage4_46[3]},
      {stage5_47[4],stage5_46[4],stage5_45[7],stage5_44[10]}
   );
   gpc135_4 gpc10517 (
      {stage4_44[21], stage4_44[22], stage4_44[23], stage4_44[24], stage4_44[25]},
      {stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_46[4]},
      {stage5_47[5],stage5_46[5],stage5_45[8],stage5_44[11]}
   );
   gpc606_5 gpc10518 (
      {stage4_45[21], stage4_45[22], stage4_45[23], stage4_45[24], stage4_45[25], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[6],stage5_46[6],stage5_45[9]}
   );
   gpc2135_5 gpc10519 (
      {stage4_46[5], stage4_46[6], stage4_46[7], stage4_46[8], stage4_46[9]},
      {stage4_47[6], stage4_47[7], stage4_47[8]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[7],stage5_46[7]}
   );
   gpc2135_5 gpc10520 (
      {stage4_46[10], stage4_46[11], stage4_46[12], stage4_46[13], stage4_46[14]},
      {stage4_47[9], stage4_47[10], stage4_47[11]},
      {stage4_48[1]},
      {stage4_49[2], stage4_49[3]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[8],stage5_46[8]}
   );
   gpc2135_5 gpc10521 (
      {stage4_46[15], stage4_46[16], stage4_46[17], stage4_46[18], stage4_46[19]},
      {stage4_47[12], stage4_47[13], stage4_47[14]},
      {stage4_48[2]},
      {stage4_49[4], stage4_49[5]},
      {stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[9],stage5_46[9]}
   );
   gpc615_5 gpc10522 (
      {stage4_46[20], stage4_46[21], stage4_46[22], stage4_46[23], stage4_46[24]},
      {stage4_47[15]},
      {stage4_48[3], stage4_48[4], stage4_48[5], stage4_48[6], stage4_48[7], stage4_48[8]},
      {stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[10],stage5_46[10]}
   );
   gpc615_5 gpc10523 (
      {stage4_47[16], stage4_47[17], stage4_47[18], stage4_47[19], stage4_47[20]},
      {stage4_48[9]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[0],stage5_50[4],stage5_49[5],stage5_48[5],stage5_47[11]}
   );
   gpc615_5 gpc10524 (
      {stage4_47[21], stage4_47[22], stage4_47[23], stage4_47[24], stage4_47[25]},
      {stage4_48[10]},
      {stage4_49[12], stage4_49[13], stage4_49[14], stage4_49[15], stage4_49[16], stage4_49[17]},
      {stage5_51[1],stage5_50[5],stage5_49[6],stage5_48[6],stage5_47[12]}
   );
   gpc7_3 gpc10525 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[6]}
   );
   gpc7_3 gpc10526 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11], stage4_50[12], stage4_50[13]},
      {stage5_52[1],stage5_51[3],stage5_50[7]}
   );
   gpc615_5 gpc10527 (
      {stage4_50[14], stage4_50[15], stage4_50[16], stage4_50[17], stage4_50[18]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[2],stage5_51[4],stage5_50[8]}
   );
   gpc615_5 gpc10528 (
      {stage4_50[19], stage4_50[20], stage4_50[21], stage4_50[22], stage4_50[23]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[3],stage5_51[5],stage5_50[9]}
   );
   gpc117_4 gpc10529 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6], stage4_51[7], stage4_51[8]},
      {stage4_52[12]},
      {stage4_53[0]},
      {stage5_54[2],stage5_53[2],stage5_52[4],stage5_51[6]}
   );
   gpc606_5 gpc10530 (
      {stage4_51[9], stage4_51[10], stage4_51[11], stage4_51[12], stage4_51[13], stage4_51[14]},
      {stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5], stage4_53[6]},
      {stage5_55[0],stage5_54[3],stage5_53[3],stage5_52[5],stage5_51[7]}
   );
   gpc606_5 gpc10531 (
      {stage4_51[15], stage4_51[16], stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20]},
      {stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11], stage4_53[12]},
      {stage5_55[1],stage5_54[4],stage5_53[4],stage5_52[6],stage5_51[8]}
   );
   gpc606_5 gpc10532 (
      {stage4_51[21], stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17], stage4_53[18]},
      {stage5_55[2],stage5_54[5],stage5_53[5],stage5_52[7],stage5_51[9]}
   );
   gpc606_5 gpc10533 (
      {stage4_52[13], stage4_52[14], stage4_52[15], stage4_52[16], stage4_52[17], stage4_52[18]},
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5]},
      {stage5_56[0],stage5_55[3],stage5_54[6],stage5_53[6],stage5_52[8]}
   );
   gpc606_5 gpc10534 (
      {stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23], stage4_53[24]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[1],stage5_55[4],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc10535 (
      {stage4_54[6], stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10]},
      {stage4_55[6]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[1],stage5_56[2],stage5_55[5],stage5_54[8]}
   );
   gpc615_5 gpc10536 (
      {stage4_54[11], stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15]},
      {stage4_55[7]},
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage5_58[1],stage5_57[2],stage5_56[3],stage5_55[6],stage5_54[9]}
   );
   gpc615_5 gpc10537 (
      {stage4_54[16], stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20]},
      {stage4_55[8]},
      {stage4_56[12], stage4_56[13], stage4_56[14], stage4_56[15], stage4_56[16], stage4_56[17]},
      {stage5_58[2],stage5_57[3],stage5_56[4],stage5_55[7],stage5_54[10]}
   );
   gpc615_5 gpc10538 (
      {stage4_54[21], stage4_54[22], stage4_54[23], stage4_54[24], stage4_54[25]},
      {stage4_55[9]},
      {stage4_56[18], stage4_56[19], stage4_56[20], stage4_56[21], stage4_56[22], stage4_56[23]},
      {stage5_58[3],stage5_57[4],stage5_56[5],stage5_55[8],stage5_54[11]}
   );
   gpc606_5 gpc10539 (
      {stage4_55[10], stage4_55[11], stage4_55[12], stage4_55[13], stage4_55[14], stage4_55[15]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage5_59[0],stage5_58[4],stage5_57[5],stage5_56[6],stage5_55[9]}
   );
   gpc606_5 gpc10540 (
      {stage4_55[16], stage4_55[17], stage4_55[18], stage4_55[19], stage4_55[20], stage4_55[21]},
      {stage4_57[6], stage4_57[7], stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11]},
      {stage5_59[1],stage5_58[5],stage5_57[6],stage5_56[7],stage5_55[10]}
   );
   gpc207_4 gpc10541 (
      {stage4_57[12], stage4_57[13], stage4_57[14], stage4_57[15], stage4_57[16], stage4_57[17], stage4_57[18]},
      {stage4_59[0], stage4_59[1]},
      {stage5_60[0],stage5_59[2],stage5_58[6],stage5_57[7]}
   );
   gpc207_4 gpc10542 (
      {stage4_57[19], stage4_57[20], stage4_57[21], stage4_57[22], stage4_57[23], stage4_57[24], 1'b0},
      {stage4_59[2], stage4_59[3]},
      {stage5_60[1],stage5_59[3],stage5_58[7],stage5_57[8]}
   );
   gpc606_5 gpc10543 (
      {stage4_59[4], stage4_59[5], stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[2],stage5_59[4]}
   );
   gpc606_5 gpc10544 (
      {stage4_59[10], stage4_59[11], stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[3],stage5_59[5]}
   );
   gpc606_5 gpc10545 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[2],stage5_61[2],stage5_60[4]}
   );
   gpc606_5 gpc10546 (
      {stage4_60[6], stage4_60[7], stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11]},
      {stage4_62[6], stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage5_64[1],stage5_63[3],stage5_62[3],stage5_61[3],stage5_60[5]}
   );
   gpc606_5 gpc10547 (
      {stage4_60[12], stage4_60[13], stage4_60[14], stage4_60[15], stage4_60[16], stage4_60[17]},
      {stage4_62[12], stage4_62[13], stage4_62[14], stage4_62[15], stage4_62[16], stage4_62[17]},
      {stage5_64[2],stage5_63[4],stage5_62[4],stage5_61[4],stage5_60[6]}
   );
   gpc7_3 gpc10548 (
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17], stage4_61[18]},
      {stage5_63[5],stage5_62[5],stage5_61[5]}
   );
   gpc7_3 gpc10549 (
      {stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22], stage4_61[23], stage4_61[24], stage4_61[25]},
      {stage5_63[6],stage5_62[6],stage5_61[6]}
   );
   gpc606_5 gpc10550 (
      {stage4_62[18], stage4_62[19], stage4_62[20], stage4_62[21], stage4_62[22], stage4_62[23]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[0],stage5_64[3],stage5_63[7],stage5_62[7]}
   );
   gpc606_5 gpc10551 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[4],stage5_63[8]}
   );
   gpc606_5 gpc10552 (
      {stage4_63[6], stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8], stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[5],stage5_63[9]}
   );
   gpc606_5 gpc10553 (
      {stage4_63[12], stage4_63[13], stage4_63[14], stage4_63[15], stage4_63[16], stage4_63[17]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage5_67[2],stage5_66[3],stage5_65[3],stage5_64[6],stage5_63[10]}
   );
   gpc135_4 gpc10554 (
      {stage4_64[6], stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10]},
      {stage4_65[18], stage4_65[19], stage4_65[20]},
      {stage4_66[0]},
      {stage5_67[3],stage5_66[4],stage5_65[4],stage5_64[7]}
   );
   gpc135_4 gpc10555 (
      {stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15]},
      {stage4_65[21], stage4_65[22], 1'b0},
      {stage4_66[1]},
      {stage5_67[4],stage5_66[5],stage5_65[5],stage5_64[8]}
   );
   gpc1163_5 gpc10556 (
      {stage4_66[2], stage4_66[3], stage4_66[4]},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage4_68[0]},
      {stage4_69[0]},
      {stage5_70[0],stage5_69[0],stage5_68[0],stage5_67[5],stage5_66[6]}
   );
   gpc1163_5 gpc10557 (
      {stage4_66[5], stage4_66[6], stage4_66[7]},
      {stage4_67[6], stage4_67[7], stage4_67[8], stage4_67[9], stage4_67[10], stage4_67[11]},
      {stage4_68[1]},
      {stage4_69[1]},
      {stage5_70[1],stage5_69[1],stage5_68[1],stage5_67[6],stage5_66[7]}
   );
   gpc1163_5 gpc10558 (
      {stage4_66[8], stage4_66[9], stage4_66[10]},
      {stage4_67[12], stage4_67[13], stage4_67[14], stage4_67[15], stage4_67[16], 1'b0},
      {stage4_68[2]},
      {stage4_69[2]},
      {stage5_70[2],stage5_69[2],stage5_68[2],stage5_67[7],stage5_66[8]}
   );
   gpc1_1 gpc10559 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc10560 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc10561 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc10562 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc10563 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc10564 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc10565 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc10566 (
      {stage4_3[18]},
      {stage5_3[4]}
   );
   gpc1_1 gpc10567 (
      {stage4_3[19]},
      {stage5_3[5]}
   );
   gpc1_1 gpc10568 (
      {stage4_3[20]},
      {stage5_3[6]}
   );
   gpc1_1 gpc10569 (
      {stage4_3[21]},
      {stage5_3[7]}
   );
   gpc1_1 gpc10570 (
      {stage4_4[23]},
      {stage5_4[7]}
   );
   gpc1_1 gpc10571 (
      {stage4_4[24]},
      {stage5_4[8]}
   );
   gpc1_1 gpc10572 (
      {stage4_5[38]},
      {stage5_5[12]}
   );
   gpc1_1 gpc10573 (
      {stage4_5[39]},
      {stage5_5[13]}
   );
   gpc1_1 gpc10574 (
      {stage4_5[40]},
      {stage5_5[14]}
   );
   gpc1_1 gpc10575 (
      {stage4_5[41]},
      {stage5_5[15]}
   );
   gpc1_1 gpc10576 (
      {stage4_5[42]},
      {stage5_5[16]}
   );
   gpc1_1 gpc10577 (
      {stage4_5[43]},
      {stage5_5[17]}
   );
   gpc1_1 gpc10578 (
      {stage4_5[44]},
      {stage5_5[18]}
   );
   gpc1_1 gpc10579 (
      {stage4_5[45]},
      {stage5_5[19]}
   );
   gpc1_1 gpc10580 (
      {stage4_5[46]},
      {stage5_5[20]}
   );
   gpc1_1 gpc10581 (
      {stage4_6[18]},
      {stage5_6[11]}
   );
   gpc1_1 gpc10582 (
      {stage4_6[19]},
      {stage5_6[12]}
   );
   gpc1_1 gpc10583 (
      {stage4_6[20]},
      {stage5_6[13]}
   );
   gpc1_1 gpc10584 (
      {stage4_11[28]},
      {stage5_11[14]}
   );
   gpc1_1 gpc10585 (
      {stage4_11[29]},
      {stage5_11[15]}
   );
   gpc1_1 gpc10586 (
      {stage4_11[30]},
      {stage5_11[16]}
   );
   gpc1_1 gpc10587 (
      {stage4_11[31]},
      {stage5_11[17]}
   );
   gpc1_1 gpc10588 (
      {stage4_11[32]},
      {stage5_11[18]}
   );
   gpc1_1 gpc10589 (
      {stage4_11[33]},
      {stage5_11[19]}
   );
   gpc1_1 gpc10590 (
      {stage4_12[16]},
      {stage5_12[10]}
   );
   gpc1_1 gpc10591 (
      {stage4_12[17]},
      {stage5_12[11]}
   );
   gpc1_1 gpc10592 (
      {stage4_12[18]},
      {stage5_12[12]}
   );
   gpc1_1 gpc10593 (
      {stage4_12[19]},
      {stage5_12[13]}
   );
   gpc1_1 gpc10594 (
      {stage4_13[26]},
      {stage5_13[7]}
   );
   gpc1_1 gpc10595 (
      {stage4_13[27]},
      {stage5_13[8]}
   );
   gpc1_1 gpc10596 (
      {stage4_14[26]},
      {stage5_14[11]}
   );
   gpc1_1 gpc10597 (
      {stage4_14[27]},
      {stage5_14[12]}
   );
   gpc1_1 gpc10598 (
      {stage4_14[28]},
      {stage5_14[13]}
   );
   gpc1_1 gpc10599 (
      {stage4_14[29]},
      {stage5_14[14]}
   );
   gpc1_1 gpc10600 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc10601 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc10602 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc10603 (
      {stage4_15[22]},
      {stage5_15[15]}
   );
   gpc1_1 gpc10604 (
      {stage4_16[27]},
      {stage5_16[8]}
   );
   gpc1_1 gpc10605 (
      {stage4_16[28]},
      {stage5_16[9]}
   );
   gpc1_1 gpc10606 (
      {stage4_16[29]},
      {stage5_16[10]}
   );
   gpc1_1 gpc10607 (
      {stage4_16[30]},
      {stage5_16[11]}
   );
   gpc1_1 gpc10608 (
      {stage4_16[31]},
      {stage5_16[12]}
   );
   gpc1_1 gpc10609 (
      {stage4_16[32]},
      {stage5_16[13]}
   );
   gpc1_1 gpc10610 (
      {stage4_19[17]},
      {stage5_19[11]}
   );
   gpc1_1 gpc10611 (
      {stage4_19[18]},
      {stage5_19[12]}
   );
   gpc1_1 gpc10612 (
      {stage4_19[19]},
      {stage5_19[13]}
   );
   gpc1_1 gpc10613 (
      {stage4_21[26]},
      {stage5_21[10]}
   );
   gpc1_1 gpc10614 (
      {stage4_23[21]},
      {stage5_23[9]}
   );
   gpc1_1 gpc10615 (
      {stage4_23[22]},
      {stage5_23[10]}
   );
   gpc1_1 gpc10616 (
      {stage4_23[23]},
      {stage5_23[11]}
   );
   gpc1_1 gpc10617 (
      {stage4_24[21]},
      {stage5_24[6]}
   );
   gpc1_1 gpc10618 (
      {stage4_24[22]},
      {stage5_24[7]}
   );
   gpc1_1 gpc10619 (
      {stage4_24[23]},
      {stage5_24[8]}
   );
   gpc1_1 gpc10620 (
      {stage4_25[15]},
      {stage5_25[8]}
   );
   gpc1_1 gpc10621 (
      {stage4_25[16]},
      {stage5_25[9]}
   );
   gpc1_1 gpc10622 (
      {stage4_25[17]},
      {stage5_25[10]}
   );
   gpc1_1 gpc10623 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc10624 (
      {stage4_25[19]},
      {stage5_25[12]}
   );
   gpc1_1 gpc10625 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc10626 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc10627 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc10628 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc10629 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc10630 (
      {stage4_26[19]},
      {stage5_26[15]}
   );
   gpc1_1 gpc10631 (
      {stage4_26[20]},
      {stage5_26[16]}
   );
   gpc1_1 gpc10632 (
      {stage4_27[17]},
      {stage5_27[5]}
   );
   gpc1_1 gpc10633 (
      {stage4_27[18]},
      {stage5_27[6]}
   );
   gpc1_1 gpc10634 (
      {stage4_27[19]},
      {stage5_27[7]}
   );
   gpc1_1 gpc10635 (
      {stage4_27[20]},
      {stage5_27[8]}
   );
   gpc1_1 gpc10636 (
      {stage4_28[29]},
      {stage5_28[9]}
   );
   gpc1_1 gpc10637 (
      {stage4_28[30]},
      {stage5_28[10]}
   );
   gpc1_1 gpc10638 (
      {stage4_28[31]},
      {stage5_28[11]}
   );
   gpc1_1 gpc10639 (
      {stage4_29[20]},
      {stage5_29[11]}
   );
   gpc1_1 gpc10640 (
      {stage4_29[21]},
      {stage5_29[12]}
   );
   gpc1_1 gpc10641 (
      {stage4_29[22]},
      {stage5_29[13]}
   );
   gpc1_1 gpc10642 (
      {stage4_29[23]},
      {stage5_29[14]}
   );
   gpc1_1 gpc10643 (
      {stage4_30[24]},
      {stage5_30[7]}
   );
   gpc1_1 gpc10644 (
      {stage4_30[25]},
      {stage5_30[8]}
   );
   gpc1_1 gpc10645 (
      {stage4_31[14]},
      {stage5_31[9]}
   );
   gpc1_1 gpc10646 (
      {stage4_31[15]},
      {stage5_31[10]}
   );
   gpc1_1 gpc10647 (
      {stage4_31[16]},
      {stage5_31[11]}
   );
   gpc1_1 gpc10648 (
      {stage4_32[20]},
      {stage5_32[11]}
   );
   gpc1_1 gpc10649 (
      {stage4_32[21]},
      {stage5_32[12]}
   );
   gpc1_1 gpc10650 (
      {stage4_32[22]},
      {stage5_32[13]}
   );
   gpc1_1 gpc10651 (
      {stage4_32[23]},
      {stage5_32[14]}
   );
   gpc1_1 gpc10652 (
      {stage4_34[18]},
      {stage5_34[9]}
   );
   gpc1_1 gpc10653 (
      {stage4_34[19]},
      {stage5_34[10]}
   );
   gpc1_1 gpc10654 (
      {stage4_34[20]},
      {stage5_34[11]}
   );
   gpc1_1 gpc10655 (
      {stage4_34[21]},
      {stage5_34[12]}
   );
   gpc1_1 gpc10656 (
      {stage4_34[22]},
      {stage5_34[13]}
   );
   gpc1_1 gpc10657 (
      {stage4_34[23]},
      {stage5_34[14]}
   );
   gpc1_1 gpc10658 (
      {stage4_34[24]},
      {stage5_34[15]}
   );
   gpc1_1 gpc10659 (
      {stage4_34[25]},
      {stage5_34[16]}
   );
   gpc1_1 gpc10660 (
      {stage4_34[26]},
      {stage5_34[17]}
   );
   gpc1_1 gpc10661 (
      {stage4_34[27]},
      {stage5_34[18]}
   );
   gpc1_1 gpc10662 (
      {stage4_34[28]},
      {stage5_34[19]}
   );
   gpc1_1 gpc10663 (
      {stage4_34[29]},
      {stage5_34[20]}
   );
   gpc1_1 gpc10664 (
      {stage4_36[33]},
      {stage5_36[14]}
   );
   gpc1_1 gpc10665 (
      {stage4_36[34]},
      {stage5_36[15]}
   );
   gpc1_1 gpc10666 (
      {stage4_36[35]},
      {stage5_36[16]}
   );
   gpc1_1 gpc10667 (
      {stage4_36[36]},
      {stage5_36[17]}
   );
   gpc1_1 gpc10668 (
      {stage4_36[37]},
      {stage5_36[18]}
   );
   gpc1_1 gpc10669 (
      {stage4_40[22]},
      {stage5_40[13]}
   );
   gpc1_1 gpc10670 (
      {stage4_40[23]},
      {stage5_40[14]}
   );
   gpc1_1 gpc10671 (
      {stage4_40[24]},
      {stage5_40[15]}
   );
   gpc1_1 gpc10672 (
      {stage4_40[25]},
      {stage5_40[16]}
   );
   gpc1_1 gpc10673 (
      {stage4_40[26]},
      {stage5_40[17]}
   );
   gpc1_1 gpc10674 (
      {stage4_40[27]},
      {stage5_40[18]}
   );
   gpc1_1 gpc10675 (
      {stage4_40[28]},
      {stage5_40[19]}
   );
   gpc1_1 gpc10676 (
      {stage4_42[19]},
      {stage5_42[10]}
   );
   gpc1_1 gpc10677 (
      {stage4_42[20]},
      {stage5_42[11]}
   );
   gpc1_1 gpc10678 (
      {stage4_42[21]},
      {stage5_42[12]}
   );
   gpc1_1 gpc10679 (
      {stage4_42[22]},
      {stage5_42[13]}
   );
   gpc1_1 gpc10680 (
      {stage4_42[23]},
      {stage5_42[14]}
   );
   gpc1_1 gpc10681 (
      {stage4_42[24]},
      {stage5_42[15]}
   );
   gpc1_1 gpc10682 (
      {stage4_42[25]},
      {stage5_42[16]}
   );
   gpc1_1 gpc10683 (
      {stage4_42[26]},
      {stage5_42[17]}
   );
   gpc1_1 gpc10684 (
      {stage4_42[27]},
      {stage5_42[18]}
   );
   gpc1_1 gpc10685 (
      {stage4_42[28]},
      {stage5_42[19]}
   );
   gpc1_1 gpc10686 (
      {stage4_44[26]},
      {stage5_44[12]}
   );
   gpc1_1 gpc10687 (
      {stage4_44[27]},
      {stage5_44[13]}
   );
   gpc1_1 gpc10688 (
      {stage4_44[28]},
      {stage5_44[14]}
   );
   gpc1_1 gpc10689 (
      {stage4_44[29]},
      {stage5_44[15]}
   );
   gpc1_1 gpc10690 (
      {stage4_44[30]},
      {stage5_44[16]}
   );
   gpc1_1 gpc10691 (
      {stage4_44[31]},
      {stage5_44[17]}
   );
   gpc1_1 gpc10692 (
      {stage4_44[32]},
      {stage5_44[18]}
   );
   gpc1_1 gpc10693 (
      {stage4_44[33]},
      {stage5_44[19]}
   );
   gpc1_1 gpc10694 (
      {stage4_44[34]},
      {stage5_44[20]}
   );
   gpc1_1 gpc10695 (
      {stage4_44[35]},
      {stage5_44[21]}
   );
   gpc1_1 gpc10696 (
      {stage4_44[36]},
      {stage5_44[22]}
   );
   gpc1_1 gpc10697 (
      {stage4_44[37]},
      {stage5_44[23]}
   );
   gpc1_1 gpc10698 (
      {stage4_44[38]},
      {stage5_44[24]}
   );
   gpc1_1 gpc10699 (
      {stage4_44[39]},
      {stage5_44[25]}
   );
   gpc1_1 gpc10700 (
      {stage4_48[11]},
      {stage5_48[7]}
   );
   gpc1_1 gpc10701 (
      {stage4_48[12]},
      {stage5_48[8]}
   );
   gpc1_1 gpc10702 (
      {stage4_48[13]},
      {stage5_48[9]}
   );
   gpc1_1 gpc10703 (
      {stage4_48[14]},
      {stage5_48[10]}
   );
   gpc1_1 gpc10704 (
      {stage4_48[15]},
      {stage5_48[11]}
   );
   gpc1_1 gpc10705 (
      {stage4_48[16]},
      {stage5_48[12]}
   );
   gpc1_1 gpc10706 (
      {stage4_48[17]},
      {stage5_48[13]}
   );
   gpc1_1 gpc10707 (
      {stage4_48[18]},
      {stage5_48[14]}
   );
   gpc1_1 gpc10708 (
      {stage4_48[19]},
      {stage5_48[15]}
   );
   gpc1_1 gpc10709 (
      {stage4_48[20]},
      {stage5_48[16]}
   );
   gpc1_1 gpc10710 (
      {stage4_48[21]},
      {stage5_48[17]}
   );
   gpc1_1 gpc10711 (
      {stage4_49[18]},
      {stage5_49[7]}
   );
   gpc1_1 gpc10712 (
      {stage4_49[19]},
      {stage5_49[8]}
   );
   gpc1_1 gpc10713 (
      {stage4_49[20]},
      {stage5_49[9]}
   );
   gpc1_1 gpc10714 (
      {stage4_49[21]},
      {stage5_49[10]}
   );
   gpc1_1 gpc10715 (
      {stage4_49[22]},
      {stage5_49[11]}
   );
   gpc1_1 gpc10716 (
      {stage4_49[23]},
      {stage5_49[12]}
   );
   gpc1_1 gpc10717 (
      {stage4_49[24]},
      {stage5_49[13]}
   );
   gpc1_1 gpc10718 (
      {stage4_49[25]},
      {stage5_49[14]}
   );
   gpc1_1 gpc10719 (
      {stage4_49[26]},
      {stage5_49[15]}
   );
   gpc1_1 gpc10720 (
      {stage4_49[27]},
      {stage5_49[16]}
   );
   gpc1_1 gpc10721 (
      {stage4_52[19]},
      {stage5_52[9]}
   );
   gpc1_1 gpc10722 (
      {stage4_52[20]},
      {stage5_52[10]}
   );
   gpc1_1 gpc10723 (
      {stage4_52[21]},
      {stage5_52[11]}
   );
   gpc1_1 gpc10724 (
      {stage4_52[22]},
      {stage5_52[12]}
   );
   gpc1_1 gpc10725 (
      {stage4_53[25]},
      {stage5_53[8]}
   );
   gpc1_1 gpc10726 (
      {stage4_53[26]},
      {stage5_53[9]}
   );
   gpc1_1 gpc10727 (
      {stage4_53[27]},
      {stage5_53[10]}
   );
   gpc1_1 gpc10728 (
      {stage4_53[28]},
      {stage5_53[11]}
   );
   gpc1_1 gpc10729 (
      {stage4_54[26]},
      {stage5_54[12]}
   );
   gpc1_1 gpc10730 (
      {stage4_54[27]},
      {stage5_54[13]}
   );
   gpc1_1 gpc10731 (
      {stage4_54[28]},
      {stage5_54[14]}
   );
   gpc1_1 gpc10732 (
      {stage4_54[29]},
      {stage5_54[15]}
   );
   gpc1_1 gpc10733 (
      {stage4_54[30]},
      {stage5_54[16]}
   );
   gpc1_1 gpc10734 (
      {stage4_55[22]},
      {stage5_55[11]}
   );
   gpc1_1 gpc10735 (
      {stage4_55[23]},
      {stage5_55[12]}
   );
   gpc1_1 gpc10736 (
      {stage4_55[24]},
      {stage5_55[13]}
   );
   gpc1_1 gpc10737 (
      {stage4_55[25]},
      {stage5_55[14]}
   );
   gpc1_1 gpc10738 (
      {stage4_55[26]},
      {stage5_55[15]}
   );
   gpc1_1 gpc10739 (
      {stage4_55[27]},
      {stage5_55[16]}
   );
   gpc1_1 gpc10740 (
      {stage4_55[28]},
      {stage5_55[17]}
   );
   gpc1_1 gpc10741 (
      {stage4_56[24]},
      {stage5_56[8]}
   );
   gpc1_1 gpc10742 (
      {stage4_56[25]},
      {stage5_56[9]}
   );
   gpc1_1 gpc10743 (
      {stage4_56[26]},
      {stage5_56[10]}
   );
   gpc1_1 gpc10744 (
      {stage4_56[27]},
      {stage5_56[11]}
   );
   gpc1_1 gpc10745 (
      {stage4_56[28]},
      {stage5_56[12]}
   );
   gpc1_1 gpc10746 (
      {stage4_58[0]},
      {stage5_58[8]}
   );
   gpc1_1 gpc10747 (
      {stage4_58[1]},
      {stage5_58[9]}
   );
   gpc1_1 gpc10748 (
      {stage4_58[2]},
      {stage5_58[10]}
   );
   gpc1_1 gpc10749 (
      {stage4_58[3]},
      {stage5_58[11]}
   );
   gpc1_1 gpc10750 (
      {stage4_58[4]},
      {stage5_58[12]}
   );
   gpc1_1 gpc10751 (
      {stage4_58[5]},
      {stage5_58[13]}
   );
   gpc1_1 gpc10752 (
      {stage4_58[6]},
      {stage5_58[14]}
   );
   gpc1_1 gpc10753 (
      {stage4_58[7]},
      {stage5_58[15]}
   );
   gpc1_1 gpc10754 (
      {stage4_58[8]},
      {stage5_58[16]}
   );
   gpc1_1 gpc10755 (
      {stage4_58[9]},
      {stage5_58[17]}
   );
   gpc1_1 gpc10756 (
      {stage4_58[10]},
      {stage5_58[18]}
   );
   gpc1_1 gpc10757 (
      {stage4_58[11]},
      {stage5_58[19]}
   );
   gpc1_1 gpc10758 (
      {stage4_58[12]},
      {stage5_58[20]}
   );
   gpc1_1 gpc10759 (
      {stage4_58[13]},
      {stage5_58[21]}
   );
   gpc1_1 gpc10760 (
      {stage4_58[14]},
      {stage5_58[22]}
   );
   gpc1_1 gpc10761 (
      {stage4_58[15]},
      {stage5_58[23]}
   );
   gpc1_1 gpc10762 (
      {stage4_60[18]},
      {stage5_60[7]}
   );
   gpc1_1 gpc10763 (
      {stage4_60[19]},
      {stage5_60[8]}
   );
   gpc1_1 gpc10764 (
      {stage4_60[20]},
      {stage5_60[9]}
   );
   gpc1_1 gpc10765 (
      {stage4_60[21]},
      {stage5_60[10]}
   );
   gpc1_1 gpc10766 (
      {stage4_60[22]},
      {stage5_60[11]}
   );
   gpc1_1 gpc10767 (
      {stage4_60[23]},
      {stage5_60[12]}
   );
   gpc1_1 gpc10768 (
      {stage4_60[24]},
      {stage5_60[13]}
   );
   gpc1_1 gpc10769 (
      {stage4_61[26]},
      {stage5_61[7]}
   );
   gpc1_1 gpc10770 (
      {stage4_61[27]},
      {stage5_61[8]}
   );
   gpc1_1 gpc10771 (
      {stage4_61[28]},
      {stage5_61[9]}
   );
   gpc1_1 gpc10772 (
      {stage4_64[16]},
      {stage5_64[9]}
   );
   gpc1_1 gpc10773 (
      {stage4_64[17]},
      {stage5_64[10]}
   );
   gpc1_1 gpc10774 (
      {stage4_64[18]},
      {stage5_64[11]}
   );
   gpc1_1 gpc10775 (
      {stage4_64[19]},
      {stage5_64[12]}
   );
   gpc1_1 gpc10776 (
      {stage4_64[20]},
      {stage5_64[13]}
   );
   gpc1_1 gpc10777 (
      {stage4_64[21]},
      {stage5_64[14]}
   );
   gpc1_1 gpc10778 (
      {stage4_64[22]},
      {stage5_64[15]}
   );
   gpc1_1 gpc10779 (
      {stage4_64[23]},
      {stage5_64[16]}
   );
   gpc1_1 gpc10780 (
      {stage4_64[24]},
      {stage5_64[17]}
   );
   gpc1_1 gpc10781 (
      {stage4_64[25]},
      {stage5_64[18]}
   );
   gpc1_1 gpc10782 (
      {stage4_64[26]},
      {stage5_64[19]}
   );
   gpc1_1 gpc10783 (
      {stage4_66[11]},
      {stage5_66[9]}
   );
   gpc1_1 gpc10784 (
      {stage4_66[12]},
      {stage5_66[10]}
   );
   gpc1_1 gpc10785 (
      {stage4_66[13]},
      {stage5_66[11]}
   );
   gpc1_1 gpc10786 (
      {stage4_66[14]},
      {stage5_66[12]}
   );
   gpc1_1 gpc10787 (
      {stage4_68[3]},
      {stage5_68[3]}
   );
   gpc1_1 gpc10788 (
      {stage4_68[4]},
      {stage5_68[4]}
   );
   gpc1_1 gpc10789 (
      {stage4_68[5]},
      {stage5_68[5]}
   );
   gpc1_1 gpc10790 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc10791 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc10792 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc10793 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc10794 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc10795 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc10796 (
      {stage4_70[0]},
      {stage5_70[3]}
   );
   gpc615_5 gpc10797 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc207_4 gpc10798 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc10799 (
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc606_5 gpc10800 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], stage5_5[16], stage5_5[17]},
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10], 1'b0},
      {stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc117_4 gpc10801 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {1'b0},
      {stage5_8[0]},
      {stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[4]}
   );
   gpc615_5 gpc10802 (
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12], stage5_6[13]},
      {1'b0},
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[5],stage6_6[5]}
   );
   gpc606_5 gpc10803 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[4],stage6_8[4]}
   );
   gpc606_5 gpc10804 (
      {stage5_8[13], stage5_8[14], stage5_8[15], 1'b0, 1'b0, 1'b0},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], 1'b0, 1'b0},
      {stage6_12[1],stage6_11[1],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc207_4 gpc10805 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5], stage5_9[6]},
      {stage5_11[0], stage5_11[1]},
      {stage6_12[2],stage6_11[2],stage6_10[3],stage6_9[6]}
   );
   gpc606_5 gpc10806 (
      {stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11], stage5_9[12]},
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7]},
      {stage6_13[0],stage6_12[3],stage6_11[3],stage6_10[4],stage6_9[7]}
   );
   gpc1406_5 gpc10807 (
      {stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[4],stage6_11[4]}
   );
   gpc1406_5 gpc10808 (
      {stage5_11[14], stage5_11[15], stage5_11[16], stage5_11[17], stage5_11[18], stage5_11[19]},
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7]},
      {stage5_14[1]},
      {stage6_15[1],stage6_14[1],stage6_13[2],stage6_12[5],stage6_11[5]}
   );
   gpc117_4 gpc10809 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage5_13[8]},
      {stage5_14[2]},
      {stage6_15[2],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc117_4 gpc10810 (
      {stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {1'b0},
      {stage5_14[3]},
      {stage6_15[3],stage6_14[3],stage6_13[4],stage6_12[7]}
   );
   gpc1343_5 gpc10811 (
      {stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[4],stage6_14[4]}
   );
   gpc1343_5 gpc10812 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[5],stage6_14[5]}
   );
   gpc1343_5 gpc10813 (
      {stage5_14[10], stage5_14[11], stage5_14[12]},
      {stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage5_16[6], stage5_16[7], stage5_16[8]},
      {stage5_17[2]},
      {stage6_18[2],stage6_17[2],stage6_16[2],stage6_15[6],stage6_14[6]}
   );
   gpc1343_5 gpc10814 (
      {stage5_14[13], stage5_14[14], 1'b0},
      {stage5_15[12], stage5_15[13], stage5_15[14], stage5_15[15]},
      {stage5_16[9], stage5_16[10], stage5_16[11]},
      {stage5_17[3]},
      {stage6_18[3],stage6_17[3],stage6_16[3],stage6_15[7],stage6_14[7]}
   );
   gpc207_4 gpc10815 (
      {stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7], 1'b0, 1'b0, 1'b0},
      {stage5_19[0], stage5_19[1]},
      {stage6_20[0],stage6_19[0],stage6_18[4],stage6_17[4]}
   );
   gpc7_3 gpc10816 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage6_20[1],stage6_19[1],stage6_18[5]}
   );
   gpc7_3 gpc10817 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13]},
      {stage6_20[2],stage6_19[2],stage6_18[6]}
   );
   gpc2135_5 gpc10818 (
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[3],stage6_19[3]}
   );
   gpc7_3 gpc10819 (
      {stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13]},
      {stage6_21[1],stage6_20[4],stage6_19[4]}
   );
   gpc1415_5 gpc10820 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_21[1]},
      {stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[2],stage6_20[5]}
   );
   gpc207_4 gpc10821 (
      {stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5], stage5_21[6], stage5_21[7], stage5_21[8]},
      {stage5_23[1], stage5_23[2]},
      {stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[3]}
   );
   gpc606_5 gpc10822 (
      {stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[3]}
   );
   gpc606_5 gpc10823 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3]}
   );
   gpc1343_5 gpc10824 (
      {stage5_26[6], stage5_26[7], stage5_26[8]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[2],stage6_26[2]}
   );
   gpc1343_5 gpc10825 (
      {stage5_26[9], stage5_26[10], stage5_26[11]},
      {stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage5_29[1]},
      {stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc10826 (
      {stage5_26[12], stage5_26[13], stage5_26[14], stage5_26[15], stage5_26[16]},
      {stage5_27[8]},
      {stage5_28[6], stage5_28[7], stage5_28[8], stage5_28[9], stage5_28[10], stage5_28[11]},
      {stage6_30[2],stage6_29[2],stage6_28[3],stage6_27[4],stage6_26[4]}
   );
   gpc606_5 gpc10827 (
      {stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6], stage5_29[7]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[3],stage6_29[3]}
   );
   gpc606_5 gpc10828 (
      {stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11], stage5_29[12], stage5_29[13]},
      {stage5_31[6], stage5_31[7], stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11]},
      {stage6_33[1],stage6_32[1],stage6_31[1],stage6_30[4],stage6_29[4]}
   );
   gpc7_3 gpc10829 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage6_32[2],stage6_31[2],stage6_30[5]}
   );
   gpc1415_5 gpc10830 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4]},
      {stage5_33[0]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3]},
      {stage5_35[0]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[2],stage6_32[3]}
   );
   gpc1415_5 gpc10831 (
      {stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage5_33[1]},
      {stage5_34[4], stage5_34[5], stage5_34[6], stage5_34[7]},
      {stage5_35[1]},
      {stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[3],stage6_32[4]}
   );
   gpc606_5 gpc10832 (
      {stage5_32[10], stage5_32[11], stage5_32[12], stage5_32[13], stage5_32[14], 1'b0},
      {stage5_34[8], stage5_34[9], stage5_34[10], stage5_34[11], stage5_34[12], stage5_34[13]},
      {stage6_36[2],stage6_35[2],stage6_34[2],stage6_33[4],stage6_32[5]}
   );
   gpc615_5 gpc10833 (
      {stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_34[14]},
      {stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5], stage5_35[6], stage5_35[7]},
      {stage6_37[0],stage6_36[3],stage6_35[3],stage6_34[3],stage6_33[5]}
   );
   gpc615_5 gpc10834 (
      {stage5_34[15], stage5_34[16], stage5_34[17], stage5_34[18], stage5_34[19]},
      {stage5_35[8]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[4],stage6_35[4],stage6_34[4]}
   );
   gpc2135_5 gpc10835 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10]},
      {stage5_37[0], stage5_37[1], stage5_37[2]},
      {stage5_38[0]},
      {stage5_39[0], stage5_39[1]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[2],stage6_36[5]}
   );
   gpc2135_5 gpc10836 (
      {stage5_36[11], stage5_36[12], stage5_36[13], stage5_36[14], stage5_36[15]},
      {stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage5_38[1]},
      {stage5_39[2], stage5_39[3]},
      {stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[3],stage6_36[6]}
   );
   gpc606_5 gpc10837 (
      {stage5_36[16], stage5_36[17], stage5_36[18], 1'b0, 1'b0, 1'b0},
      {stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5], stage5_38[6], 1'b0},
      {stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[4],stage6_36[7]}
   );
   gpc606_5 gpc10838 (
      {stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10], 1'b0},
      {stage5_39[4], stage5_39[5], stage5_39[6], stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage6_41[0],stage6_40[3],stage6_39[3],stage6_38[4],stage6_37[5]}
   );
   gpc606_5 gpc10839 (
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[1],stage6_40[4]}
   );
   gpc606_5 gpc10840 (
      {stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9], stage5_40[10], stage5_40[11]},
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10], stage5_42[11]},
      {stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[2],stage6_40[5]}
   );
   gpc1325_5 gpc10841 (
      {stage5_40[12], stage5_40[13], stage5_40[14], stage5_40[15], stage5_40[16]},
      {stage5_41[0], stage5_41[1]},
      {stage5_42[12], stage5_42[13], stage5_42[14]},
      {stage5_43[0]},
      {stage6_44[2],stage6_43[2],stage6_42[2],stage6_41[3],stage6_40[6]}
   );
   gpc615_5 gpc10842 (
      {stage5_42[15], stage5_42[16], stage5_42[17], stage5_42[18], stage5_42[19]},
      {stage5_43[1]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[0],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc7_3 gpc10843 (
      {stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5], stage5_43[6], stage5_43[7], 1'b0},
      {stage6_45[1],stage6_44[4],stage6_43[4]}
   );
   gpc7_3 gpc10844 (
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11], stage5_44[12]},
      {stage6_46[1],stage6_45[2],stage6_44[5]}
   );
   gpc7_3 gpc10845 (
      {stage5_44[13], stage5_44[14], stage5_44[15], stage5_44[16], stage5_44[17], stage5_44[18], stage5_44[19]},
      {stage6_46[2],stage6_45[3],stage6_44[6]}
   );
   gpc606_5 gpc10846 (
      {stage5_44[20], stage5_44[21], stage5_44[22], stage5_44[23], stage5_44[24], stage5_44[25]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[3],stage6_45[4],stage6_44[7]}
   );
   gpc606_5 gpc10847 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc10848 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], 1'b0, 1'b0},
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10], stage5_47[11]},
      {stage6_49[1],stage6_48[2],stage6_47[2],stage6_46[5],stage6_45[6]}
   );
   gpc615_5 gpc10849 (
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10]},
      {stage5_47[12]},
      {stage5_48[0], stage5_48[1], stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5]},
      {stage6_50[0],stage6_49[2],stage6_48[3],stage6_47[3],stage6_46[6]}
   );
   gpc606_5 gpc10850 (
      {stage5_48[6], stage5_48[7], stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[1],stage6_49[3],stage6_48[4]}
   );
   gpc606_5 gpc10851 (
      {stage5_48[12], stage5_48[13], stage5_48[14], stage5_48[15], stage5_48[16], stage5_48[17]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], 1'b0, 1'b0},
      {stage6_52[1],stage6_51[1],stage6_50[2],stage6_49[4],stage6_48[5]}
   );
   gpc207_4 gpc10852 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5], stage5_49[6]},
      {stage5_51[0], stage5_51[1]},
      {stage6_52[2],stage6_51[2],stage6_50[3],stage6_49[5]}
   );
   gpc207_4 gpc10853 (
      {stage5_49[7], stage5_49[8], stage5_49[9], stage5_49[10], stage5_49[11], stage5_49[12], stage5_49[13]},
      {stage5_51[2], stage5_51[3]},
      {stage6_52[3],stage6_51[3],stage6_50[4],stage6_49[6]}
   );
   gpc606_5 gpc10854 (
      {stage5_51[4], stage5_51[5], stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[0],stage6_52[4],stage6_51[4]}
   );
   gpc606_5 gpc10855 (
      {stage5_52[0], stage5_52[1], stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5]},
      {stage5_54[0], stage5_54[1], stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5]},
      {stage6_56[0],stage6_55[1],stage6_54[1],stage6_53[1],stage6_52[5]}
   );
   gpc606_5 gpc10856 (
      {stage5_52[6], stage5_52[7], stage5_52[8], stage5_52[9], stage5_52[10], stage5_52[11]},
      {stage5_54[6], stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage6_56[1],stage6_55[2],stage6_54[2],stage6_53[2],stage6_52[6]}
   );
   gpc606_5 gpc10857 (
      {stage5_53[6], stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11]},
      {stage5_55[0], stage5_55[1], stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5]},
      {stage6_57[0],stage6_56[2],stage6_55[3],stage6_54[3],stage6_53[3]}
   );
   gpc1163_5 gpc10858 (
      {stage5_54[12], stage5_54[13], stage5_54[14]},
      {stage5_55[6], stage5_55[7], stage5_55[8], stage5_55[9], stage5_55[10], stage5_55[11]},
      {stage5_56[0]},
      {stage5_57[0]},
      {stage6_58[0],stage6_57[1],stage6_56[3],stage6_55[4],stage6_54[4]}
   );
   gpc1163_5 gpc10859 (
      {stage5_54[15], stage5_54[16], 1'b0},
      {stage5_55[12], stage5_55[13], stage5_55[14], stage5_55[15], stage5_55[16], stage5_55[17]},
      {stage5_56[1]},
      {stage5_57[1]},
      {stage6_58[1],stage6_57[2],stage6_56[4],stage6_55[5],stage6_54[5]}
   );
   gpc606_5 gpc10860 (
      {stage5_56[2], stage5_56[3], stage5_56[4], stage5_56[5], stage5_56[6], stage5_56[7]},
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage6_60[0],stage6_59[0],stage6_58[2],stage6_57[3],stage6_56[5]}
   );
   gpc606_5 gpc10861 (
      {stage5_56[8], stage5_56[9], stage5_56[10], stage5_56[11], stage5_56[12], 1'b0},
      {stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9], stage5_58[10], stage5_58[11]},
      {stage6_60[1],stage6_59[1],stage6_58[3],stage6_57[4],stage6_56[6]}
   );
   gpc606_5 gpc10862 (
      {stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5], stage5_57[6], stage5_57[7]},
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage6_61[0],stage6_60[2],stage6_59[2],stage6_58[4],stage6_57[5]}
   );
   gpc606_5 gpc10863 (
      {stage5_58[12], stage5_58[13], stage5_58[14], stage5_58[15], stage5_58[16], stage5_58[17]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[1],stage6_60[3],stage6_59[3],stage6_58[5]}
   );
   gpc606_5 gpc10864 (
      {stage5_58[18], stage5_58[19], stage5_58[20], stage5_58[21], stage5_58[22], stage5_58[23]},
      {stage5_60[6], stage5_60[7], stage5_60[8], stage5_60[9], stage5_60[10], stage5_60[11]},
      {stage6_62[1],stage6_61[2],stage6_60[4],stage6_59[4],stage6_58[6]}
   );
   gpc1343_5 gpc10865 (
      {stage5_61[0], stage5_61[1], stage5_61[2]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3]},
      {stage5_63[0], stage5_63[1], stage5_63[2]},
      {stage5_64[0]},
      {stage6_65[0],stage6_64[0],stage6_63[0],stage6_62[2],stage6_61[3]}
   );
   gpc1343_5 gpc10866 (
      {stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage5_62[4], stage5_62[5], stage5_62[6], stage5_62[7]},
      {stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage5_64[1]},
      {stage6_65[1],stage6_64[1],stage6_63[1],stage6_62[3],stage6_61[4]}
   );
   gpc606_5 gpc10867 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], 1'b0, 1'b0},
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], 1'b0},
      {stage6_65[2],stage6_64[2],stage6_63[2],stage6_62[4],stage6_61[5]}
   );
   gpc117_4 gpc10868 (
      {stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5], stage5_64[6], stage5_64[7], stage5_64[8]},
      {stage5_65[0]},
      {stage5_66[0]},
      {stage6_67[0],stage6_66[0],stage6_65[3],stage6_64[3]}
   );
   gpc606_5 gpc10869 (
      {stage5_64[9], stage5_64[10], stage5_64[11], stage5_64[12], stage5_64[13], stage5_64[14]},
      {stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], stage5_66[5], stage5_66[6]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[4],stage6_64[4]}
   );
   gpc615_5 gpc10870 (
      {stage5_64[15], stage5_64[16], stage5_64[17], stage5_64[18], stage5_64[19]},
      {stage5_65[1]},
      {stage5_66[7], stage5_66[8], stage5_66[9], stage5_66[10], stage5_66[11], stage5_66[12]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[5],stage6_64[5]}
   );
   gpc2135_5 gpc10871 (
      {stage5_67[0], stage5_67[1], stage5_67[2], stage5_67[3], stage5_67[4]},
      {stage5_68[0], stage5_68[1], stage5_68[2]},
      {stage5_69[0]},
      {stage5_70[0], stage5_70[1]},
      {stage6_71[0],stage6_70[0],stage6_69[0],stage6_68[2],stage6_67[3]}
   );
   gpc2135_5 gpc10872 (
      {stage5_67[5], stage5_67[6], stage5_67[7], 1'b0, 1'b0},
      {stage5_68[3], stage5_68[4], stage5_68[5]},
      {stage5_69[1]},
      {stage5_70[2], stage5_70[3]},
      {stage6_71[1],stage6_70[1],stage6_69[1],stage6_68[3],stage6_67[4]}
   );
   gpc1_1 gpc10873 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc10874 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc10875 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc10876 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc10877 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc10878 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc10879 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc10880 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc10881 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc10882 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc10883 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc10884 (
      {stage5_3[5]},
      {stage6_3[1]}
   );
   gpc1_1 gpc10885 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc10886 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc10887 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc10888 (
      {stage5_5[18]},
      {stage6_5[4]}
   );
   gpc1_1 gpc10889 (
      {stage5_5[19]},
      {stage6_5[5]}
   );
   gpc1_1 gpc10890 (
      {stage5_5[20]},
      {stage6_5[6]}
   );
   gpc1_1 gpc10891 (
      {stage5_16[12]},
      {stage6_16[4]}
   );
   gpc1_1 gpc10892 (
      {stage5_16[13]},
      {stage6_16[5]}
   );
   gpc1_1 gpc10893 (
      {stage5_21[9]},
      {stage6_21[4]}
   );
   gpc1_1 gpc10894 (
      {stage5_21[10]},
      {stage6_21[5]}
   );
   gpc1_1 gpc10895 (
      {stage5_22[6]},
      {stage6_22[3]}
   );
   gpc1_1 gpc10896 (
      {stage5_22[7]},
      {stage6_22[4]}
   );
   gpc1_1 gpc10897 (
      {stage5_22[8]},
      {stage6_22[5]}
   );
   gpc1_1 gpc10898 (
      {stage5_22[9]},
      {stage6_22[6]}
   );
   gpc1_1 gpc10899 (
      {stage5_22[10]},
      {stage6_22[7]}
   );
   gpc1_1 gpc10900 (
      {stage5_22[11]},
      {stage6_22[8]}
   );
   gpc1_1 gpc10901 (
      {stage5_22[12]},
      {stage6_22[9]}
   );
   gpc1_1 gpc10902 (
      {stage5_22[13]},
      {stage6_22[10]}
   );
   gpc1_1 gpc10903 (
      {stage5_22[14]},
      {stage6_22[11]}
   );
   gpc1_1 gpc10904 (
      {stage5_23[9]},
      {stage6_23[4]}
   );
   gpc1_1 gpc10905 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc10906 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc10907 (
      {stage5_24[6]},
      {stage6_24[4]}
   );
   gpc1_1 gpc10908 (
      {stage5_24[7]},
      {stage6_24[5]}
   );
   gpc1_1 gpc10909 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc10910 (
      {stage5_25[6]},
      {stage6_25[2]}
   );
   gpc1_1 gpc10911 (
      {stage5_25[7]},
      {stage6_25[3]}
   );
   gpc1_1 gpc10912 (
      {stage5_25[8]},
      {stage6_25[4]}
   );
   gpc1_1 gpc10913 (
      {stage5_25[9]},
      {stage6_25[5]}
   );
   gpc1_1 gpc10914 (
      {stage5_25[10]},
      {stage6_25[6]}
   );
   gpc1_1 gpc10915 (
      {stage5_25[11]},
      {stage6_25[7]}
   );
   gpc1_1 gpc10916 (
      {stage5_25[12]},
      {stage6_25[8]}
   );
   gpc1_1 gpc10917 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc10918 (
      {stage5_30[7]},
      {stage6_30[6]}
   );
   gpc1_1 gpc10919 (
      {stage5_30[8]},
      {stage6_30[7]}
   );
   gpc1_1 gpc10920 (
      {stage5_33[7]},
      {stage6_33[6]}
   );
   gpc1_1 gpc10921 (
      {stage5_33[8]},
      {stage6_33[7]}
   );
   gpc1_1 gpc10922 (
      {stage5_34[20]},
      {stage6_34[5]}
   );
   gpc1_1 gpc10923 (
      {stage5_39[10]},
      {stage6_39[4]}
   );
   gpc1_1 gpc10924 (
      {stage5_40[17]},
      {stage6_40[7]}
   );
   gpc1_1 gpc10925 (
      {stage5_40[18]},
      {stage6_40[8]}
   );
   gpc1_1 gpc10926 (
      {stage5_40[19]},
      {stage6_40[9]}
   );
   gpc1_1 gpc10927 (
      {stage5_41[2]},
      {stage6_41[4]}
   );
   gpc1_1 gpc10928 (
      {stage5_41[3]},
      {stage6_41[5]}
   );
   gpc1_1 gpc10929 (
      {stage5_41[4]},
      {stage6_41[6]}
   );
   gpc1_1 gpc10930 (
      {stage5_41[5]},
      {stage6_41[7]}
   );
   gpc1_1 gpc10931 (
      {stage5_41[6]},
      {stage6_41[8]}
   );
   gpc1_1 gpc10932 (
      {stage5_41[7]},
      {stage6_41[9]}
   );
   gpc1_1 gpc10933 (
      {stage5_41[8]},
      {stage6_41[10]}
   );
   gpc1_1 gpc10934 (
      {stage5_49[14]},
      {stage6_49[7]}
   );
   gpc1_1 gpc10935 (
      {stage5_49[15]},
      {stage6_49[8]}
   );
   gpc1_1 gpc10936 (
      {stage5_49[16]},
      {stage6_49[9]}
   );
   gpc1_1 gpc10937 (
      {stage5_52[12]},
      {stage6_52[7]}
   );
   gpc1_1 gpc10938 (
      {stage5_57[8]},
      {stage6_57[6]}
   );
   gpc1_1 gpc10939 (
      {stage5_60[12]},
      {stage6_60[5]}
   );
   gpc1_1 gpc10940 (
      {stage5_60[13]},
      {stage6_60[6]}
   );
   gpc1_1 gpc10941 (
      {stage5_65[2]},
      {stage6_65[6]}
   );
   gpc1_1 gpc10942 (
      {stage5_65[3]},
      {stage6_65[7]}
   );
   gpc1_1 gpc10943 (
      {stage5_65[4]},
      {stage6_65[8]}
   );
   gpc1_1 gpc10944 (
      {stage5_65[5]},
      {stage6_65[9]}
   );
   gpc1_1 gpc10945 (
      {stage5_68[6]},
      {stage6_68[4]}
   );
   gpc1_1 gpc10946 (
      {stage5_68[7]},
      {stage6_68[5]}
   );
   gpc1_1 gpc10947 (
      {stage5_68[8]},
      {stage6_68[6]}
   );
   gpc1_1 gpc10948 (
      {stage5_68[9]},
      {stage6_68[7]}
   );
   gpc1_1 gpc10949 (
      {stage5_68[10]},
      {stage6_68[8]}
   );
   gpc1_1 gpc10950 (
      {stage5_68[11]},
      {stage6_68[9]}
   );
   gpc1_1 gpc10951 (
      {stage5_69[2]},
      {stage6_69[2]}
   );
   gpc135_4 gpc10952 (
      {stage6_4[0], stage6_4[1], stage6_4[2], 1'b0, 1'b0},
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc615_5 gpc10953 (
      {stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_7[0]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1],stage7_6[1]}
   );
   gpc15_3 gpc10954 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc623_5 gpc10955 (
      {stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[2]}
   );
   gpc23_3 gpc10956 (
      {stage6_11[2], stage6_11[3], stage6_11[4]},
      {stage6_12[6], stage6_12[7]},
      {stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc117_4 gpc10957 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage6_15[0]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1]}
   );
   gpc7_3 gpc10958 (
      {stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5], stage6_15[6], stage6_15[7]},
      {stage7_17[1],stage7_16[1],stage7_15[1]}
   );
   gpc15_3 gpc10959 (
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4]},
      {stage6_18[0]},
      {stage7_19[0],stage7_18[0],stage7_17[2]}
   );
   gpc606_5 gpc10960 (
      {stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5], stage6_18[6]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[1],stage7_18[1]}
   );
   gpc1163_5 gpc10961 (
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_23[0]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1]}
   );
   gpc1163_5 gpc10962 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[6], stage6_22[7], stage6_22[8], stage6_22[9], stage6_22[10], stage6_22[11]},
      {stage6_23[1]},
      {stage6_24[1]},
      {stage7_25[1],stage7_24[1],stage7_23[1],stage7_22[2],stage7_21[2]}
   );
   gpc15_3 gpc10963 (
      {stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5], stage6_24[6]},
      {stage6_25[0]},
      {stage7_26[0],stage7_25[2],stage7_24[2]}
   );
   gpc606_5 gpc10964 (
      {stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5], stage6_25[6]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], 1'b0},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[3]}
   );
   gpc606_5 gpc10965 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], 1'b0, 1'b0},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[1]}
   );
   gpc1406_5 gpc10966 (
      {stage6_29[0], stage6_29[1], stage6_29[2], stage6_29[3], stage6_29[4], stage6_29[5]},
      {stage6_31[0], stage6_31[1], stage6_31[2], 1'b0},
      {stage6_32[0]},
      {stage7_33[0],stage7_32[1],stage7_31[1],stage7_30[1],stage7_29[2]}
   );
   gpc135_4 gpc10967 (
      {stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage6_33[0], stage6_33[1], stage6_33[2]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[1],stage7_32[2]}
   );
   gpc15_3 gpc10968 (
      {stage6_33[3], stage6_33[4], stage6_33[5], stage6_33[6], stage6_33[7]},
      {stage6_34[1]},
      {stage7_35[1],stage7_34[1],stage7_33[2]}
   );
   gpc117_4 gpc10969 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage6_37[0]},
      {stage6_38[0]},
      {stage7_39[0],stage7_38[0],stage7_37[0],stage7_36[0]}
   );
   gpc15_3 gpc10970 (
      {stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_38[1]},
      {stage7_39[1],stage7_38[1],stage7_37[1]}
   );
   gpc3_2 gpc10971 (
      {stage6_38[2], stage6_38[3], stage6_38[4]},
      {stage7_39[2],stage7_38[2]}
   );
   gpc2135_5 gpc10972 (
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], stage6_39[4]},
      {stage6_40[0], stage6_40[1], stage6_40[2]},
      {stage6_41[0]},
      {stage6_42[0], stage6_42[1]},
      {stage7_43[0],stage7_42[0],stage7_41[0],stage7_40[0],stage7_39[3]}
   );
   gpc207_4 gpc10973 (
      {stage6_40[3], stage6_40[4], stage6_40[5], stage6_40[6], stage6_40[7], stage6_40[8], stage6_40[9]},
      {stage6_42[2], stage6_42[3]},
      {stage7_43[1],stage7_42[1],stage7_41[1],stage7_40[1]}
   );
   gpc7_3 gpc10974 (
      {stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4], stage6_41[5], stage6_41[6], stage6_41[7]},
      {stage7_43[2],stage7_42[2],stage7_41[2]}
   );
   gpc215_4 gpc10975 (
      {stage6_43[0], stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4]},
      {stage6_44[0]},
      {stage6_45[0], stage6_45[1]},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[3]}
   );
   gpc207_4 gpc10976 (
      {stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], stage6_44[5], stage6_44[6], stage6_44[7]},
      {stage6_46[0], stage6_46[1]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1]}
   );
   gpc615_5 gpc10977 (
      {stage6_47[0], stage6_47[1], stage6_47[2], stage6_47[3], 1'b0},
      {stage6_48[0]},
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage7_51[0],stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1]}
   );
   gpc7_3 gpc10978 (
      {stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5], 1'b0, 1'b0},
      {stage7_50[1],stage7_49[1],stage7_48[1]}
   );
   gpc615_5 gpc10979 (
      {stage6_50[0], stage6_50[1], stage6_50[2], stage6_50[3], stage6_50[4]},
      {stage6_51[0]},
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4], stage6_52[5]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[2]}
   );
   gpc1343_5 gpc10980 (
      {stage6_52[6], stage6_52[7], 1'b0},
      {stage6_53[0], stage6_53[1], stage6_53[2], stage6_53[3]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc15_3 gpc10981 (
      {stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4], stage6_55[5]},
      {stage6_56[0]},
      {stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1423_5 gpc10982 (
      {stage6_56[1], stage6_56[2], stage6_56[3]},
      {stage6_57[0], stage6_57[1]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3]},
      {stage6_59[0]},
      {stage7_60[0],stage7_59[0],stage7_58[0],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc10983 (
      {stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5], stage6_57[6]},
      {stage6_58[4], stage6_58[5], stage6_58[6]},
      {stage6_59[1]},
      {stage7_60[1],stage7_59[1],stage7_58[1],stage7_57[2]}
   );
   gpc606_5 gpc10984 (
      {stage6_59[2], stage6_59[3], stage6_59[4], 1'b0, 1'b0, 1'b0},
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4], stage6_61[5]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[2],stage7_59[2]}
   );
   gpc606_5 gpc10985 (
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3], stage6_60[4], stage6_60[5]},
      {stage6_62[0], stage6_62[1], stage6_62[2], stage6_62[3], stage6_62[4], 1'b0},
      {stage7_64[0],stage7_63[1],stage7_62[1],stage7_61[1],stage7_60[3]}
   );
   gpc3_2 gpc10986 (
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage7_65[0],stage7_64[1]}
   );
   gpc3_2 gpc10987 (
      {stage6_64[3], stage6_64[4], stage6_64[5]},
      {stage7_65[1],stage7_64[2]}
   );
   gpc1163_5 gpc10988 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[0]}
   );
   gpc117_4 gpc10989 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc1_1 gpc10990 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc10991 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc10992 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc10993 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc10994 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc10995 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc10996 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc10997 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc10998 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc10999 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc11000 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc11001 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc11002 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc11003 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc11004 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc11005 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc11006 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc11007 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc11008 (
      {stage6_5[6]},
      {stage7_5[4]}
   );
   gpc1_1 gpc11009 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc11010 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc11011 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc11012 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc11013 (
      {stage6_7[5]},
      {stage7_7[6]}
   );
   gpc1_1 gpc11014 (
      {stage6_9[5]},
      {stage7_9[2]}
   );
   gpc1_1 gpc11015 (
      {stage6_9[6]},
      {stage7_9[3]}
   );
   gpc1_1 gpc11016 (
      {stage6_9[7]},
      {stage7_9[4]}
   );
   gpc1_1 gpc11017 (
      {stage6_10[4]},
      {stage7_10[3]}
   );
   gpc1_1 gpc11018 (
      {stage6_11[5]},
      {stage7_11[3]}
   );
   gpc1_1 gpc11019 (
      {stage6_13[0]},
      {stage7_13[2]}
   );
   gpc1_1 gpc11020 (
      {stage6_13[1]},
      {stage7_13[3]}
   );
   gpc1_1 gpc11021 (
      {stage6_13[2]},
      {stage7_13[4]}
   );
   gpc1_1 gpc11022 (
      {stage6_13[3]},
      {stage7_13[5]}
   );
   gpc1_1 gpc11023 (
      {stage6_13[4]},
      {stage7_13[6]}
   );
   gpc1_1 gpc11024 (
      {stage6_14[7]},
      {stage7_14[2]}
   );
   gpc1_1 gpc11025 (
      {stage6_16[1]},
      {stage7_16[2]}
   );
   gpc1_1 gpc11026 (
      {stage6_16[2]},
      {stage7_16[3]}
   );
   gpc1_1 gpc11027 (
      {stage6_16[3]},
      {stage7_16[4]}
   );
   gpc1_1 gpc11028 (
      {stage6_16[4]},
      {stage7_16[5]}
   );
   gpc1_1 gpc11029 (
      {stage6_16[5]},
      {stage7_16[6]}
   );
   gpc1_1 gpc11030 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc11031 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc11032 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc11033 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc11034 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc11035 (
      {stage6_23[2]},
      {stage7_23[2]}
   );
   gpc1_1 gpc11036 (
      {stage6_23[3]},
      {stage7_23[3]}
   );
   gpc1_1 gpc11037 (
      {stage6_23[4]},
      {stage7_23[4]}
   );
   gpc1_1 gpc11038 (
      {stage6_23[5]},
      {stage7_23[5]}
   );
   gpc1_1 gpc11039 (
      {stage6_23[6]},
      {stage7_23[6]}
   );
   gpc1_1 gpc11040 (
      {stage6_25[7]},
      {stage7_25[4]}
   );
   gpc1_1 gpc11041 (
      {stage6_25[8]},
      {stage7_25[5]}
   );
   gpc1_1 gpc11042 (
      {stage6_26[0]},
      {stage7_26[2]}
   );
   gpc1_1 gpc11043 (
      {stage6_26[1]},
      {stage7_26[3]}
   );
   gpc1_1 gpc11044 (
      {stage6_26[2]},
      {stage7_26[4]}
   );
   gpc1_1 gpc11045 (
      {stage6_26[3]},
      {stage7_26[5]}
   );
   gpc1_1 gpc11046 (
      {stage6_26[4]},
      {stage7_26[6]}
   );
   gpc1_1 gpc11047 (
      {stage6_30[6]},
      {stage7_30[2]}
   );
   gpc1_1 gpc11048 (
      {stage6_30[7]},
      {stage7_30[3]}
   );
   gpc1_1 gpc11049 (
      {stage6_34[2]},
      {stage7_34[2]}
   );
   gpc1_1 gpc11050 (
      {stage6_34[3]},
      {stage7_34[3]}
   );
   gpc1_1 gpc11051 (
      {stage6_34[4]},
      {stage7_34[4]}
   );
   gpc1_1 gpc11052 (
      {stage6_34[5]},
      {stage7_34[5]}
   );
   gpc1_1 gpc11053 (
      {stage6_35[0]},
      {stage7_35[2]}
   );
   gpc1_1 gpc11054 (
      {stage6_35[1]},
      {stage7_35[3]}
   );
   gpc1_1 gpc11055 (
      {stage6_35[2]},
      {stage7_35[4]}
   );
   gpc1_1 gpc11056 (
      {stage6_35[3]},
      {stage7_35[5]}
   );
   gpc1_1 gpc11057 (
      {stage6_35[4]},
      {stage7_35[6]}
   );
   gpc1_1 gpc11058 (
      {stage6_36[7]},
      {stage7_36[1]}
   );
   gpc1_1 gpc11059 (
      {stage6_41[8]},
      {stage7_41[3]}
   );
   gpc1_1 gpc11060 (
      {stage6_41[9]},
      {stage7_41[4]}
   );
   gpc1_1 gpc11061 (
      {stage6_41[10]},
      {stage7_41[5]}
   );
   gpc1_1 gpc11062 (
      {stage6_45[2]},
      {stage7_45[2]}
   );
   gpc1_1 gpc11063 (
      {stage6_45[3]},
      {stage7_45[3]}
   );
   gpc1_1 gpc11064 (
      {stage6_45[4]},
      {stage7_45[4]}
   );
   gpc1_1 gpc11065 (
      {stage6_45[5]},
      {stage7_45[5]}
   );
   gpc1_1 gpc11066 (
      {stage6_45[6]},
      {stage7_45[6]}
   );
   gpc1_1 gpc11067 (
      {stage6_46[2]},
      {stage7_46[2]}
   );
   gpc1_1 gpc11068 (
      {stage6_46[3]},
      {stage7_46[3]}
   );
   gpc1_1 gpc11069 (
      {stage6_46[4]},
      {stage7_46[4]}
   );
   gpc1_1 gpc11070 (
      {stage6_46[5]},
      {stage7_46[5]}
   );
   gpc1_1 gpc11071 (
      {stage6_46[6]},
      {stage7_46[6]}
   );
   gpc1_1 gpc11072 (
      {stage6_49[6]},
      {stage7_49[2]}
   );
   gpc1_1 gpc11073 (
      {stage6_49[7]},
      {stage7_49[3]}
   );
   gpc1_1 gpc11074 (
      {stage6_49[8]},
      {stage7_49[4]}
   );
   gpc1_1 gpc11075 (
      {stage6_49[9]},
      {stage7_49[5]}
   );
   gpc1_1 gpc11076 (
      {stage6_51[1]},
      {stage7_51[2]}
   );
   gpc1_1 gpc11077 (
      {stage6_51[2]},
      {stage7_51[3]}
   );
   gpc1_1 gpc11078 (
      {stage6_51[3]},
      {stage7_51[4]}
   );
   gpc1_1 gpc11079 (
      {stage6_51[4]},
      {stage7_51[5]}
   );
   gpc1_1 gpc11080 (
      {stage6_54[3]},
      {stage7_54[2]}
   );
   gpc1_1 gpc11081 (
      {stage6_54[4]},
      {stage7_54[3]}
   );
   gpc1_1 gpc11082 (
      {stage6_54[5]},
      {stage7_54[4]}
   );
   gpc1_1 gpc11083 (
      {stage6_56[4]},
      {stage7_56[3]}
   );
   gpc1_1 gpc11084 (
      {stage6_56[5]},
      {stage7_56[4]}
   );
   gpc1_1 gpc11085 (
      {stage6_56[6]},
      {stage7_56[5]}
   );
   gpc1_1 gpc11086 (
      {stage6_60[6]},
      {stage7_60[4]}
   );
   gpc1_1 gpc11087 (
      {stage6_63[0]},
      {stage7_63[2]}
   );
   gpc1_1 gpc11088 (
      {stage6_63[1]},
      {stage7_63[3]}
   );
   gpc1_1 gpc11089 (
      {stage6_63[2]},
      {stage7_63[4]}
   );
   gpc1_1 gpc11090 (
      {stage6_65[0]},
      {stage7_65[2]}
   );
   gpc1_1 gpc11091 (
      {stage6_65[1]},
      {stage7_65[3]}
   );
   gpc1_1 gpc11092 (
      {stage6_65[2]},
      {stage7_65[4]}
   );
   gpc1_1 gpc11093 (
      {stage6_65[3]},
      {stage7_65[5]}
   );
   gpc1_1 gpc11094 (
      {stage6_65[4]},
      {stage7_65[6]}
   );
   gpc1_1 gpc11095 (
      {stage6_65[5]},
      {stage7_65[7]}
   );
   gpc1_1 gpc11096 (
      {stage6_65[6]},
      {stage7_65[8]}
   );
   gpc1_1 gpc11097 (
      {stage6_65[7]},
      {stage7_65[9]}
   );
   gpc1_1 gpc11098 (
      {stage6_65[8]},
      {stage7_65[10]}
   );
   gpc1_1 gpc11099 (
      {stage6_65[9]},
      {stage7_65[11]}
   );
   gpc1_1 gpc11100 (
      {stage6_68[8]},
      {stage7_68[2]}
   );
   gpc1_1 gpc11101 (
      {stage6_68[9]},
      {stage7_68[3]}
   );
   gpc1_1 gpc11102 (
      {stage6_69[2]},
      {stage7_69[2]}
   );
   gpc1_1 gpc11103 (
      {stage6_70[1]},
      {stage7_70[2]}
   );
   gpc1_1 gpc11104 (
      {stage6_71[0]},
      {stage7_71[1]}
   );
   gpc1_1 gpc11105 (
      {stage6_71[1]},
      {stage7_71[2]}
   );
   gpc615_5 gpc11106 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], 1'b0, 1'b0, 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1415_5 gpc11107 (
      {stage7_3[0], stage7_3[1], stage7_3[2], stage7_3[3], 1'b0},
      {stage7_4[0]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc7_3 gpc11108 (
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5], stage7_7[6]},
      {stage8_9[0],stage8_8[0],stage8_7[1]}
   );
   gpc1415_5 gpc11109 (
      {stage7_9[0], stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4]},
      {stage7_10[0]},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc3_2 gpc11110 (
      {stage7_10[1], stage7_10[2], stage7_10[3]},
      {stage8_11[1],stage8_10[1]}
   );
   gpc7_3 gpc11111 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], stage7_13[6]},
      {stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc623_5 gpc11112 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[0], stage7_15[1]},
      {stage7_16[0], stage7_16[1], stage7_16[2], stage7_16[3], stage7_16[4], stage7_16[5]},
      {stage8_18[0],stage8_17[0],stage8_16[0],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc11113 (
      {stage7_17[0], stage7_17[1], stage7_17[2]},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc2223_5 gpc11114 (
      {stage7_21[0], stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1]},
      {stage7_23[0], stage7_23[1]},
      {stage7_24[0], stage7_24[1]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1]}
   );
   gpc615_5 gpc11115 (
      {stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[2]},
      {stage7_25[0], stage7_25[1], stage7_25[2], stage7_25[3], stage7_25[4], stage7_25[5]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc117_4 gpc11116 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], stage7_26[6]},
      {stage7_27[0]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[0],stage8_27[1],stage8_26[1]}
   );
   gpc15_3 gpc11117 (
      {stage7_29[0], stage7_29[1], stage7_29[2], 1'b0, 1'b0},
      {stage7_30[0]},
      {stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc2223_5 gpc11118 (
      {stage7_30[1], stage7_30[2], stage7_30[3]},
      {stage7_31[0], stage7_31[1]},
      {stage7_32[0], stage7_32[1]},
      {stage7_33[0], stage7_33[1]},
      {stage8_34[0],stage8_33[0],stage8_32[0],stage8_31[1],stage8_30[1]}
   );
   gpc207_4 gpc11119 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc207_4 gpc11120 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], stage7_35[6]},
      {stage7_37[0], stage7_37[1]},
      {stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc3_2 gpc11121 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage8_39[0],stage8_38[1]}
   );
   gpc2116_5 gpc11122 (
      {stage7_39[0], stage7_39[1], stage7_39[2], stage7_39[3], 1'b0, 1'b0},
      {stage7_40[0]},
      {stage7_41[0]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[0],stage8_39[1]}
   );
   gpc1415_5 gpc11123 (
      {stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4], stage7_41[5]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc207_4 gpc11124 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4], stage7_45[5], stage7_45[6]},
      {stage7_47[0], stage7_47[1]},
      {stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc11125 (
      {stage7_46[0], stage7_46[1], stage7_46[2], stage7_46[3], stage7_46[4], stage7_46[5], stage7_46[6]},
      {stage7_48[0], stage7_48[1]},
      {stage8_49[0],stage8_48[1],stage8_47[1],stage8_46[1]}
   );
   gpc207_4 gpc11126 (
      {stage7_49[0], stage7_49[1], stage7_49[2], stage7_49[3], stage7_49[4], stage7_49[5], 1'b0},
      {stage7_51[0], stage7_51[1]},
      {stage8_52[0],stage8_51[0],stage8_50[0],stage8_49[1]}
   );
   gpc1343_5 gpc11127 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage7_51[2], stage7_51[3], stage7_51[4], stage7_51[5]},
      {stage7_52[0], stage7_52[1], 1'b0},
      {stage7_53[0]},
      {stage8_54[0],stage8_53[0],stage8_52[1],stage8_51[1],stage8_50[1]}
   );
   gpc1415_5 gpc11128 (
      {stage7_54[0], stage7_54[1], stage7_54[2], stage7_54[3], stage7_54[4]},
      {stage7_55[0]},
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3]},
      {stage7_57[0]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[0],stage8_54[1]}
   );
   gpc2223_5 gpc11129 (
      {stage7_56[4], stage7_56[5], 1'b0},
      {stage7_57[1], stage7_57[2]},
      {stage7_58[0], stage7_58[1]},
      {stage7_59[0], stage7_59[1]},
      {stage8_60[0],stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc215_4 gpc11130 (
      {stage7_60[0], stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4]},
      {stage7_61[0]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[0],stage8_61[0],stage8_60[1]}
   );
   gpc606_5 gpc11131 (
      {stage7_63[0], stage7_63[1], stage7_63[2], stage7_63[3], stage7_63[4], 1'b0},
      {stage7_65[0], stage7_65[1], stage7_65[2], stage7_65[3], stage7_65[4], stage7_65[5]},
      {stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[0],stage8_63[1]}
   );
   gpc1163_5 gpc11132 (
      {stage7_64[0], stage7_64[1], stage7_64[2]},
      {stage7_65[6], stage7_65[7], stage7_65[8], stage7_65[9], stage7_65[10], stage7_65[11]},
      {stage7_66[0]},
      {stage7_67[0]},
      {stage8_68[0],stage8_67[1],stage8_66[1],stage8_65[1],stage8_64[1]}
   );
   gpc606_5 gpc11133 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], 1'b0, 1'b0},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc11134 (
      {stage7_69[0], stage7_69[1], stage7_69[2], 1'b0, 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], stage7_71[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc11135 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc11136 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc11137 (
      {stage7_5[4]},
      {stage8_5[1]}
   );
   gpc1_1 gpc11138 (
      {stage7_6[1]},
      {stage8_6[1]}
   );
   gpc1_1 gpc11139 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc11140 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc11141 (
      {stage7_16[6]},
      {stage8_16[1]}
   );
   gpc1_1 gpc11142 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc11143 (
      {stage7_20[0]},
      {stage8_20[1]}
   );
   gpc1_1 gpc11144 (
      {stage7_22[2]},
      {stage8_22[1]}
   );
   gpc1_1 gpc11145 (
      {stage7_28[1]},
      {stage8_28[1]}
   );
   gpc1_1 gpc11146 (
      {stage7_32[2]},
      {stage8_32[1]}
   );
   gpc1_1 gpc11147 (
      {stage7_33[2]},
      {stage8_33[1]}
   );
   gpc1_1 gpc11148 (
      {stage7_40[1]},
      {stage8_40[1]}
   );
   gpc1_1 gpc11149 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc11150 (
      {stage7_53[1]},
      {stage8_53[1]}
   );
   gpc1_1 gpc11151 (
      {stage7_55[1]},
      {stage8_55[1]}
   );
   gpc1_1 gpc11152 (
      {stage7_59[2]},
      {stage8_59[1]}
   );
   gpc1_1 gpc11153 (
      {stage7_61[1]},
      {stage8_61[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor_CLA512_64 compressor_CLA512_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485] + src32[486] + src32[487] + src32[488] + src32[489] + src32[490] + src32[491] + src32[492] + src32[493] + src32[494] + src32[495] + src32[496] + src32[497] + src32[498] + src32[499] + src32[500] + src32[501] + src32[502] + src32[503] + src32[504] + src32[505] + src32[506] + src32[507] + src32[508] + src32[509] + src32[510] + src32[511])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485] + src33[486] + src33[487] + src33[488] + src33[489] + src33[490] + src33[491] + src33[492] + src33[493] + src33[494] + src33[495] + src33[496] + src33[497] + src33[498] + src33[499] + src33[500] + src33[501] + src33[502] + src33[503] + src33[504] + src33[505] + src33[506] + src33[507] + src33[508] + src33[509] + src33[510] + src33[511])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485] + src34[486] + src34[487] + src34[488] + src34[489] + src34[490] + src34[491] + src34[492] + src34[493] + src34[494] + src34[495] + src34[496] + src34[497] + src34[498] + src34[499] + src34[500] + src34[501] + src34[502] + src34[503] + src34[504] + src34[505] + src34[506] + src34[507] + src34[508] + src34[509] + src34[510] + src34[511])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485] + src35[486] + src35[487] + src35[488] + src35[489] + src35[490] + src35[491] + src35[492] + src35[493] + src35[494] + src35[495] + src35[496] + src35[497] + src35[498] + src35[499] + src35[500] + src35[501] + src35[502] + src35[503] + src35[504] + src35[505] + src35[506] + src35[507] + src35[508] + src35[509] + src35[510] + src35[511])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485] + src36[486] + src36[487] + src36[488] + src36[489] + src36[490] + src36[491] + src36[492] + src36[493] + src36[494] + src36[495] + src36[496] + src36[497] + src36[498] + src36[499] + src36[500] + src36[501] + src36[502] + src36[503] + src36[504] + src36[505] + src36[506] + src36[507] + src36[508] + src36[509] + src36[510] + src36[511])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485] + src37[486] + src37[487] + src37[488] + src37[489] + src37[490] + src37[491] + src37[492] + src37[493] + src37[494] + src37[495] + src37[496] + src37[497] + src37[498] + src37[499] + src37[500] + src37[501] + src37[502] + src37[503] + src37[504] + src37[505] + src37[506] + src37[507] + src37[508] + src37[509] + src37[510] + src37[511])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485] + src38[486] + src38[487] + src38[488] + src38[489] + src38[490] + src38[491] + src38[492] + src38[493] + src38[494] + src38[495] + src38[496] + src38[497] + src38[498] + src38[499] + src38[500] + src38[501] + src38[502] + src38[503] + src38[504] + src38[505] + src38[506] + src38[507] + src38[508] + src38[509] + src38[510] + src38[511])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485] + src39[486] + src39[487] + src39[488] + src39[489] + src39[490] + src39[491] + src39[492] + src39[493] + src39[494] + src39[495] + src39[496] + src39[497] + src39[498] + src39[499] + src39[500] + src39[501] + src39[502] + src39[503] + src39[504] + src39[505] + src39[506] + src39[507] + src39[508] + src39[509] + src39[510] + src39[511])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485] + src40[486] + src40[487] + src40[488] + src40[489] + src40[490] + src40[491] + src40[492] + src40[493] + src40[494] + src40[495] + src40[496] + src40[497] + src40[498] + src40[499] + src40[500] + src40[501] + src40[502] + src40[503] + src40[504] + src40[505] + src40[506] + src40[507] + src40[508] + src40[509] + src40[510] + src40[511])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485] + src41[486] + src41[487] + src41[488] + src41[489] + src41[490] + src41[491] + src41[492] + src41[493] + src41[494] + src41[495] + src41[496] + src41[497] + src41[498] + src41[499] + src41[500] + src41[501] + src41[502] + src41[503] + src41[504] + src41[505] + src41[506] + src41[507] + src41[508] + src41[509] + src41[510] + src41[511])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485] + src42[486] + src42[487] + src42[488] + src42[489] + src42[490] + src42[491] + src42[492] + src42[493] + src42[494] + src42[495] + src42[496] + src42[497] + src42[498] + src42[499] + src42[500] + src42[501] + src42[502] + src42[503] + src42[504] + src42[505] + src42[506] + src42[507] + src42[508] + src42[509] + src42[510] + src42[511])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485] + src43[486] + src43[487] + src43[488] + src43[489] + src43[490] + src43[491] + src43[492] + src43[493] + src43[494] + src43[495] + src43[496] + src43[497] + src43[498] + src43[499] + src43[500] + src43[501] + src43[502] + src43[503] + src43[504] + src43[505] + src43[506] + src43[507] + src43[508] + src43[509] + src43[510] + src43[511])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485] + src44[486] + src44[487] + src44[488] + src44[489] + src44[490] + src44[491] + src44[492] + src44[493] + src44[494] + src44[495] + src44[496] + src44[497] + src44[498] + src44[499] + src44[500] + src44[501] + src44[502] + src44[503] + src44[504] + src44[505] + src44[506] + src44[507] + src44[508] + src44[509] + src44[510] + src44[511])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485] + src45[486] + src45[487] + src45[488] + src45[489] + src45[490] + src45[491] + src45[492] + src45[493] + src45[494] + src45[495] + src45[496] + src45[497] + src45[498] + src45[499] + src45[500] + src45[501] + src45[502] + src45[503] + src45[504] + src45[505] + src45[506] + src45[507] + src45[508] + src45[509] + src45[510] + src45[511])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485] + src46[486] + src46[487] + src46[488] + src46[489] + src46[490] + src46[491] + src46[492] + src46[493] + src46[494] + src46[495] + src46[496] + src46[497] + src46[498] + src46[499] + src46[500] + src46[501] + src46[502] + src46[503] + src46[504] + src46[505] + src46[506] + src46[507] + src46[508] + src46[509] + src46[510] + src46[511])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485] + src47[486] + src47[487] + src47[488] + src47[489] + src47[490] + src47[491] + src47[492] + src47[493] + src47[494] + src47[495] + src47[496] + src47[497] + src47[498] + src47[499] + src47[500] + src47[501] + src47[502] + src47[503] + src47[504] + src47[505] + src47[506] + src47[507] + src47[508] + src47[509] + src47[510] + src47[511])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485] + src48[486] + src48[487] + src48[488] + src48[489] + src48[490] + src48[491] + src48[492] + src48[493] + src48[494] + src48[495] + src48[496] + src48[497] + src48[498] + src48[499] + src48[500] + src48[501] + src48[502] + src48[503] + src48[504] + src48[505] + src48[506] + src48[507] + src48[508] + src48[509] + src48[510] + src48[511])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485] + src49[486] + src49[487] + src49[488] + src49[489] + src49[490] + src49[491] + src49[492] + src49[493] + src49[494] + src49[495] + src49[496] + src49[497] + src49[498] + src49[499] + src49[500] + src49[501] + src49[502] + src49[503] + src49[504] + src49[505] + src49[506] + src49[507] + src49[508] + src49[509] + src49[510] + src49[511])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485] + src50[486] + src50[487] + src50[488] + src50[489] + src50[490] + src50[491] + src50[492] + src50[493] + src50[494] + src50[495] + src50[496] + src50[497] + src50[498] + src50[499] + src50[500] + src50[501] + src50[502] + src50[503] + src50[504] + src50[505] + src50[506] + src50[507] + src50[508] + src50[509] + src50[510] + src50[511])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485] + src51[486] + src51[487] + src51[488] + src51[489] + src51[490] + src51[491] + src51[492] + src51[493] + src51[494] + src51[495] + src51[496] + src51[497] + src51[498] + src51[499] + src51[500] + src51[501] + src51[502] + src51[503] + src51[504] + src51[505] + src51[506] + src51[507] + src51[508] + src51[509] + src51[510] + src51[511])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485] + src52[486] + src52[487] + src52[488] + src52[489] + src52[490] + src52[491] + src52[492] + src52[493] + src52[494] + src52[495] + src52[496] + src52[497] + src52[498] + src52[499] + src52[500] + src52[501] + src52[502] + src52[503] + src52[504] + src52[505] + src52[506] + src52[507] + src52[508] + src52[509] + src52[510] + src52[511])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485] + src53[486] + src53[487] + src53[488] + src53[489] + src53[490] + src53[491] + src53[492] + src53[493] + src53[494] + src53[495] + src53[496] + src53[497] + src53[498] + src53[499] + src53[500] + src53[501] + src53[502] + src53[503] + src53[504] + src53[505] + src53[506] + src53[507] + src53[508] + src53[509] + src53[510] + src53[511])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485] + src54[486] + src54[487] + src54[488] + src54[489] + src54[490] + src54[491] + src54[492] + src54[493] + src54[494] + src54[495] + src54[496] + src54[497] + src54[498] + src54[499] + src54[500] + src54[501] + src54[502] + src54[503] + src54[504] + src54[505] + src54[506] + src54[507] + src54[508] + src54[509] + src54[510] + src54[511])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485] + src55[486] + src55[487] + src55[488] + src55[489] + src55[490] + src55[491] + src55[492] + src55[493] + src55[494] + src55[495] + src55[496] + src55[497] + src55[498] + src55[499] + src55[500] + src55[501] + src55[502] + src55[503] + src55[504] + src55[505] + src55[506] + src55[507] + src55[508] + src55[509] + src55[510] + src55[511])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485] + src56[486] + src56[487] + src56[488] + src56[489] + src56[490] + src56[491] + src56[492] + src56[493] + src56[494] + src56[495] + src56[496] + src56[497] + src56[498] + src56[499] + src56[500] + src56[501] + src56[502] + src56[503] + src56[504] + src56[505] + src56[506] + src56[507] + src56[508] + src56[509] + src56[510] + src56[511])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485] + src57[486] + src57[487] + src57[488] + src57[489] + src57[490] + src57[491] + src57[492] + src57[493] + src57[494] + src57[495] + src57[496] + src57[497] + src57[498] + src57[499] + src57[500] + src57[501] + src57[502] + src57[503] + src57[504] + src57[505] + src57[506] + src57[507] + src57[508] + src57[509] + src57[510] + src57[511])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485] + src58[486] + src58[487] + src58[488] + src58[489] + src58[490] + src58[491] + src58[492] + src58[493] + src58[494] + src58[495] + src58[496] + src58[497] + src58[498] + src58[499] + src58[500] + src58[501] + src58[502] + src58[503] + src58[504] + src58[505] + src58[506] + src58[507] + src58[508] + src58[509] + src58[510] + src58[511])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485] + src59[486] + src59[487] + src59[488] + src59[489] + src59[490] + src59[491] + src59[492] + src59[493] + src59[494] + src59[495] + src59[496] + src59[497] + src59[498] + src59[499] + src59[500] + src59[501] + src59[502] + src59[503] + src59[504] + src59[505] + src59[506] + src59[507] + src59[508] + src59[509] + src59[510] + src59[511])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485] + src60[486] + src60[487] + src60[488] + src60[489] + src60[490] + src60[491] + src60[492] + src60[493] + src60[494] + src60[495] + src60[496] + src60[497] + src60[498] + src60[499] + src60[500] + src60[501] + src60[502] + src60[503] + src60[504] + src60[505] + src60[506] + src60[507] + src60[508] + src60[509] + src60[510] + src60[511])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485] + src61[486] + src61[487] + src61[488] + src61[489] + src61[490] + src61[491] + src61[492] + src61[493] + src61[494] + src61[495] + src61[496] + src61[497] + src61[498] + src61[499] + src61[500] + src61[501] + src61[502] + src61[503] + src61[504] + src61[505] + src61[506] + src61[507] + src61[508] + src61[509] + src61[510] + src61[511])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485] + src62[486] + src62[487] + src62[488] + src62[489] + src62[490] + src62[491] + src62[492] + src62[493] + src62[494] + src62[495] + src62[496] + src62[497] + src62[498] + src62[499] + src62[500] + src62[501] + src62[502] + src62[503] + src62[504] + src62[505] + src62[506] + src62[507] + src62[508] + src62[509] + src62[510] + src62[511])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485] + src63[486] + src63[487] + src63[488] + src63[489] + src63[490] + src63[491] + src63[492] + src63[493] + src63[494] + src63[495] + src63[496] + src63[497] + src63[498] + src63[499] + src63[500] + src63[501] + src63[502] + src63[503] + src63[504] + src63[505] + src63[506] + src63[507] + src63[508] + src63[509] + src63[510] + src63[511])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h58fe0c67938d5a7747c9753bc288794fca6ddfebab9bfd379e7c35f7ae0892faf0ed4c74a8ed23ad541cbe3f89b989327fedef72bde04d97cfecbd82012125379c0eb4b786f07fca081261d886ce01d8c77296825cceecc54922f41fa2d8db9162347516f293d4f5215eae34d779f0c8872dfdf9295e9fa58dedef52f18e93743d15bf949a52b77ff391c43127d8b5856a3ae2595328fbb53b932747cbe536ba1d256a226433108b4e117516e54ef6aaae46fa5921bcb20abb76ee63b60f3fb57ee2ab5853a33301fd09fbf206183df782a3e5c687363a849b5fe2ddbde25b0fe162706aae529280b806481c92ed994a6dcbe0ee771af04917537297226f2b71c82c506e763992a03c63a8d2d912394def5a74735a1c36fd8d6c8de2fa330d176dcd0efaffcb8613e0163af99f8ebc31fcf2f2dca8deab6239d9cc9865a99465e18ea78aa2ae968047ec7f5bcc789b733de6b2482dd57be95232ed774621fbf4c6ba95d549cbfca59bdf62abcef805ca7bbcd6f48f006b56e88f35313017318c0c340dbe6614d66fb786725244f947c93b23c52b5ce74c24f3feaf9044b4813cede8b96b77854245fc205750c8f65d7b21b415c491e7381613030b6ced4f72c04762604c5bc8cab39f39388808aa08685a790bdc4f94bbf278524e4b7fdc5babeef5cdfaa7f907d24398af514b254b4972d94d8da1302389342e5da79eadd0b24151ef8b7d410c7435dba71a86378f2b7f87434e44f1819960c21b79dbf399c999ef9eff3a1ed34a97f39c71d4b299740cdb54078a4236374c7422e6e2ebea1844f921e7aef6cbe0cd8bff4f1324fc7df6a3a900af0c15d1148008443d98f5c672849225dce459b1c67884ec8eb9929d26d988ec55b07be3f234c04d729307985dfd719b47f854aec2b22fb5a068e009f7176b7c7e87a84c3c68e0f34d158e7f7d5ec4f650741c1e3398309365b2481f96210004508328e4a89d845dd1c7768fe2b5fe73a471ccd9f608921d8e637dfad5b20caaabd68a2f859f2e231b7c65e2ba6ee142a9c70a5a0347f87422430a82aa930afc9e53b9f3d243584b4317924859e72ff07934cdc2da1e145d5cb9bf193202380b0d5c8d8198d093aed996c0136f8aa2e0f36271b50d5d06ff63718aaec1edbed55cad290174ec045941de9b8359d5513189d9b4e57eadb8d927eaac74c32d143491f7f3bbd5a0691db39e4b71385abaf3efa3a5ff007c1c49718fa9929c1d5d30b5427b5e798aaa47fc1c0bbba0de02946bbc7ee9716fde8bdcaa173b3c2315857e68c87d701abdff0c6856d791c85ce7b8fc3d580b82622a5153c4f96319849b4377fd5d0c5d5db89e8092d4b982ad09c1a2633b0976d21dba5e7061544f5fbe4aa3b90e4c4045fb28654fa2c76d324689304ee5834a94a4c81cb3b9d3382361511ec2f4d4762ebf5a6969618389dadbb1dd3f7a92316aac16e496e3c9c8dd214bd0cb27e0471794270e458fedf54a934f704c9ed5df543106bea0a3cd270745cd12d4249de9942d185991e14976f8adc283d2bdc3a158fada28b8c8ea527f42f2312dcf06e4e577319cabf8cd11f1f29c89ea3040b82a64147ab357337f388e69f382a7cb5ba412f65b943aafa7c8f8a5ffc869a9bc425f65a7801a938af40c2561aafcda845844a051404499276717d9184265091e6bfe4091720c72967e1f759ad3bc810c9349889c033971054308ae10d1494467c3c169fd9eb844b4753301dc006454a34ee22258cbd0dcb2b8e43ab2312775c70fd283d1a7c69a23a193a83753a6be632f6c740d388941f8703ffc2f682630c8123b9c8e7f55a5be0d83226b078cd134693f262b49b49dedd16618b33f04850785d388216d832885ab8e17d49232b23722e3237f00530218ca39e336c3df29ca4ec4a1936f010a5de433f1b02d1cfe85bcfe7c0eac89811731a94487dfee71f4c593d0aec26984bb042429412e1442a9004dc6eda221e08d2f8f1a5559ce8068e12c84dd4538d25d71fb8e3d19bfd8c6b56b07d77a555cebdae8bf06f630aa1c516186618bb682b8c37529a178f0556834ae04bbc39582d978871dc052556a41d582454881c80cfd2e2faa0b9ef7589329429ec6fb9cc05b58ec1c7b7b206e8a2e213f20b59e1b836873ff56f89bce561a41b0f92ff200be6ace59610f5d00c873f4eeaa52a5c177e662bebb38c0ca6e71f25103c8b59f61fedab73d4efd6fbc64ad499ecf60de4196d74aad892af02400fe02d92405d2814de261e4ebb37348a8c40acd16fcafde231721321e7537b52ce569c1758ed2e1578f2bb16466d723fa365315c2f4e5d4ae1b27db91e1645711968ada168a32e4555ab240370485abc097015b90a8deca34039b50ca02af9d2576001661972514f93fd243920cdd681ddbbc66b78c00600ce671524cc1edefb6cfd1eb7663262cfcfd7379c5d8fac748d8bf8c353318da04dc967fc49f48314196a06819ee1ca131a30f7abf6897aabc5211f5353955b69c4b326a3f93f1a4a508a8dcb8689f9452f6523d6d7fddd5fa89774677fded6660ae53752544fdf9edc38ba8f8e480f14f958b524a8f9e4daee1a66821b5bef798c4b7e8e7a06ffd0a0239bbe50c3d31cd0997fc7dce16ae80a36de416d790fcd90d70f20065e2ee32fea357da43b0aa3581662a56a6d3fcf02d183d0d582b65afd2437b57162fd4123688e08c07e06ba02c2ad01a1e50df2a8a71bcd7ad183041ad4d4f7ba0554ceb5c80e9ffd0188cb96559dd73d073ba025cb438a40ea211cc2ff0133a937801ac2a83406fbe697a21cb28871f9b34d0d90715c1ee0769afb3b1c5d8d9975ad6aee697c1f64e3349e6c5b8e0e717be317e93e7e9223b9bd8e9bd84fb4a1d6df62f0a06d1f5acbba173c367d829220a17a9135def7ca1b21dff14bec343f5e012c8ce1c1a9dde772b53f94b3da0575fee1458530597f078f2bc69cce19c0e0ff203587c7714579ae9d00efc7e1bf379ad1961bea27dfeda6f3e0086e3ef726e40809fcb5f3a3f87631a84a8ae46678642e667a2b9af932088308646b409c26cfc87e60b2d57351d2235f145d20d3e53b5fd9e5ff9a9680c17e86a42fc6e974ee01bed9eb19418e2263b238824a71087308cd7b333ed7a48bc0f45d72d96192d2c8ed460b3693a17bd592dd711b86b6aef815259b08438d70311634615ea19216927fd5ae2e8f85adb553629000d207512542473ebdf3ab3e7fc18f973c64a8405096ca5d0ecd89e057aa3df633290bf1d0b42a0bbc07ba0b4a1d2896e1dc75cd432b42992eb4e40615813957d5a4fd7d2ff7bf36adfbdc1938ea27361006ca496182e5a5267bd8c858a3b12c04be9f9761f3267147a23d27a6082e974d7c3bfe662d4998703e8e438d81289d94c8fffcfe5bbe22fec33884b951e0d6483d39747596f6d31b1711f7966526458a70f283a9decfdab71bd419de12b0bd26807494606ceeb350bcbe349b636e328ad47854f94d82faecfbae5bc090333e8473f8ce78bc47814a3971b033460e97d760363b2bb56b54006b87993006d2c69e11716b067db0ef8c3690a63628f458e24929e3fbfe86d42e9aac9a773e42520fa8e66b22bc1c9a7eaedb1533d702b9a838061cf16e173cfb8b849b909b8452bfeb6a31714f59af55ff7b5ca4b1cb8f01f9cd5ec5b813c826220774489c666758754039d7108ddfb187b5bbb308dd007171ed37de1b20d2412ede6c87602f095d37574c0563a5bb16da36b826af64445e074ab931a2a22035cede11488eefdaf3abf5b3cc2879c1193d233eb1097a510923010c0eddc6b69cd2ba63682e105e00bc9b48b6b4bb57c49ba518fcf68533a4851538cf3898d87d493f320bbf4113a9a767b0f30e5cf35d7601685193211f905b1c9a77a2315055839adb1aa37d35078f37e0889c6464cdfd16a3577ba02f8d9e1d18fdec081e703040eafa7127187acb55a0afa2c2e5f74d890b52147a371a528aba28d344e8a1c4c7bbbb0c7d3a2ab1bfc94f609493a9d5d4b0b6a49d0263ce730e5822a32c7c61232520ebbd4695d77cc29979891a0c8632880bd3fbc1aaf4ca2ad5db2963a08a626d630273ecefbaf99c04c760f8902d6cbbb45f8ec13df3af659b4d576f5f5e4fa0c2030bca61fc7e879e247feb1405d30ca18f8d9f37b82adc3a0cb0d60f5db810e4b2708efaf1bc157b9b01f91e57cc39604a9e9717eba70ca6dfce4a99d6872f2cd6e58307ae26197bca959fe924dc0d7b73763816058f2da9f4e330ac95d45a25807ed7255bed7beacdb42e5fcfee87a54323835092767adaa32c19b9172dfd75f4bc4522229c740ba314bd19172a1df7bedf98bf5c1513949ea5b1a86cca9e66fa9839898d3eb4464054499c910c040aba7c660ed619bea17a665a4ed5605f100b3f10fb6c9aa8801d7c6d326715b36b800b6c0cedff70351b56c82242ac8c1e7fdb4d60c90cc2f8f7a02c6affdbdec5e61b50f922a4b48495b626ea1644ff579636d5173279277214d4031a42edefb4cf4d307e58d40c6846463ae8c9bdd04ba093385666e10ae7d3fadaaf03be18397eaa40a5a66860f46b2fb8676a83ecc63a810fc21a1814896b2f86cfce65ae38c452a859e38817fcf92b8b01d1e26b85cf60d242745b03be661228d3b1fc731c278af215ba1c43acc8281cb8a1cf8a893818adca1ede98bd8d999516eee79cfcf00d005a9f644648e22ba008f17de013c9b9e47a596f313ea98fe7c76ce8b49dea30771e7f0e5c593c3ce18e8451be7bad0f6bbf78576e3afb98649c89f11b7691d1e9928b5b97c0095cd95b1e269aa436433833da43c26ee64b4c91555269a38899c028133d9ea87c966192f6af69f40bfffafcbc4a687524aa90b74cc4abecc7eb1364e6ca0f6b2da3bcfc585a7efc4e1c146405e3c1887c773bec77b84b9106ad25d69eb9baa8c03613698ffebd9c56edde74a7ab87eee93d0942cd32c820af9190a18e4e9b431c78bee7a8922ebb7835c36a1c8fe3660716312608a6f2f0519673c876d412c1486845bd6c17615d5eec4d2767c38f52aa69f0b445e7dcacbfc06c610c5fdefa1cb486f56cb1cc1a198760b44d2427f7d9f80c4024d4589afc379ad362b7ee04256258140f2c6a14ac97a73423df5c60384c3b809eabf344b46432ae9a1a861a3f8b0328ae12973c27274eb5c417f7bd82b5d8b78bcf83483738725a7d7dd4d195872555ce7e82f43c483b3eda1ebe105c35d33f5617cdda99b1ef94e087cc58bb2791756bad737ebc1a67cc493caf00a5fd3613721f709fb8f891d9c4dc6846d77bc6a88424a38962ba138ab32695e99b6a822a7b5d7a06c7f28886be1d31e3700c94744e16135daa7c5080906a5643181e2067cd72e28018f26104704ebacdd518c46d8f1e5b44df54e6a368a4b56b68d0039b94af1efb29865854d35e6d62ab052d9a66d0f7135ae4191a39bcb072d947152f39e519a02bb7c95c7c65d9d00b88ab54160df4dc48d2a1e0ad902ac96861ac580430ed70efdeb900ea3f8eb54b4711e7559694645a60fead27dfc5295597a411168917b3aa23e9c9382142f92414870a6ebb9bc78f9a31fbf8eb65c592cd3cf734e5f5fcf3763e1b672666cf2678ecf4892c7fe72ac1b4abeec8186cdab759f27e3a5338d283935ed5f9fc742a0842f02d68639ae8b68d57cafa18d2a3fd45c4ffad1152dd7e813dafc17ec6edb362d7af964eba0afae9966ef03a6a81539af84debdbbb0c105e908e6f86f4c7d7599165ec1adc329225cc2c1011f87551d6b6b9c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h474df06f7c47189981b252da08aa16a5b85e8c56d5e51128704acc6f185826d658cc294b94847cc850ce7fa0d33390ea27ab1703638c317080539be7a869e41b86ed4271eef84e661cb4ef418869a0e329e6b6c74f650a8a86b79edbecb2265123843cf22443befec170a16714c5f95891f0200698a156ee930d2c07110503186389e2556a01905a60fa7e53d30060225df570328640c2d1fc61d5ec43fbbd50faa0e820732c56ca8d483dc07e64fff77700f42a7f46ac8eeffb1ba048b192eec2ecc2095ede79a50b087e80d973fbf58cb08d7d87b95c9a3b6a05f91896953e5e00509bbaf7c8f64df02f540960c04752424f27ae4091ce62329ae94987cea638380bffa3d91e647cdea657e2aef3f5a93329468bfe6cf95aeabc2828f6caef553408f2c0c0f0279609a4023cad210737efccb3a42ffecb0930e2750db8197cfabcb402f5f65c73d3dd698648538a9a0f0b5dffe86c6fc5e0d372c448a63ac20ea7f7252bb67598f213521b1e3b0ccf6eab305a0ecd1f86f30116e466cc23ceed15eae675e6c1987912286405b53513172ad18107eef1e97ee6c52e6546b2b753b95ee4c477702f9aa65e0ec47a25a3737c859da5a551658a869739215b30e1c537a137faabaab6effe8e492b350977f4c57a2c44adddfc6f18d5fcefdf241c60eb3ad43e930dcdd68582e7281b91ccb45a111106ff83bd125110881059d51013cf1b46853ded6972afcd8c248bcabc3d4785812eb08f1a1a970960568d7dc8ada40e58200a81e55d4922cf5aeef6c48ba4d60d5f5b5462acfd4ee3dc809046284d048bb39bf9b61e963c932d3f7a15a096d21955f7f0618a8c86f92419c6f4f54f5f62061049890105fac39e0df674a75afa505353d7cac3ec30b4c931a9b468b440ef6d0119ffca79fce0ab8cdcb6663348e6de2b2d0a68ead19611cbd16c69fe5ba8072d619114ea02207fc1d453750f8736611103b3b42c3fd36ef6058780a3c17cbcc69bbaf70ad8bde8526a7ce082a7ac9c26324b9fce5da6585c48e0a1e22d645fb257a97afada105002656a88975dbfc9883864a8bca9830c41194a6b484f1c97a7d24facd223a905ad6d29fe7198771a192e615e1e1acc8585b3de0071262100548046099c37ffaee94935087046fa972248653d98821d31b48449ebe35471da3da65e6b86ec403ac63f48992b6875c24df2670daf3ad4456a9a096d2cca29b8761bc67fb1c0bab008630dca289451d086b234ebba7a0f7bf164084be263684a7701e6b93ddb2778f34f50fac43a255a9cf8c41ba9c49d6ff05cf88e7aac1ab6b2437d30b65e55769e5aafc447223a05338f55e9f327ac2699353a675dcc134173ba9e9292096a11c0d7b0e1ddcc183688f1cd530fbdef0a40d0bff67a451259a45724e978e62db366a434ada33a746d5ba904d0c5f6c98b430cdba6a39ef90799bce0bdb5268b737fd27824ff92c48fb035ed7dae39a023da956f0210501ef2016d6695ea14a93ee14dd58a092124b2dcfc774aa9099ffebcf206f437855e8b69255483fb5d1652797b499796e40ff408ee6be7249869a7ba3f8bb18eba74128435437b289a217e587785398ace62626fb8689b036a4fa3292d01835311909b4fd91af0c60bc8bfae4747fab50739e0d490991d5bd83437b287299069227e97e48b933a0c08f83cb1af8b4aff32351be68417ea3f20309d1c3410f8afc31e541360a8933a029795f4075c507444b10106e7518a7a00adc8bb7520862c015a144b01dfade6172ecf6b4f7d725fe23d541bbca80eda53df80aec8b10e0f56c61940ab557d0240fe9c719ecb77af8be5ffc8fc9a31fed769cf0ae176d1458482316144de1ff76bddb7223c6d0214400aeff7365349864525c2533ffd6eabd4deac1d4a7ba34c32ea35b8520d1ecf24805aa467ff25400509bf09e2677dfa59a23ad0366909d04fdfa3f5ba20108e91e3d976351c4b803aba3a5d62f4f45e9864de0b9273e6d6672b7b59b259d022426c25e97551f924c7332db192f0008517a19608019b86587f811dee2c811c24c9a2ed2a4ebcc60997db8f609ff8f3b50327c6598daaaec793b0d14183e451b9b3ba3187f3ef8a2ff9bfb5ce078d8916cbe8ea659bbef7d273f08ed734843993c916bcf6dad33c701c48fbfc20bad1e7948cbfafc56ec7c573811ad3e09d9c0b9b0d0e4fb531fd1cc11d6b5c7c10e77f58b0ffbe68687bf1b7b4054d3890ba8f848e2e61a68f1d6ba437fceb6f0921a1a2b0d3d2ad3a02dfafd04811d53e66388d91b683b1c86081f30df3156113e9654bce52b8ea74e2bf222a3f8fb7fe0b65c70b24420f0b9087a2eb2fdd933169181bc3cb75f346cb37e73be453e0a0ab635b9003b7f46ebd79536bdcd38ea5f4926877ec69d47476537047defab23a34307dceb8cdbc2043c7aff9f4242531f92e027b8d3f2d334482dabe2f326cd8f3f82bc5048506dffa724cdaeede1cff823aa2d143f3df1696c07465ba7d8d13e3fbc2a7717fe381d8a7b8098deb161aa5e447dd9aa8f4655c2a226a21ee7fbde420171a4442b4fe99e29cea43cae0b7ee16c8b1085d0959d4f54e7ddcc4a1d4b7cded4e3a09f3251852c318237bfa693c53ff79821458a6d96b7903c6c5cebd19c2c725f9d0810b9186262f71886a78aa7e2dae7305e526a3920d03929113034ad4229aa780b25fe93364b6b22d551bdf176e54f122990218c582a5a09aad192b1c7b887f3a9c5c9607fdf332190f1963f2624f08d3be31a1de5f92a500436d9b05e44e0d4d4ded5b65f40545b7c5e49b7b25f25d5fbf0bc4645a6a25d2389ef8f57720a1cc71fb97ce2e99c0e8b0ddb534f97f1994a9949c5c6805d90e5c9e7c06ed56753cdd2111699dd57f9b019e04ff42991a287995c18c8074c90f5d6bc7788a4074abdb90bf271a6739a288023ca2d28ee77d07c8baa58d0209e01bdf885fb9b03bf5f4b95c32e25ab5423973913efddb6f6b26a122424e14c6ec30984bbfeb5c0f2b58922c0871192f81d265e88e795ca098a65a3bba75a4321b3ba7a7a88da68e4cd17f35d2fbdcb240c4172f959a0637ebe449758db7fc38b4d93d138d42a6faffe989a6b868eae1d133e147f020131150fd539d4f3d17e822c315b3baedc9edce9703a62822455c6d0cd8b289470a6ae8f0a0e8ec239e7c7d16d32f6ee32c93a5b51549cc68752ff892d41eedfe838b1bdf5e6a8a3b9fc5507be7249d0c00e5a90a613ba92a58551a6e3c809ee067b724299c76b71c948991cdf93cab33ef6d2dd7466a8bc3ab6de75346b689db63af01631825b90daca629c595214d9fb543a1a77572747a8dca37c2586191fcbc9968adb52cf1d1600ba9dfa751879a36790217b900e05eab73b503c0eed66644574daa414f823cb56660cd40aa4fa9efcc2db5bd119306c593dab9c60bdb14bb769f5ac3f171269ce08f767de219dbf1c9de7fa6a6bc0c138844f23fe09e37aa0e8860c29758bd70ba6ba8eb29774fdbe4a24fd01a42d6d5295dbbf706ed7c11ae894308d55f60a743a91b60346868a3f12e8a008ff07e8ce873d96e456325cf678158750844e06fc2c4855b5f053cee5a8085c275199159b0d225333a2e5d7789fe89f81ccb620aef4f94635427eea44a3a36eb287ce1107658fd795000c87613baabbd3ce4639af871f8edd764cae4d6a8ff3df41d78eb356f1668c99bd237eeb8b37689570c14846d0636190f3a740b040577f14c9e3b31b02734f8888e6cf62ff32f3125217e5e8e9ca43b5973dd2b1095640318b3007008a4db7c4edb71b10cba871f0656d36892395f046a574ee3cb6fe2bb9f9295e63f0c8c42509702e74238756bc39751dfdef30fd46939af21925bbd764a92fdcfd4304f13797bc1eaafb220c8b222d5913a1f42b7dbbca0d6e3a7daa72d8d9962237ab8b1c3f4cb979049389ec25d1727ce55de37f029168bc318dacafe81a898fdff2792918672525781d69bff6a855ab297caa58d2b6ead1f6d2e3a3ffc65ea5781c333aa37470cd53cd6bcdeb1e6d2a2bb6f8563a02abfe0e3a9103a8c8860e8b8d200ab9de7b7dd8fe64558c414316d193784618289e88f8f803d9221fbff5fc09a255a332c1b1a65d4358390003632e9c9806536e9be9405ff42e7bcb6aa972d97b5948b280a0608d3142c79cd7fc5b2819871b90a1a90eb79535ef0d6db38863a41a3163aef51d05b1417f2a4094ec21aae11f7f40abe6be78617a634ee436765b84d18978412100fe26ead533717004ee08e4fdd72b5f006b6d2394c45f924fb56e3b033a8af22ee376fc005617f2ac44a41f37f85497213bc18f2c842d2297e1c246280173b34be491f2c1ad15434c214562d77aa4ad968ed62a926e5e3b06bb96aa836f6ee4be2428ed5f6982c9d1f0096ac72341e7101e5e502695e7505cabc71e27cf2b77606c059c81b8d9106ac4bb1ed21d733a61bc902986deea1b8933c600b64b0fbf124203a1392b0cbfabef06896d6e6bf3d0203afbbd0b84e084ed32b86f177171ff8eee0efa0a921f4fcc322a86237370f5255278c3f457feadca7ce524f37a1b9827ed83364e45acc3cccb2272a8510162a6c124fceb87d4cebbed3c8e964b1fb10267adaf1da4e70e6286241f1aba82c32d562c01296eb5b49dc29c728c2097494c3db88790be26144e873e335af3acdd38fc57d960cd96a9e9d66a11f8ea91a958c51fcf80fef418786708b4b4a1d2facd8b062b2fe2b53c4f5fa43e85147be523f764590954939a5c435d16ff36b320788454eab730e42eeade1db388c0b639c0eba4dc04e0ec832362587344dd25b15ed2e0342d55b8587a9707d163dd50b4ad38930ea8ae21a93e613d6fedb9fed9365e3dce1a5bbd7ed9d278074cea244d9d7747f536f7beeb52093a419512d9dce89cd05e325bb5faab565ce8e57e852e3e8da668a55c72ffb4d6b875d85e85c1e8c440ebd3cbb62e1ba641c182ee80c4158346aa7bdcd7f3ab7f2461910b5fb302c92c4cff992780a0685ce73ca5146dced0e283260007ecc04a42de2f3b6d0ad166cf1bd88f06b5dc6eebf9deb0a120224319a65c0c758386ff2ce4a11a4c94a2ce92946047b328a7f22ca30b05bc70f8fe83bd1916be02b87c1365a739188d79a7395240ee0d7e17e1f273afc691e1d37e3d6ef7e459aec8786c1f51a5a56ee10a75f6707847de60ece21a8dfbe1703da82ec42e0251bc980aeecdfec8cb4ab6b9d8152625691aaf493be1a45c66af2eaf6b048be77944eba5ceedb187f9581f13604441f3ad8af6c375b8e4238d5ebbbedb164f711db0c8d17f9ccae1d82b28b86276a84f7f49734fb9b3f4440eb92639699519727057ec934b75027acdcc9476c1328b280753c008051714563c1f89fad1aad09099f489fdae97b75505e7a2876ef8563a52d99a069300cece40e21b4abe57219d3ebc7269d73faede0fa68cc3f723f1e7997534e47f1f78f711d8fcde4d735ea035df4d311334792b2f7b21c49e4b59137380373111e2daf827e5450751e83837087eb41388c085a8eb4f4adec28d4fc50b0b87a9261c8cd7a0959307e7dcb3afb6b5129790202da43bc6eeefdecd57d2cbad7d812b9d25810eee7e5b148a3d4a53d5ad6bae94373e277b4fbb57da806088ae9cbbaadd9171a45304acca993ca77a78b42b9f4e80ada9a571ace0e38cf3bc598d07ed5fb99457b81f7b8c8d7c37a491d01faba33fe233ffca8ad3768bfb498435ea5d1396b547627de3d668331df51ffed72c035c8f085a154093e974d7303f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h328fe7209bb1f6556c7759bc23af0cdcc475d9d603564fec1e04ddddb2be9a5a84295b7d84c4281a80793305ad0232a74c2882cce0aabc81f9ad7952cb3d08f22a71675d2082aa5dc1d1ccc0a70f02eb2cf68aa0b7f3a6879d230895527305ac26ed36c8ea66833680e08f31d4ea7b1a9bd73474c0bea25bd925cdf04c59088c24a955fab867c71fdf20606e2a2a8de27a252f9bf754fb135b4bd5c7ddc8ff7474720fb80332509cbb96d120b4e0f9848b4d5b1dcfef5fc8f44554bfababd4470e10b566338ffa18c70527b6acaec8b281b79ec0e88d9857c134bfe2c51e0c68660b4e3e75f988b6b1c49d7be194e0479cc809fb1245d96a4018e25f93f71fbe7e9fbc4c45759e959b5a0e30b6e44fe2fedcae1aab22cc33f1087306a89becea25975f1162dcacee29a63994794561e3165ee733d9250e4e3a02f0fcc808c5384a178f9cc79ba303f28327e2a0ae2f19b8d655c379d468a0ffac5b78df1ba9e7df372c0ee20cdcc9912561e52d162fcd0b7b93ae609486a6e4cade39a8bd9432ea2173da933e38ec586677bfba20626c1fe5734d9741b821fbf36d0fd9bd833bde166e45461da0c2d50ed4bf90d19b737d76a4ec56454610fb80939ab80ae02a6d48a130bd750e7e3bd1c2ec5200c01557224edede5684d15a6167e758ffeb82d7e68b80b44a24d6ae1cf339098a6d46a6a0cec8d8c42e49bf7f0747c0351da1f6aa7998ed3a117fe0ad93e3278da7d5db24781d5e1ea84c35086bca3b69bdb68e48430bf2c062b516ebe01cc5ccca9e0037570fa21cbc6b4379daec06a8984d08c5287c3447bfaa91eaa3e6392a2ecaebb00c266692ebdfaeefdd89fc6107679a2dc22c8ea1c7405c79120e6f0e5dc54bf803fe7d7cb46a472c8400b443ec41d8596378505c49590089350b6ddc125a5045f4415acd3e715b52f02882812edf2ebdeeb3d820d37a43b92e78fa74ee0ff504ad30a25e37637e7eeb0eb73af2328fd4690aa8096325be5f9e7038612ae95370943568e4f5aaa2c4aec2d335b16ccb0d45e460ed17a9086d3751c7d7222d4ba55ea0b1681d8bc7354cac0328fb7933fec9464bcb148ab1b1ffdc10f4fae88faa1f0f4f6054dd324b91f316fd04fa1c37a28cfb3a97521b81b56aad783cb1c5bcb6a14b00e97c5f4b04b52877fc7cf06b9184ed5fa4bc804c5f2b3dd35a86d5b010b8b939fffe8e47f70abb1ad759b99040561a0dc44b76874b38b430292515ecdb5631b5fc16243dfea7b8a61b8bf7688eb22813dd47c1a5f9f80177e5f3c3b72665ab1ace37f4d597da361823d7a7a0b1154df5f38378eb865d92f47ba4d93ddc416e0fb056cb4f87a66a766a31c7e0f8a9037c79336ed9a56eb83b1f57077311d3a7ccf7f280d5c10f130c512961047fd08099da583e5f620c95a84223ebbb58fa85d32ed3616f57fc6c99c30d9948809b6faf104651d0b90a5b05b29f9f110a419e735a211efc41f9fc7ea7795af6bdb18dc79ad36e64952f15ac28b6de09b9df672c8c2e6b7a2d3c079c2726af2f6f33743d4dbd4f95c4f84f7a10c65a07a44065880d281d3fa9ebdc2ee74321898f17d0d7414f49f4792f7f4759177493745e94b5b13b74f3bffeacb436dd6168dbaeb153199cf1d84412b342bcadf785558204a0a389d6be165a1a90b62fb6e20e47627ac5147f1b0890f4e38760a809bf439f34dfc81a824d25ecf4c21945bbe0315f596aec9ad219cbf33a056173b3682380b03535481ba4c49ba616a9df8ed62c914b5f08b01d06579a35d9aaa644249fea3aad39f2870f02ed9faef6e73c738ee39bb91ce520607e3123af7e72a0da739f501fd3ec0d14cfd074e72106e660c8242f2e74e31249a4292ee749ea54aad64aea28798fee719ecb34a39c7e00b28a95ae2fd0e926b8915b3ddffd183e3372ced02d2de4ef654662bf0099d1f7c1453a3424cff573151f8826cf115782aaabf6ac205f8d04d88abd316e5530a3cb996bc591ad477974e8da222c9c4708abf1d3190f323dfe5aadf0784bedb3b46b6dbff25fc21582406b8cdfb4f48d3d8f450a326406148995083f8ca3f41894345566a340ee9f7a1baaa11aac7575d5e4bd0a3229ea136d8d0ce9af7f4599a2cf846ea1fc7680921f266c4d0ff84652068a6300bd03ea7d335b7299ebf0e30325150992e3db77a65bddb94d1c638441edcc656a7c6df0c0abb7e5bf69721a20794b0c84629e605111e0da7ea1a107e9e92175d864689e9618c345c9d96bbcd5eab47f0a7386c49c18ae48e85dc9577bf49029bf6623c8b38b42f3ac32b4dca4a99063c259643b6e614c9a458cb5260d59ba961e8b621ed552b1193766bb8f6b9a1e24f34b7311fd4dddade2b7c27b954ffdcc75d40d0bea4fb180e30d1676e0751ff56d7d4d9d935f5e3fcf204cf7b362adf4aca491e36b3c187855eae3967ab21426c05913b611adaa22b5a7330a0fec959cc8d511531041f037b4f3a25a903e897f8f6fead61bc1b34580f740eaaa55deff7152c4bb149fcae7ec36eecc31df20d07bdab488fab05eaaf54c4feb60fa568fc8c602464b43509f056760c41b35fe2ab045b6ad2f447e3107ea6bb5cdadd983ce806a8e16f70346a570db2a9dc7d00942a2b27f34cd7b61d79e0986ebb64102e9bf6d3cd7c252184cfbfeb7875d72b886b0788b389307e3702c9dd7f6bb99a4e184338b83e3a8c553ec1dc02effe06a0d91649623a9d780041dadbbf963157c2bd69effeb821349ebc8c294fb62ded32986b292f4f543126a4025d5a385f41dbebffe5ae80e13608880e0da0fb849e48db51494e587231095a9ef4716a9d03098a886a0b5aaffa46a1b0ca3ff962666c6161cb7b053a291d317d746f547c7e174fba55e47af33bb7adcd30fc52da6e9185f25f5be853ad014c9e4916a54c3e74a67d8c80c34592ae60d96cf095b7637422c77d8d1194bed905cec62750cf243f88f1ee404cbf36bc719702bb08164f4de19f8a5ba7419c953074085cba24e2c42350856e27c53f34d715d67471e82cf8a09bd36acf0d205adf2a564d3350f89d3697ee4870c6fafd205127f1ddfe1c5831ffcf5a0e3a6370f449169be37248339ba9d2f22bcb8b4de7167f197e4e5d2d9228eb433283db1b3a572652d33a4fe6a3b0438a4bcd7b54fa8d384a6b9d5eac8a44cd0bc875bafdfa37e90ef184148c1d8524b53e57015a9e4d10aff03f0194839feefecfbb24073a95babb9d920320c7bd2c0235024cfe075a756fd31e55bf4be27ffc01587bc0e25310f0f8361dd832558800c7188312060c27f69a087ab69fad965fabcf6b5dc1cff83b9392c6f69b52f40ee6125f65b11607ccc8abb68107eeddb4e245a33b74209fa8e72c2424fb45375c527ec8f12f4640e33ab188b550ca741cc8ab69e30747a6576d5cb08299e2d4ed289f008c608f041758616dc8945c2c3b45ccd041a6cfb0fdf11d0496760d4db4eca8f7f5c8be19f4ddae607ed6d6676701da9cd6846a913015a96b1210c1463c1850d2b9fdcaefed90255a3bf344fe0ddbd870226742f95a94ae2d937821a567bb9a9a3d00828f80359cb0724d9c70e4aaba5e924f18e29de6b83e20614aa47aa1a33f29c1d97f566482f693d0d366a00ff362c8433dc4d72431aa0e3a0ffe9b2e83a5c63fe7f39d2e1116a59f14be5983968adc314a52da338807f928c5ec837bfc5a4775201c17bbad9cc48fc244cf3bb6081c702993ec97db4341da8fb89eb7c09bbf3ca9c47bf24741da3903b94bcda804f3826d0cc3e291816dc6f8faa1cc9e7d1efa58f78adcfcd22d6b5cf2cba2854949699ef56ecdeb934c0ca89494c472805213a2ed5e37e1cc32d0161d359428416e3b9583c90b83a4bf4efcca89c0fe84f3f8571441bf55050c0a0ad01ea29a76faa7ba619c58c79dd0cbb4d7e4f26260a2691c230d65684898e2e011b68ddb429b3de7f3331c67c68523d8b417541d7947ddef2492bf41e005ba4b3045b92f623054e3fd508626544e1043828b993cc40865a7ba446d80ba8e1158f47b89439c3ab3b3bde075c0525b1d69d75361b0818c2d16a3931433d1e0bf6d30966ec88561bd217786b671ac33732c672fcc7453717a6c070073f1ecc573e6b16fe9e690853d446c821c49ff2a93228e8ab30d979caa8d2f87b2fb1db9392678c24b94b4c8dd6f1b45ad9ee19c16a98aee41956cf407412fc3b5910906be48ebe700e51546cc37beb47cc43e955bddd47d61a40ee56a5d9ef27194cd9652e21c1c727380d0ad28da61c7102ccf2acd125210686b1e2fb5ea155474b384843d88adfd5aba8302eb4358ebbc973f54a1592f41f09dbc5100d66411f65dacb95c736daef8a594e119bc9a216c7de279f42907ed3e576adb5b263726ea2de4125b7ce070d16f0b5a2006b9b97a70118982fe2b8b4f66fe5ecd7dc3986abdbc88c4fc184c4a7bb0987d9f44e1211ea8c94364c3a17187ba4d82c30bd5d6e059a06f72f06473af096e4f548c757db1879663593b939042a976b2fbabef4efb21bbcd0fe987c8ba848e66dfb4995958d2cac9656329072fdf065e89aadd1ee02de7ffa50fb2295089e60599b30c4747c11284bf81bcba5ef0d69d6f6b8f36e2d4ba101eb43c7ec261c61903676f0d9578b5c0cef323232ea4877fd285cdd3fd72a512b6dea9420caeeec4a1fd2ed1918e122a3c1661746211b6f55febbc64750839597977385c2f5c79147f8efd4802af7d199b6089c57f7845cd68837c175011c76c4017f48135eeaeed9223980337b9e2ee30f28ed5d6f312af89f6e41c05799cfb63af66bf7c3bc353c37ff446cb988f71a19c987a93f0fc2ff72408c38ac24a0749efc4892112d6a326a527551907b7fa28b5c1f71af117f0c6bd955599159cedab2b3eed056be4f78e4469526a4a7577d7778158b70c82b139203b5a7db3d276ed5449bc10369a7602e10a08ebc91e725c7878a9b6aeeaee3adaae5e6bb6b6e9cfaa95d56f51d6abcebac97510581d39d91ff4cdd9a68a9ef19714d333652c2da00ac1a426f882ddcaec8b66dae4f0db8a4ce1817dab0b5db42a5e2e761f6c6071181cdf478ee2f07860d6724965fee04765b431b1b24de76ac830eb296d8bdf1fe92c07fe3f69e0060f6ceacb2f4e16d10460dc9184cebb80301387126e94c75835baf98b7febb677a3478354c5d2621d397fb0dfd9527980b7893863f22cfb74bc029a45189f9e2f543b059f5c2a965752b86ecdafc16bba843d41c2ef2eaf3535797cf534ca7515b171b4280ab20101e3a47efe7969ce711032810d4a2ad9c3bb9733cffa7f32a3f6dd26b9582a49ff8b07392e2b4ad8b1dff6f1d2d440f880e14698835d45070d39a957a8d7fc3259d17025fa405125e6c40903049ca030f5f5c502f0e070895d1c0a81dc187b2577f17991d0d484bd519914974a9d00100d35db869672972c7fabfb0917e59ea27ec9e134bca753270f857058c9e5fe821934f0e3a8e12a2bf946b9f555d2020eb092bdd0419dd9ef00e3d8d608c9ec73b3f75e071f63ecaee7a9e5d67881c1b37d08b6b553e0f88803f1d47ad99a90b9693cbb04810269e63da8fd2a7c332f95914bfe2920b726bf4646bf3c6e12bb922f3228806fee60b69c051c57138720345e64ded453aec031d9c923935722098d1c5a507372c4508bc39c6e1e05f88c1aafafe19c155e9be39f1e743c8c68d02c2c15fc40e84931962c4ba60b85665f92c90d2ac64a0276f7a2c457ed0ceccc862f35b09c223dae7531ddaf70db870ab90eab0887f8515e00b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h389ca380e73fa2caf249592d368942d196b6810c898e96406c1db08891f91223e8fec68304639dd51fe43aed790cd44b5ac133dddf294f8b75f8e8a51d06c28f4b4e519de0c34b1c2b0c3c6704aaf83ea5d756d29f4cd7ad2077a8439d8ff0f1f86fc4cca7957ff59fef1f6a5ab8d1847e35fa17ead2e8a82d2b2a2b1ce5f1495a79c0e5c1acf5ecc09ded397b7a7f65cce4657d11d20f61d2f7402eb74b264057272b5421c27199fdd46d1f744c6457608a398979ecf768c3becde7460cc614cd86fd118e27135d007c71d9c5e781122b7d4fb4a6c802ee8907d67490b4ca9b63e8234643927880f275b6dbd494633aded9ff01e4d0b9697c61246cad2f999c8d15f0199c72c4927c53361afaff15b0808a12fe90bc75a6b808a9b49359c28c928bcbb0a69839b29a7387e9a86773940152a1be45c81f4fcca55ba7c4d73bdc996eb28bc3758641f090eedebb2c633fa0032d6b79c496b4c164e13f6746c965f6582aa9749750b33365a770cf23e153099b19a84033f7d31901a8659205c69e7f1f678e9cbe30adea4e0596e07a98a76f79071c6746a26319b962b6e515e9ac30dba195d6132487f1071f6bab1348d476ba9d120ebc8ff6ab797969ebf20241a0d9e167f555c50e1743f2a7a1b54abb5c7f579d76c89600f0b1cc8f097a12076f832ee8bfe2ba4e06638535ff60875db0e0ebbea59b7529d6eadde5ae61c3f26debf0adf30ec14536b82f2ff03ceaab3ef21a5ad17cee5ebc491066ce45ae57f27a4034b410cf1d62bf2b4f67c47f579dc1976befc173d0f9bcf2bd831e80d8a9b8113d00db7ccb205d1e16c1ff2cdac8e5f57db4b77dd517d52f3fd31be8e5200c492378518dd8cc420db4b3e1b97e6408572b742e3c2b432f5669485cd73e7c770c470e4de27cea818c8f233e25d04d6cadd50157e4a0a86bf2d0fe2bccf618485b138500c40a9d277b4a8a36548a03fca114176a85ed639481dd4f21df25c3bc9470d06af21968424123e2be81ed649aea50c77729f787b8215bd42d7924266a9d9a04b43e6938133191f4e0afa45c95dd3d0563e316d9a3f1f986fcd32f83a1b2708c338809a78a8266856359b4ecca96578a0351b6eaee21d42a18406703bf728f531aca8d0f751dc0595918470f2e3874c2460416d8bc4cc81fb5b675ffbd71cd1597864bf7ef1078e30d105802a3082266a3bc675a841c8a714168dfac090cce938db62b4eba87ba833c710acfee688ca6af116ea9bf38b886d793decd2cee8d78105de9691d28ed3e96d91a88a77f8f7b04a97a033c9e4e39c61b8bb60f675e08b675e31a60721f8a1b6059f218bc3d56580ce3ab2eff45fc5cb77cf628c8ccd48d01feea254286899bf36a61547fbcfb6776aacab901712c9b5afbe067abaf88a702ddf8b6866fa2409bcb1345fb4b0bef6cd998111e5b7d9498aa8b3fd5889f22fec697b080142eaef5de3098dbe5a0a0fb629c4ab30de57273004e6af621fc3dc5fb8e263fb22009f99045ddb799535487fba03fd15fa81f70ad91c3d87ef3f0eabad3d3b4204f6823854e425ebf35efb4e4a14c2874ceb6ac9db2e09dde425f179be619c5ee7025b08212a7d3d8bb1253eb641db9920ee3174b798cae4f51d8943cb7100586c596acfa0af0176c19b401e977b76b4909bd3b48ca8b0166b0898bf6982c08aa0dcd3bdd9084c8bb51722d7bf29ff4dedf1c5d840506f32f6f0442be29e278eb8f52afa4ccf45ebdd14a44b72c7e47d7a1cfdf7f37444aa797f1ff7f6faa790f39f4ac8cbaa8363b37fcebe8464cea6950369baddf9fc76f027d9f7b30ae9f09826fbb1a03c7b62fb6aa11f9a30985925eeff93e640cc88387756c7b379f5eb8d194e3a20a40e1b63d1edfbfab5b00ebd2115b14a670bc876d1f1d3434e963356fe3a2c8cfea024bc77f8e97822db63dada3cd1d414dca743f435404618de5e90656848a496b2dc05be39cf191dcf8b98fdd413ecb3e353499cb5e4e19201ace0528771d95b4d8c638f77c5893b9d427f5432ed55a2d3e778011578f215d6d2db9df43ae6792bfc5194f0912a414e28293eab423d0410078dbbe172ca143a24acd37c90322869ca7a249c6cd21f85d150462bb55aae7ed61fe13a00c0d37527a0c7f5c1c8c96c33768643da2650fd4d088884d78eac18352724b7ecb424ec1dc93fd1fe9606d31f2bfb726bc7b674204b3ee061af90bef25e35baa4c4d154e90791ae7de136679333a880b122a8a196e4c8ad5c1dbef176e5fa34cd76db331508a9945a8bb356e12d7bd0145442002a88553ae0cd7f19b8a797dba2e5e18260d4bfa065da5787fe47ee64bb83db3a547009e4665021929289b9e26b735dda092275f430b058865643317e1e11e664547546f8be8e955aeec5356bdcdcefe232569e809ffdd3194b23e6007866d0885e9a7b07de660882e3e792d363addb150b2bf94a763d7af231f70d2ac63408c1e3d7d42155af0e3a1e1277cbd6ae45b39cda4e754e1c391cf43a723f5985d622f171afb781c4c38c712d3e6997fb88fff60afe67d4002e6b99058ba6765aa740bf122ea046fecea6a2da9a228b15d5bf7b8b27188381e8279d1d1a7824c764ad20039e3631c1947e30a52675191069b37a564eb2aa8e052d62b7c47fab1b045ce96cef7f80604cf6ff0c0162709bc1d428024c359ff08e3105e40193acb61b277d2ee017bb0887da7b87d7ad9d9179fe795910453460976e0f793185f74e188d81497597d8944e184b38f25bb8b8e124c6f55e15d1d32091f88890b0329b260102e48fd742d2b85770ae14812dfd77bcffadec1eadc4bd37647f9526fb62726af2db5187d2312e09c995801478532f8abf3f26ca0758dd19f5c6fa00a55c2ad4b9d0e2256e71db5b6082b1baa7f4242b30b1635a612d39febc2b39ef159e1529181d13d6797692204266e239bf64ba4ff6406f61699082f8e5b52626005398b5ffa98842f3546274849ae1b169cafb006ccfa86959dc87149be0208d633dea2b408bcd3ac88fe0fc0c2b8bea396de3ba4d29ad1f6741e08fce4625f5657baec2367f37aed451b2213c1cbc29c1646579a866bc3f57c83b8e0af3a49eb5865489f8b5efa277eda23b597c42a2b8aa2765770654966386ce5767af2f08e4335d5f76f5f961ca4178b6b1f7aa4ccdc8bbf0e9bd2242394dabd2883367a9a9f73891c152448bcc6df3e73618ec157c3e49f2731fc4609ef5b957022e22dc6dc02ed2228cdf06c2be97bef8abe13b5fa008b0a4c0720afe69292a65dcb6076fc239fa113f261203bca6942521cf34cec71adb1056aa5e395e89e5996f6ecf692a5ff221be4eded62156e2a7cc44841bd54190f37d427e925a4b09e63f15027eace20726dee8d724804b322b54569625c1ee8e756edde7caf22d576d5a6fb5864fd9a13323bf936a3218334021ab1c607acf4f26ab77d3a0493a7a082f63c683d8a205a3c3824d6bf9821b5459c6141220ac1b7fa45f1cc8c21d1e4c0b93478c99e3224cb1a78e8ae7ee7b1ff272cce5137695cbf871f98f0a1692fa696935c26ff3c60fa152d9a0c78a054c4dd3bfd1e7152a1d9e5ea02e43e72f581c4a9b126d1a30eeabb4e2b443c0d041bbe87e29d12b9da38915561b2952a2ada3a48c6d5ada147dbdfe54ff2a678939999d6b813fab73147ece22e130760906eb80a564e4be63d684b672b57f478591741893fd91ee22fe3c934127df2bc28619aa4ba74c5b554ad0f97167a18e93bb5d751f7dd09b712c4e23d2c9e0d86b05be31547cbd79f3bf35c2740d6186086ee0e1c29a77a8c5528bfbe23cb17f868996cfa27de11a39846595d8b39d1cfdbd865671e0a938e20e49686bebb465880f5cd4d7f2f0daf27c09d379ad8947f932229a4dd7d270a991512070b6459921bfe93d76522b625c7fe68326e6795b43562a8f62b8a4546a1aa94f6f87cd09c7c13f4554c65c0a3d94ef428ac4aa84f842b8a5bfda82ee83143d6dc516ab270e3e98c5d36ce47dec746cac4f03ee0f81130cf3812b2d16e8799afe60ab7408eed0c08ff432f1cfa5c44903a488d1d8f1ddbb6ca799f8bc933b2b6df0a390b01873636a625d4cc0786ec7bee8ab2cba014b1caf6640accfb69f66e888ee9626d0b0c5a3f1e146ec7674766637bc83721741ccbe619877da2f4bbe41f0768da2de73358e0d0c5db09bee587aeb1574a6f6e425ff3c9a738d20d233266ee142cbd6fd566d1da72b5fb2ca62ec3b0b085f888a56b793805a8e28f6377b4f2aaa7b8d6077589948f2aea205063d8c91087abf208e9f3012d4b45e9935e74941941cfc371a84602a105bdb7f70e647b316ea2d24d3f17a5792000511d6001080126526446c61c7a91165d0fbf84d7dde1b71773eb9375ee7157ab57523a45dce5457a81c94dd5421125224305d3282cd3d9a4c776134700ac62675a0e2e68abd62f6991edba60ea3864856df2601d4835f69dace7dd8cb705ce65d01c3a23ab8b5529f48f94bd22a0ef81a7421d2cf27a1140b27adea19289ace8ff6c55b8c7b337c25a5b1808ec994df92b25d004755482116aeac42d15b124b328511e4d4527ca4226c2a9afe46833312035fb4aad49ff4641c4eec975600e2845ee0f38f6e24307d45e20c39fde98b50ac8fbe9ffa229e2c0939c4beb07124afcf5d1d8da1c40e56d9d138750de19a88bf569f05427f7dcaf507d3ff466e64116083c25e91a9ba244c48e3ca7a01200bc28033bc7f561654a945472c5155fd24e61258e13487c60fc380907ade3767b90dd02bc8e428f6a75c044def7f53094d311204859f4e9023c8aef655b695e5fedbfea551fe685516a39db2a729db5dc9d7f11eae7d78e15f158808183ad66e70d69ce240db3114a308513b8772246e51e3d793114e89dd3b98633a8164cba760c29c5954e975dbae0cbc7667cd4bb31f687a1149e830122b5d0b7486bf05f09862a37774ddcfc2f8bd1beecba3ccdda8cf1aa3cce2543b1bf7dc746f06bd5664d375b7d97e2ff07163db72e076ba160f182501d6dff54a0eab1b584b04999e7ede49566059dc35047ac6f018b2d470707b7434903550a70fbe0243f6b580a87e848c130e3ddad9a1e3d9487af0ad52ec0a33df272d265f2a8fb10e74ff3207b0e4fe5174eb1f6e30b75dd6524a154e237ac9a82a2313895b4e2ee530c20d69e55e0559ebc26993cf14724c0854869aefa86f18c1e6c0affc3e3ecaf326ca629275fe252d8b163a167415cf37d78cfa4fcc84127f43135cfb23bcbe62208f93bc57cafdad589b8520c5f72e986624899e5fd3cfb972a46648eb6af14997c8ee37acd705b418cbaf9d3e768517c56dd4655601c2111b544dc44bc1533ba6dc83f785e6056cc53df677400c5bf52ae45cd70da68f84ae38478bf07b89396357f5c789e67bb1fe2929acf9913fe9ff08d671356bf81c6abe4464fce9f79a354e17c480bddefb74818ed8c0e859c7fdde00fff1b208a80b8f15fb97f90ca19d31f1ef5089a6a4723a9539e5f7b356e9ad55eca8342d7daa5e9f016a7c069df2830c07974114167d04f1401b1eb95b5c212b8f0d49325dbab3a702cd1fa62035ae20ca6c180fdb0b70215a51cdb90d63e3cd153e385cff3280a14381aa06dee530b849622af332b4dffb114bd5b935dac9fdf71cbb4b635a088124cb6d52417b83e01ea9adb91d396e458a4e062da0bde750f5b146a2d23b45f613b615559608b4a22654cd6d55c88982ef0d68f75876c59bfb850cf84ad46c8fd97d3a4bcb011a576e7c36ca3886c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h17ff4d314b515c97dbf24a0bf93939b1ce89efbbf21dad821619194898ddedfd6e9c20a51dd62491e75745e9c9f8c16841c1d33314a20faa6cf9d50d706ddaca99fbc28d67d9755a8f43f54a9f158b74e6de98f4a8971a7e92626fed02c3f98ae628d47f1023d3756bf6396443b051e6c120acec35d4570b99cd3b8288943dc49e5eedb0126f69a79c5568d32422661cd804f485077edf9872b836f6706d0531c767303ec5fe7e2f95e87c64ad09af013e654339193c2f46990b7554554bafe182fe350f5587eec204bded5156105dbb8b85f569f966affa7538701597c4d987a1d1ef4a18316d306319290e008ee0cde8e8ac03bb8d25ae8dd7202669a66be2369d4559e5e0fef1879d4a3eba7e273791e04cce239e2cc2b8262c7cbfa14634a4b5376081da645e5086aa9fce0766bf27774d682638ae81f22e7e88ffacc50b56a26306ecdad4ec03f711ae09f7bfa9db6d4ebcc8c5ac20d88c3abc7330f0417d3e26735aa9f5bac9146a34709b00e86715d7803847e8eae12d594e1f2b424815eb731bc01512f2b80ed6694cce716cf5cce010ca73a1d96222d53d93a3fbddf3a7235b2ca5d03e2c5c2794583fe6f267a6fbd396e3d863d4b09bd20bae5653c9652e8586e76333ee8ebec867fe2859c9982f502f95efbc7e3ab42c6f92530e7a17a114f4d6c9b6f60b84caa57b778ba22167bf79c8e2b2850f8dafa26af67b846f921ab3eadecae4d922a5b841a28d5d147ad3246fff1fd739c02cc8910a544c07f786c43097ce4b63ebbf93c74853ac2349e895dab29f818f62be73b7b8bbc0f7f9c0a0bf76ef9643cfba2f99e4ed3b7d41aeee21090a434d5cdfd6fb13db903446b13cf414f5de7ca567c3b770285fabb51be0423f0cd37667288cf842b13e06ab170ce93e818ade367d094e5e2e6166e170e54ec91b02b171dbb8421f7403a2bfd13f68d64e42498d27b519e0598db05ce41a34fba7e17fe4954f3a571e60a6b447fbc133502a9b2c5800779e74c04e12e0d4a210d1c2d1b59277706ab6f208abd31e1cff2091efbcd031474a2e44aa82de04b1bfac11a4e043d8a14a0eefdfd3f5b5393ea7fd1f1d7b074b9e622caba9998933dd8f8df8bb0a89ce49765da24c4230e9d7c317a46cada5f569311b2831fe516abbe6a8b035dd9796eee567f2ad1f7627483d14231ce00f24be4248377671d99efc82bf1447aa80d0f996c15539a2ed06ca0b7622bf9609f509e61f6b5e28d555336e032fa1c9ee604678c21562b6fa52eb0151e8c1a6efc881e5f03cd0f6c0654b1da3848d653b2cdca9d9b4745ef3305972e38f90dd09c20c72809e72092bdc590a2936499424c89a090a74be14ac81c5e8f72b20284b42bc2416f1bdc0d762057f980c82a843f92314edc7589ce2b01694bfd12a774fa6b53d677c26974f7fd7641825302a8b81f328bfcdedb7defd1c1e752ff9540290ff75399928b39c9c051810e879500716f2ff5e36e86d758f6c45e24f0fe76b9e893daecb2a15eafcd3a606a66444e8a1e01cb989bf42dae9b31f689b537cf8e98c638c32f4d078b9969b25b851142c3b0b1a8e5f54019acc0b85f6a078ae80fc91ae850b7bb4c9136127d6bd68bba0c0c2249a178f17d8b46e3a9f146a43313aeb0cb2040a0d6800a5e1373042682c67ba59f0759662d9ed0afac06d52c1e5d2fbeb69c3ab6ed5108758905b02c8242b4cd8400bb20af867c50c872ae102f34f64c4b606e16ff95b62c1591dca1db782f19febbab06f4e5cfb94d194b448b9091028a717ddb55d8ba8782b45f49a889f7c1aad88588054411f13f3309cdcd4b4430baa650200dd884a996f37aef939ece06a11aacec39d23014975031c6625a51587c3ce50081dbb8ce26a788565fce370d05e38c06bd4800a2863a924ef67da272f0b92cbbc33091f0579884a5d81514d6788c649ded122614df337fe9a1f586235c88c8f9878d524618c3015067c6a27db6bc815cfb60d2b51e7036cddf490f154b4dc70a6cec86c0a9646a93f829b9272bd45a7b91b4c49ddae2a540ff6975beaa0001d9612993ccff5cddc836675a97849390ceae927176d3b1527460ca7f86920eea68aa90568dcb440243d895d6259dfbd6648635780780650db15191fecd6a2798332e366d7a61fc538f5ee5dfa62b1f7d3a29957ea098ca910f3dd83fa966abf64feadb88f83db3d10c447ef861116b071fbf3a5a3348b08781dc3d39c2f5758e5b27414f5e22e5874e1b7ce11483e0f1f78b2b4f379653f6215254bd1207ad24098396cb23e9143ff8f4645b063bedb240c8969c3b1722724a07f160b73e10cce5998f2eadf58d3125c15e5d593d72c862f3fffc034a25d25c03c23b62fb256abaac0f6bf713f0ce4b493836fa6188ad0eed57309191a7cf09781acafa9a23ab22400b4f8b708f61b1862358926f8569cd74272bb265a7e80d96000a32dfb6f8f501b00bde5c4a9a8c0c3cffd7213049b270dd673f9195f1c07b11149d71e8b1c3550cb6b57777099c6e6e28f071b3f94022630f773f06cfcf5c1ba48bfaf2db849c6a04981ff24dd6a32494a40bcb811b42cde6d2aeff18f6083bdf948e029a07edcdba8d32aaa3bea3bab07a7174e508f85c74df7c067f4fd60856187b31d1d1a81675382e3bbab6f69033aee6ad22e72d22f786e4408811b62397cba0aa292e164bb995dc5be55af51fdd8a0079f28124be9964f116b7cf77bc645563eab06582e4680257f8fdf998093d97afe65628cd655a0bdbc23011e66efdfef9ce5b70de7edb07e4be6076690df102409f09e2ef16d4144cf862df867a5e1e784788b4147baca80c97e9646f3802f35bb41cd53950801fd45f1cdc04ad078a63e3cc3de4e6acc43c98f3637657704eaedc53da0301215c7901543c8cf7b8791d1d9d44be860ffa1f62c3d1990c7588bff12439ea9b15523d4fe288c2840820fd04d8601e6a8d4deb4a4a461b24944dcde7caa9f4aeb7729055e9623a078e8e24cd04384a225b96ec13bd2e51797dbf438db0d1aaf946f147b5f70dace45fa094831298993439eeaf3107951dc04f14a374fbfb47843459f9ec65f55415b590e3c5b15a91383e211dcdc8a4b30f6337551057f1c724355c543ee631bf2cae992aaeea014cd196623c507f7f9f41d76d39b14961778be6c7ca135c165bae69038b881842e9cec3f258c627558f9cbbebd154437dd809e297557b4a6bf15767e079e68c08deebad473f0f4e054608af11ae0e7345ea8a8a35cbde93498e76cafc3ab0ef8fcf0bfbe82f3ebde32b33dcc56ec15254ad8b2cf6e5b829ed0d19c3ae7622b51af56f2bad61ac0c5a0ff10cba5f39d9f953dd3ba154c48b4ea05478f46797d05b4e53962b3f52ce0658b099dc74da0d95dedd882c09c7da9a6e0d279187e8110ea47f550cd4174c05a862620f68c3bece26ca35818e81d933b8c1c119c9efaf6af0ef330daaba10365ddad23f3e0473cd31b2c8656a0f5ba5f85d8940e5f1f9c56f119db9b33ad9c666783a5d392f5db4891a8580d7985a1168bc0c5064d118728ddc5d6823ed4385d78c874b363be31fa16a21bab56845cad5b0ece33ea17dd1223b9510bd50f302543b00763b8a2349b710c0aab027c0a2a7f647098db1540baa14c2bc9ee3a986e999c1125870f40a9c175dc194835364cb25ade4e087d08eab61411250f090e3ece0dc97cff87a2a1a6dde8d75a2d2be5ef5ae2aa11226406b487824f096e04660a6f9f60fcbcd140218bebed11c60e3e517aca6538d7d7e61ee4fa4dc31dbe157170599df1c09f8edde2b56f15c0e4fab9927ace2dd7761f1b930c2d784e7f6174b0db7263bdd2e9dd5dba12f8fadcd9c41f03cfca9b2c999561b0c3932bb6c3ec80bf4b61395bc5e884c9c3b423ca8201ea22852b7a2ff83c15e1fe762d6a94da3e3e38c0e28b4762cdc0e46a7f7e4c497af3110e47e90daaa14a8443604c094a32767f1398728eb71c764fe0fa7122dea76718935dfe654f9942de87db3ba5068f3e1ced38758e6fc53e27bb0dea48efae0089dc1784b641aac466b8e6148fc4db912ad3be4a334dd909d515de233321621c3dc0be6b761394009e30d723138c187d3f83abbfb30582a76d6cf8c732dc0addb5b77f203171d4ae8a53459fb8ba3988977af9db1ac617b45c18b3b70dea325b86a2f185d049d7cc3b92d708cf58cdd0565c5fde7499e138c1f628b734661767fb9eadb9514b7b7c23ed9fd41e98bd4ade066e1cca161f45c2329cbf4027be9678cccb4578cb87afb86cb2e547b52de0dbda6140b1384ce59de9a4115fc03d1505dc0bec19df4ff23215914fcea0eb17d2594307b2dd88361f3f728283897da4b28f3f27967056f744dc232ec0556ccf9320cc6be8ed65a0442cb7d63d452bb45133d9be70218b1eb19047b12fe4dde8652bb267b9b1988c3b3273e96361a486ef2a3799b309a4162e63dd97927247ba461c50a4f4d22bef3dafbf27be133e31284f8399c3256f76f50c20f69d36059eaa5b6a394315612b6ecfd9698967879e629014bb0215d885ec60384509bd48288ff0b818548f72c3cd1e0d73be8467de36842e5b42d9e163a9014813315b8f763b7289e78f56a73f49469fd83af246fd68cdcceaec7ae3e7dafbad8df146455041c5d303c17d2fe6f7259a5235dc91611a53d5179b267faa88ae21b096e2feed23738c0c8eb51c42cef819f4d7b3ba6507c6e2183f5a5644535fea010d480bc9d94e10fc2d13fe269b74df03b43e4c7b1a6f24a3b75941b3388d84306e4d7ca49bc4df4d0a2a9243dcd93f54b56ee2877c3fa01ed4b479b32c67c02e0c49a4d6d37a592f026b422e66f3a6006da6e87cfdfbf0123f1748806cf763aa753f292e15674a556a0e9705c40cb1eb5400f7e3999bb4cfae1a9effa925f65e099964706a2436e7fcd636adff3c96f89ffd06a8fd944cd69cf21ca83973c2cc293c723cc9ade9df4e989fb16248944673c58f85f4f198e8328549b3d66d338914a682ea49f3008ff7b70642302235c586a0eb90419bf2076a31d4cf102b972b3e1f66ff04d158912365030da95c2a7b0b1dad06f82092ec487f84a7ea059d1037705aa71e2a532bdbcc0b5d3dab03004a8c2c6c89144d7fe5e988e04dc2d4111430406e2b02f55ae92d67a0a640090f23f984b88c0debbf0c25bc03387d85350697fd62adbec72197a526ff870b6ec675abe2abca1607202bf50b11cb34a90ae723615ea2e2282d5216c00c6f96d5e84cfb0b03aebc2dc8eff1cd26a48f6e562c2472162ef82e78955d1cf0e8a02bc7e7acc8f44415e78511408ef8b8255a1de48fd8ec82a878b36662b2f4ef3728a2ec86a25f8bef5cb49b48aa68fb48263b7970bf49af2716990b8bb249eb7c57f9b9a1efb636bf97604a451201075f2ef958eb6beb80c245181cb0879c857bdcd644c087d39daa93c0218af471677ea8217b0b17713d2f101ef37b30cf59ae67d20c67dab3f0c1758ca9df49312a4b0394144b8981a82bcfcaa8537d0bbfe99edf1792ab563bc378c0b1e9675a134fe5e5a3f0fb58ee3c04a857ea2ff05534459c2e35f3fd13b160e27d26f8b19c8905f6682d887a96314e2acda191d50a736c3a070829f2710857bbc4807839ba2770c4204ae75bbc863b6dc1b82c4bfb44b4f601c8ea578ff2186ea0545fbeeda03cb09dd683efa97e658f1087dd781b0d48533648888eb07f41f40fca45edbd2e9beb244ff859b3cbcb31f8cae2292edb2d7f748f970bd9f77362eb550760f3d72c994096374297;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hebe95b3afe39b9ec9de4f5276b90ef329ff7bfc3ed4457fea56479da295e67e164449982933365a27ca820963a25f6d15e6ca506f61286ecea2eafc4d75ce5b429eead8784909e7108717c498a23910356db2f938ad87bef541beb986bbef60dbe7cb610d46f4e15eafc9bd81d3433de0ba29e258c55d688733185401bc5b0b54222afbcecc9f3e5eaa64247eef8c0c66f179fcf9f38bd1a0d6d15d5839945f4497acb1eb4929e32d8395fe09694b8e4b9b3c7c94347d63e9f0feb0f263bd6a07b143f32936f3f20629d061516a3112955c174ac28d5bcaf30b6d1553673aa2d0cce8319948d896b01e85cbaeb6a0c3a3df4d0e789828bb91f02c3b1b1dc760cd8d0a5c09bbb7ba03e577ba69a8829d620f25d2a9514ed041706659f8a7cadb581dab62fd5df6f0f3a272665b873d508dbb83690e8788c4be0bb368bb54c73c1f6ec54663551cfba5ddf9f4111a54f8dba7b6b068e2ec9378d1ca30bd609ddeab321c60711c303e34ee5576c00c840bbdf31cd45869cb5d7f0b28ea731e39710cd117ebde8a2b173f7ec688247357cc6af040ef83dd4f1fea821e7416dff1aa40e640450aef52c7e819294c6210b39b7605d4532d196c88e196f1aa0c2e1d2cc87fd950eb71180c0ce4e62aa63fd7249401e298a3e5ca080e3928151139f92960dcd584d33483ea8ae10684ffee2c7e8d5bf8e2ef923f09425ec60ae5e454715378e46e95cbfea46f3954e18caf2e4ac6e715c2e1ffe6591fe1a97bf22c6cfa4c484b795f7f7bbc3aaf6f64e901cd254920b0ea9628f5ad16d8951b90e280b786d353cc7b15fea81d923a4932e90fe3a67bec5d712531f37c8ac9305bb385c70235762c997c8e5c6ecba846b5a3b02f5cb9dafe807b2fc1d71aa6435fe95bdc4de6c187d2452c0342e04cbc95f72702d1685a0379498df6efe7fb2751ca82429794e3891b1ec1e4e637cdf38fec9dd76e6371639fecda47c4790997471314a239c7f5ad9ed66b87f2b067d470d3b9cb5defa8e437037dda48a135e3c99c8c14816c879ff625adbaef33c90f973962efc4e9e12924539cae3de556061e6b8cf25784b80dd5e87339a8c81c1fbf75d11b92ddc14e969b5c163a4f6d6762f698925107327106f5f29232b7020330b188dfcaef0139c4732eb7fe9a290d4fa2f5645877d2f328f5b134225ecbb22a5c907518664338284d8dc2b49aadc4e6de0e6d6aa5491f95dbce713025105213533791f4a9f38efbb348bdf0a4e46daaad8967deb9a4d42eab5186e704c7a818ea7ae904ee78eb875b4f9f9a406e09d341768816377b0f84bc0311762088d8d6777b93c8420fda2b9caeb51dbd9524e5e8297f976ee842c3c23343bc9864d67339ca601e7443a8c57ded44697a3e7e68583c58f24ca6d7c598a58f3e32e0de640f7bd74f55200a3132814549b94da7ddeca815d43cf9036fed2e8d451c22252a30be856a93aa774b662732d83c7d033af5c34f77283fc7f4902d5d1407ca6cc4a7ad63fca048ede60db59fc13634d51798e815f9bfc1bd3183fda8ef181b228dc8053795f163f4d14094fac0e57d46142d09acf3046d44df2f572d4823f48c678767b67a625bf50a0a232d973292b17d9b87faaef2ce30995146cf491768bcc9714624680577d6b033329f80300d7161b8ca777135dcddc09665afa72e17d35312376cdb9bfa2247dcb2b10986877ef5034839a01b9bb2c12d3d3cd4903a16cb7ab4af2bf7d1c24ce2ecd65edcfaa1267785fe8a0432ec2f7ee0f8f680c7e6ca13650912457e0dca5f2b8b6184612d5598f74fc541ec856e74de4bf608d014456800c73864735d7ac049c454f6b16a09b41c27c105dc3a964bfd0ccf6f6dfd9d7127531d5eed1ea5b173c2c2efbd8c792f2ebd408bcf644ec3eb360495432505f2860dcce31036bac7256ee3c457e4c6ea861f3e495d5dec32e8906d2b9b1d5902569814bc540e5c585d45ac9e91a4f097e82c98c0e496d5a9e2ba69b04c1788e7be52c82f6701a3551e6b659c990779c23be002191f291f2ea425cb141ceb1f44887e5bff18af9c06758c6356df6e57da8416a44a438598919def4f0a7655ea2de620b2b47f42220ca4299fbcd760e9ad309eedaead67379a0927f50a70495975d7a7bec19eeeabe32e8180b856cfc769da86d539d90e4ef5eb474182132f833ec5cc30b473f8763c1ce5da7b8ac56c5f61eeaa89cf4e8bdb2039a67506fe5d6c1ea20c187dcc86bd7579570ee4964f34b07e5508e808b8373fab72b5cafa29224ae53d8ed44f634d2288384b666cd911d818dc82c4b77ed0a2683c2f89c0e36fcb994e135e8f5c938c80f2804673ab213ebce56d11fa314d0ad682bc4b90c57efa77a9b454290c45ea9a7ab9a10f4c46030b97f3487a8406471263c5284be77c15f983ea6d02c7af69c62ab56b9a3c5ddac3d7a01d0ed49908c9847b5d25ad0fb2922f4e5074320ed78eba08faef2e524d3f230f04f7820a178bbc0c6b6435807a565e23613cd2094d9782e0083335cf51492d6c12d749a7be80adbdce78c305f0bbf86bb857948501c7bd51d5629febe518db7a67a2b5dd86ee81d23a79eb2506305d63c534deb26f5856c16455758d6f197d8fca852baa71eb998bad4380ab20a2f901b72c921f2cd94ff9a40682bb9b3244677dd6fc0bb78eeafdcfe29ab4fb4f2123949499b7fb26bee5374f6eeff68bb46086856a73dde637ff68413a45e072eac2d03d6d8b0cebad97034cbcb0f6d58753e8a37e888ab2fc4206a83323b3699731bed78e81241ca587bde15629b60a33e1b99a611ffb38fba4b0e37c33d2319856145cff6e7ad73c17d676304ea97d3f8354ed6cccd43fa96c27fc1b0d6d11de725cb07c5b2ef8702ed6f311111f2bf29c454b4217ab412d626235eeed1966549ee62aa0332db43c3ac784a2cb659c2a5b73092735efbc79b0d72b9c8a029089924bfc791546c71560876e7c668f80ba604a29044fe4c3959f45903e74b4178812452c68dcd1d0beafe29acac6b760a32f71852314aee34d21b42560c491731079ada22c31eaa94ea4ac5580b503efc268b3948759c258af74c679e0b4638273bb328190b4c66a7d4cf9ba161a1e22cdcf2e3a3e5889275f3d68188161ad109eb486a1206d8496b5557942608a5ffee0701562296cba8609c01bc280243297bacfab1fe6620fa061a03d192ca35fb57d0436d3784982b00107fe9b452d13482c9bc474cfded57f1c3c27a560795aa1dd0a2b46b3c69ec910aa9a327f3231a4511e3ee113037ea2356da9229d93087a7b2470535bc0fe3184f2bcd28ccc30894ff4fe95b965b228e2df89689998c8ddbde18ca6d4e181c0b0834bae5ae4a398cbdf172b91abb5bdd81a49d9023a7610aa9ba5b01b2a71e9e128c9c7ff9fb2030de25b293765686a704e9b8a119424aa2e5ef8dd979174b3ee1f8827a8eae7d9353e69b8f4ba134cf8af2af41557fc6f749b72fd5c49f2a012b729f5d44b031fbd00a8895f16282ef58ffd8e6e065986ab8c9986629caad6786e1703f0aab435ff49a5da041dff5ac0451c966a6e378ce7323e740b5dca0db33bdd5ae5f5bd14d24b154c1a7630d205ba6ca30990945e4fd262c4a648ce57929b0e8e7595c02d00b6588e4cb7abad306bff9310d20a8c46d458cb0ef0521b2ea68429f25151c932ffbdadc56ce60ea3aea0f659f667899aa7ec845ded5c3911060a9ed9ec93b670f6f1fde76e64794b25bca143833375c37f4daeef7132e1e54e7742837359aec2fd5bf73f60bb78a1666c5550a9540ea42f7e648d987e5cb7f7968b5a891deeb7d1000497f17a86608d165c46905806073171b7508403ff3d95a8d2c7d740af290453e34d629ee0ab8c84c74e81f6168113f57bd895e1b596e0308c421cb6376248c4136889b49cf73cde2bd8c7c4135a3e0548dd4928638cd70648da9660f98bd44a67fb29d471f10a56555a1ad1773caa9410156ca2083ec058f0bd24899ce5ee1a564e7d965861c6aff07d00ae0b6c243b6a508125029c5c450ebb6886c1ce3940ba72dafd437e753b64b0d9fe2a10ca4c700f7da239fd0fb76cf4f1b816d0615a17df6369e58365a92fbb403f86bd445a134ef66afdddf6a19d112248a81f6b3cfbf19e7bf5152eb61d93f69eb95ed3000996dc20967aabe767913cb30c85e9e78fe453469bdbd42034468c685dcdf349d1138b8d0dd97c7643ba7700d720e7df87aa41733be538ca00b3814ce66585ee419f65794abd51167fc31186821ce5119a2a27bde20489dcadc902e9f8dd7e2c88eee1b7bdecd7a410585bc62b8e8938d3339c98b21409eb2ac395785abea80eb6bc46492ead0aaceff6ef99f7a0faafcacaaa0c95b53bbb1783a60d5f826eafa8b19e0a65b325e9a5b7e476c08da6c37fec9764637d9cd4a510c6a26a6eabac3512c0e4748319e62676b90ecf5d5591cca2240313aec51c0e2656db97e159f20de3d8519ee82b5541a1dc94e6712a79a74bb18f0b180f5dc880d9ff5ded30edf066b380facc9627afc47489a3d6dc73bdb078e3a90536e09cfe9ccabacd329f0d90b8e5d8c82c5dfe69fd1500a5c786d79e6840de2370996bc74720f01023d9968c9a74e2d04c655c908b28552c58c5c3475215121cbf6f157cdf3f2a746173a67093d622ffa732d1772613ccd225cbb2b721034049d9988941b7b332f1622fad5a178c75f61ffbb1ab0061e52bcf98a8cec5616e92887468ae14d43d1c9eedf103a742c5ecbb4483e017630120b2ac8f4a3b7645780cb28c020f6e025d6fe4a05d033ffe55a93190a92b602f8954711fdce383299fd888454e76b46b2d7db7daf41ce677428c2a7c42167155a7332e0d1b4b42cfc753951c3640e4838b6480eeb0930fe020e45c1c00309666d4794c8e26388a46d8b1ef124cf024f8c15d3324a5be82f5a10e76b6fbd0be2362d89f06454a550d3a2dcf334aaececd19c17e17f7c56516e949241b0d1abb0288e829a29fa20b6165995d720578a0b61ac2f8fc7bab24e0442bfc069ddd28652ce6c155cdf76513c36236bbad5e8920f038f62cf5f7dcb496c5a9cdc671d8484807fc6e6459de69c9b7b8cca0b1438ac14575fda59daba2138c18842c30ad2861ed8bf5fa1904d55ce5d7d235f4c6ef507c413b0b3a2de558ec17ce776e1708952015d841ddea47ad9de54b8cb653d8fe2fe70774c610a59b3e19c2b1b533473cf9edd129aaa4ccd0dbab8af8d1e2f84693ec031a33e01f5460072960771d49896a413b847a874e43843eecfe8630de9a22e287948aab5c03b5871e9cb2c9b1a0d34029f1d0cf690a153e862b7f0a2a109f68fdd2364617ef32b9348e4fbe7bb661285b31ac8d07bcafed09cf1a9c89ac53da009e8463570c02e52148c7320a3c121224dedbaad38aeb2c3adeefb00be16460b4edb67ba4e03274040f04214f8d3862c4b2bb36488291eb4b0e651e98ff07f4fc37caad6db092345864c2a6b402fc1da13a45f04eac3f78ad8569cefe02154ad9674136eb8d0797c579106cdca09c8a76ce875d732cdfd35b832c23c01bb92772be4cd8b4039f3236f65855e89835c59ac225d53f12f412e006ca207f4a8d4f8c8d27c3c16b601020aa36275eb4cc0a4b8e70d65444e7e9d8050d5ea3ba4d6b22f094afcdce8df4559744e56bd2188dc8f7af16963ce6785164e5e7ff2f3f06cd71e751220e2a9c2205b5b31ab9eaa03129cb2e303ec8c3e1ce021dc38a1468a804b80627e62b0f3bf8cce6006b4aa88d0a73787d827830f12e3c34bcb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcf63e3e399f07b442bfe6da93e072b6240c8bc8da73e1816524a5680ee933cc57c7a5f5d91921df5833c630d267c9739dcb960bd1dcf9ff0677c8bf20ef2e76cb7d10017140b7dc9a951335ecf8b4297c220b75d497d75ab65325b8f5a3dbf4dc218c845b4f0f2bb7aaed35a814c733a697b34ac540734c6ff37e0c382ff8720be3898dcdf02fe6eeb59b6018bc2fed3706b0c611491c20697414c1396c9b9e7a6662873560bca8521d0a56ae3224c6c92a8db01294433171d22b955d454094a2ad7670aa6e2a8ebc51c04dfc30688283060e4ed4f603b9e92b07af139916bddec156664055cdf1ece171d9a44461f848e35c4ff4fb426b92550c56f7dffba1ca8110befac2755fdb4741a0a5de0365e75d2050637b6612c141c39d1167d16b18fa2ab057d85e4dec70970aaf50cf3ffb35e2e1c006bc3a18cac537237b1dce31e019a9530914935f1da0b6066e4315ec845d3b3e4d82df809836e165b0cc26cf054e50262d604e8fbc9249aa2a2de281ba255fd356cb32a521fc7005c230429265ccb46cd52c1f2af560b92a6372dff31f24d9a75f1630d5ae836bffeace883997541cbd62b95b8c75a480af3b20a6847e3e2469198c9503a87990c4751a214559224ba483a33bed66858f5c9db31d3f6d0f1fe771ab780d52763cd22a42b81ce8c8ee10548e31fee8a882bd274f5de7e7e79dab8277d6df429dd2585c0a43857873d69ed68d45d524694ee32328a0753af7c774a755b5147ecacc7a54f2b49d6a40f90ff1fcd036bd251b5b5edcb993a2aaca525397d4b8ebfb3d664ab1bde5669c6e55b3d60827b23c5457e8f9060df2fa719afa2b4c6d7b15dae232656eb7aa6bbc3a9283342d2a7652dcaa72bc75fc5b2747a80d71ecd936306a6cd3eca6e73942fa071477e70fba34864efe43ada980baf41030a9db8fa85eeacb42c011807e8768fbac192f944ba6ffb9e378dcbba5ba7243b72b53f7ccee238e4b80dcf2057076ca53ca29a4f1093c56a6c3ee4c31d7c5ac7bc845787633a3596b32fdefdbddb338bfd4860edbfe54194bdeda919d5892a80dd12098f9e264afa936fa2d730e52e401765e6708e440296c1dce75aa749e4d929f8bb78ea7b1579e203301670f88e2de672f4b8a85511953e3dc8ac84d0f7df41459807da6adb1aaccce81f34e4ab12e8b1c60a654b11f04e66c860951f4a597d5e9eeeac0066f9b8de669c0f4c67c9d04006d62506c6329f49ce6af9a6e030f44e56535b55c4127e8b02949174215080ab410225ffcae650297533984196db746be4c61e523403d9f16f64f59c28bd989ca670abab05fcb62943fc3adc105061384cbdd688519ddfb8c5c5c67234eec6e07c416ac038605a59f39db1382261f006117c56f8af8cd9d09e09e5e3b0004d69bd4b811fc6fd28f222e3c3ae9bcebb7b11a1c6caa6b2706dd8d5019e1aae6e5e181d99806d5a20dd7e58d02b32106657358a527c6d75060ce20016f3dd124c907b8713d42d7072ed9c8f5e439411c64ebe6d623c1144caf20c9ea2a5aa671c2623093b6ece28543bca830a94921fee12100a94e4d11797f9627fd2151ac4a243d6921e63c166c8db69702c415d1283e1e292f7ba8f9469a9c931976e29044d440711515859a949639f65569dd3b2c2bf81a8d9df6f16496f0c4bb9d261e3de62161518072c7abb41e67fa48ea11274c2ba662b54f6649352652cbbcae28c549d58133f22a90ce4d8156f53d34c5bc6b51745eccfb820b98d8a345491ef17ef12d6d50e7be14872ad34085c14bcdc4e48e2b3723d8507f5ea80b6903c245b586c7ea178486500641196682d2ffee3dab4835f9c9514f4e69baea04427d69f93eee834a8f1e1b8290b9cd03d463763f7c7d0e650f7805b9b17e2ffd49c1ada5d4acfa767ed515b1232c301e266c0eb58974627f6149a0e382e4c73a4439021f541f3f2238d31b84dedd9ac5bebfd63709c6d69c6be6fccab96ddeca3dde1679bf44c2360d0c3a7ac014b60474706dc87245b630fcc2110db685eb77dee376157cdf74006b13f24a8790d5380bb41ed46ef77661d817abeaeafc6543c9fc32169bdd9a0b1032397d2818c67d14fc760b505e55cf8d0efe8a2257d752fb433e1bcaa714504f7e683fcdeb46f58ef23e1e432978d6ce68fec33bea272daa83d72823f9bd2a946b7ade35f07fe234a104cae74c325239d93e80454cb192031aaee1b7c246f917e3b5ac10fccb7a0fcbd1455acc26e779b7743120a424ccbd3e1968c91d66ecdb35b7e603888bbd3637d5215aee6efc1a14176094c1ddc7e956af0a6db277eb4b5fa29dc329a538616bd064702ba3c2e7bc1957e1924997b4a652bf92d7ddfadcb37f0403f30b96222c2c35df2b27d0eebc5e095710e66bbb5fb6fb356b2b05d1ef2662164df60aa9b54470ce28ca3064fac4ee3d11a5b593834c52171a452158cc93b968d27efd8530b991f7fb317b3b65b451f201de2aaedcbce4b050d4cf2a278270a7ca166e9557d527b9117601f363b4da609f07d1463700df41eb403bc8df18778c72fa718c972d92ea0112d1ebed9273967a8ce969833d4ca45a3a50c4433b40d3b51d5391fad441d8825ad84f05004ad4d24666d477950a51e3182a68d8cc6e26e68ed47576e010441ef29ab975afbae10a7ca2320943a71a0f1617d77b3a6d46c75da5d580f92bfd3decc6899cad8effa2c27fef23e975e7ba08f5860984bf9c36a305e258675e980baa5ed15b6bc6c0c6dd0e5589cde71f47f7f0c4c5098a53aa15b00cf492010cc8fc4b7dabc787266db0a7a346045a26c916363775701cac5f3c53a0a100240e7e6217e3776ebe4c9f6239e84d367fc84f710053a857eab4b6baaeff32ff75c7505132d01e419bbf259c833b38b080fdf3a4fddfbe504c5e615cefee91ea26f2f891fb9b47751e5e8dde2aa71967342586b13117494a8c4a91e16c8a97ebee788480d53876c3144c81fec274673b065459c167d93c769045a705b3dd5c862d7c2b6cb9953f58c39a7854bb96970e446b3b25b71cd2e628cb47db3bd6ab9f442d3f03361a0196e12102ae742034d2ab5ae1729fab87649d84a65fcdaaccf408f8e9b293c1658dad43108ad10a1c2fd4cf77e9cfee27b01fcdd1ce1cd0a21c98c8d1b4cc13ea11b32095b97f1ac5193c39167699099621241c436cace0c074521469f37a23f5a3d0643dfbe4460ab8aa5fbd41c593bff05e08b6b103efea073927316692eb9a48e570a3504e9edad5908ac9fd0040603aca313a76d7150ead0a6664729a42b0155f91b74a9f62de86791a7427465509b512b3dc1ce0eb1f48239ff5db404895027f95a973eee4f021bd5fc5fda255cedff9a676ac34fdaec1f224196277d1e6a6fb33429e6fe0991cbb086da988232944f8e7d0ea50badc41d4aa7d7bda89f9b4763fe7c68e8b6003d53b7f2838971544996961a05eb1ad1f176da89d7222c7a402fc80a765739d5df301348fbb714e0317749950fafd5b5d7c957b5ab2ce0bd4202948c17226f6eb07d3bd625d11bd71fec48c4bd1617622f98c913363f728ff95c557939e839e9f29da00802350282e633b3dcc70ba350d136cb5e273508c1b702bbd359cefedea60713f3cca957ac3e22c322ea3183c14add87e1915fe84fe55ae5355556e5121c5d75350565d7e774643a21fc4ca7d3d92000abf842ce22fa2b9e2972957a3b40a1cb94eaf95331363c19a0c32b926424aea66e7a3a4dc72579edf808f2df6e31b4376a8b88369bf44ced9d42b54a842ef1dd462c7dece34745de8671b052d108204be75181d98b951e6495a44b63a9f097b0d25cd2ea72a6577cd0ded78cf675f2e9e2d0d3b1878e220d39fe3f8093f70800606788e714b179fb8a77eeee417ab1440fb4c25957333bee80c86e23182458824688a4fa9a92e5417c391bc01adbb4f852e210c88c517b1446578af22131b01081f9792c32f34232ffd762d4f214ab7d428fead0b4cb016fba4d5aa57f2e2c9ad6170ac6f635f25d44c123b574987808df70bdedfb018bbc45b06d2dc2154cfe7d07d4d056cdeab363301c78e7e178ef541636f7c6da56256cacc2d7975002de4593295ec52cafad20605f0aea461d8553b6fa790249c97e2b0e99e9a38802d2758912ead9a8e39f2615fda9e710f0403b91fe944ed8b6eaab0a89f02ec54d2bdaf3f49c668da1a031f63975d2cc66bbe4ec23f4b3c6c3232181456567297fddc2442ea21a826d73106de92be3dbbebcc429153414a8a15982dd0f3b84a3467ad6a0bc5e4f8921f013d12e30cf0d3a7a6f2d6cbffef6b0e314647c07b9d6d77ef03a4f23a072a1abc798c142e792d744b2a2f0208af5dab42fbe74f37e06dc334dd21e7c158db65873f63d0573f72c61618a53b4f937954cc47daf991c473c134a060b85f63e3c81453fbaf216eabe1909866c59256611179b7a1c0bd7ab9245466fe6888263aad71351ad9d3f07a16fd6fac36a5be3ab4ce2110272277cab4d711c98fe3c5760d7bd2b4047b4f7cd5bc3c6631e98c2858a9c52b02811544a3e0727441b0933686663fc92afb61fabbd53de559decbb6b487e498eaf686ec0de31b68336b4d89591a41eb574b5de6150aacc06babaa1aa979dfaf7a9ab62908877ee3836ae378a9efad435400800f003e101de2d9f3c623cf56463e08a4b29453fe7d0ddca29464b8e365d371c76c53c98f0067ce68af5dc641c27ae520a5a0bc2aa80887d6880e7cd5098a9785aec7bf3a89c2e066c26d62ea1f955aa62dcb25c65a91d94161f798d214ff6ec3e1d5d60d16aed39bbb9a9d61d9d6b0760f2ec3b21b6f1b6e0828d4e6935a9c953b18855b94a665698bbeae5d92a00f872aac6c61cc16201c957d928d114dbc2971694859bb1df069ff9d7123ba897e414bc962850173f00c9f6e96246999edf1b0aa0f80332dd427c66aa81c760054a314c74eebf89b8a0b4e1cae14438e94d9a26d3fdaa1f96b03449a3044b53ec7293358c6312c740305cba5b81b92c664c7d5e6e0ea4210f46964114d9b8b284456b246f495389cdad7fb64289c3616a3cfc2aa9727c560233434ddf60d4d28614e3ecdc74ea0aad844c3aae5512dd1380701303bc9aa63a29dc693719d504bd323028997c106e5f43aaa2e04c3f7131cf7fbb7b6e7768e8d2823d433b39e1697823d3eab2f3e79b67546cd2d71f7639f244b5495611adb3904df0382e064876ab98b22e244d3828b3f8e0efa466cb626d5c193d0db08d98723d93855e2814ba3c23f820d0a97b96d68de74231acb0486da1b63a5030e92b1cf3371489d6307e18972f4e8c174ea4f8e1ffb9bcd323661f6a69b55fbad1f4709058d219eb6bf7004b8a87d7e530ade5e2d3ce77563ea2476cbe5c89a107f9924a9de8c0193bb9fe45e266fd561950553d9c086d7369d82a72f03b513ce27015808826ac0f5c54902a75838694d506a61c682c84325bf9079e32c820251e5a4a6f7fdabba3103835ac8844f51c6a7a255d5ef81b90b13ae39decf3c3e0ebea3738667fa7de62dfb9d082336a2d364944a674fc61b88241d2bef152d5a26e52f2373a6738e324917efd977a87c78e2453c63dc6161e86b9b810d84d68440f65509cdad5c3579b9c97a87c8dadedd9feed106cd8e9eb18d66182dcedf9d5e7fbed1962e30140549c19fc0a0517fbde5735b13d9e2335522e93f4cd475aca817befb07536a38394e71fe01b98ddd4df6e21e1620f20d4cc84d6216d15d3821855904fc9b8f4b4c9aafea90c9748b18c3d82386e91;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hdb3029c728397f7b8cd5f09799aa50f58018546c4e18c33c092ba7d91d0a91012dcffaef1f929a55a60da7c6f2a4384476ffcb3bd3b3188ddd0cae18b1de05349d4a7d66f463f2582a1dabcc3b3b72e5aba97f111115198fd990a1a1955a3b4598b4e21969c3c593b92007ebf1d636d4ae033c6188c79f239aa9509c0a52b72d0552305c150777cfd3b6bafc2a297acecb5add801d6d4c74edd334f27261760ab4208a5c15df89e3d903f0e45493241f7e5a0000132fd08b99a17148ed609d2f8fc9dfc9997d835e513a06836009cdb1c293c6b6bd96f4ac1182a529005ed675515b1d50af6b9e08369cccec8390a9fea3bacec8f53074371ec8c059a91b828ace87dc3859535faa592c77c83f835af12e6ba5eea008795711ec77acbc8ee94db63d306d928b42dcf185148f9bdd93e135a2971d6e52f05e35d2e6f090b2be4ee781fdb30ba00274553606f3626a9b3d7bd595b0aae9a9522956758b3301e14cabdb90fd2fc81c235ba11867dee136ea708c778b3f274e15ef49546f352433afe67084042b4290ae61ec0f98a6bb5dc067cf2732a95c76314e74b41f856e8efe49f91f2a6c605da668d988f9623950246522fa822f80f2b094d21c8ffd2b2e4c5f82636416f11d3e4490e9b81fa3abae7113bff263172c69311ce0a9540f23ad86107caccf29290f7607da93c9013cabd754dc3615c040c8cfaf6d8e2ccddcae1b17ba98cf09f5e7c1448cb5d7bcde32929a32378b176aa04ce3fa0e0ef388e25b545f90653be8f809d4e6dbe1ead5b6f00c358986d97d1cdfee05f02956ac5deeed87bcc79c3f5fc1e884601634df3f2a5449f704d4cca43d53198aa35cf76772ddab3b08f7f924a91648e56229043772d5fc49a9693e9ab9eee6c2be95da7bedd790b53be1621555d7752d852e427e34bb796b34866700e2ef75fe99d6241887cb21b58d2d27bd76644fd3a07a5f5f719338138ce38fe2d039d1058c002eb9ae9758d632cbde96119bda40068ad6679a5545263bf89bb3125f4ba01731196ac899ad6488c14e346a3f1bb1bb6a6a89bcf412a9105de43b67ec870f3970401a23b4efd0a0069a35aaa55564223c39c3e1cd3a9aac6e6d8b5f7cd423c23508469b5b9f85cc7cdf74fa84c3ba2ffafcc212f69aec557e9ea78d3ae1487c56bc7bb1f15c2f7dce8844d040f31baf92d6c42093b32bbe5a2363ac99fb08ac68ec7a1ece9e26a36e761f80fec4369923caceb72057b390afee2724a6ffa79d0024bca5db182d26bf428b7fdaa18f149586b600c65a50ccdd82d648ece2e83e35c8c014c545886ecb88330084f6c0728261bc07fb69b18e3c4d49e33b3adfae7159fbdef4ef794a16ef4f5f7cc274189f1bbf5281235b43b8954b75adefc0f8c1517028f865abd04da6c881732e2414a97861ad294c5f187083b92a39c7d1a1f5096e9071c2bc7d047c2186a01f342f04604078e3a5c727adb36853f624d4c7c2d05767b63f4acf95dad70cd047289eb4b0c8e2f41606679561bba0505e04492e784f8958bdedf65ba67ae582514c918be9c521c01f52f05de9b264542a5713266881c58130268a6f433fbedbe6ae2a39147549b5c9aa577b6a37d7f81cc7b1cba8851cc93646f7339aa59f5bb1769dfb9db6fcf4502459fe0ebe2ef3ded563e5d4abaa9623f925364bc4fa09867eb2b56afb5877bf895909fd904b89b944b76b83a631b9c8ae7b27ed007096b8fa68f09ca2fbcdb490746db6455a01e003c2234f87787faa0771bd7e86a75c1594b6c9ff083a9d237c5e12d36d8f0a6f0b2b6caa980d70dd3e0f51471b025ffb27f2d438380e6cf386796f2b62a7e2e9f83a7b4aa95f14bd6547dda774710b967cd6b7969ac5cacf91f33011875bab1d9195f69a3daa20ec00e56ef6792bba534eea8cf5b6df9e4dec386eceb6ad5475b48f8c231395fc780d55a5c1b4ee5df5dfcc932c20f2dc4d4e89d3e3758863b828530fee568042c9a3e5247c6038c5be9dbcbf6ec798fe3e23239b68235b9c73e58f1c9800ea62586a7d03db7b01e19b5bff310e66191fd2af6c80f390270efd043d7485ea7e73c607122af6783b4463272bad0c6ff4aeb091ef18502de950c0a1e7fd8360d882f6ef880f603c51d4589adf6c4fa88ee5d2a8bc73ce96604b204616bb43bfd2907e3b22e2e28bb260f7dd07dac44849a173433db098057fd265b0e92e53ccb8d3b2a4756c7c1c040195dd8f532eb941c7ea077dc0419f2be2db9b3ac3807fbcb2d031fcb2f321beb39555fed03e6c156a2f38ce0aa84e941ddf8dc9fae8b8e1cde2f4e43ddffcd28a9f72249d95b79664e5fa55896c0f13ef2b3d795c4fd656e13b98d0c14de6ef8d86fda24bf93ac6d8175e3b8ffeaff87d112b644ea294b054e1c2d56a94de47ddd0b3341e944ec336632e33405d54793bf8c949c0ba0841f4644389a3323e9f3e361c18fdbf67b97b2c16f475415a610148db132c8a8c0ba3fcfeb4fcef6bac89615d0cb9ca5a466ff9ac4491736ab6f94a2183e6d138350b19b8411b50fe748b0e666e620816c471cce2afc6f72730debac8bbd0c811b815a0c97ca89aa8db9ca392c3ebae0f545fbf69872c0d0fca0f4eaceac56ef8367774c48a48d26357e2e5f0e563b794f86f4738bacdd7bcd8cdfbe1f912404d044bcb6ab64c6c5809f373183b154c7be5156ef9d78411419ea011168a23f3064cbd0b8dc399901bcdd872406049801e80334bada1723869f6b830201cb6dfef35868fc4bf62c9b22b98f20010da323c7ee00ab54a0fc8de125c61b36261cf66462bddf7c9164ac2762f1ee8d25834f29f51b9f1117633dfac48eefb3822ed090170611918b1e11b6856386c08668edffb30c449a23268071597334b96966eaad630d0858818825a1a841ef2cb4eeb9d45b2270a2215fba727db836657bef63269ee728f1152ed4451a1b1198bde7e613d9fbf1b1c6d1289e07a40ac34eed8a5a57e4effc957b317fb49598c2f57723665459de2dd1c07ec21da9b04f46fe73002acacce833dcbe8b359e5788f0530845b6083644c36bf6ac5e93194c7df9f61bddb8438c53e7bd3b47571a07330dd4e16cbfb9037d5301f42ae764ca97eba4122c73e119aaeb34cee629daa5b01c9ba4215aa73db3e8c2e75b067d692d08d1adf9a1dc0a08a60af938ff57f35261c0b51a8a60525145cdff08a7aac72515c2551b90dbf4c94deaf6b67e33d84d40098aa871d32fd5c67b402984685c9a88721c764bfedcf07869488a3f1147d2bd0a3b762b6b4729bd05b11b1712455e1fec0e864bf8d649f17d375282dbd7aba86908e61f9ddc835f5f0c68154cccae6c74a1de28354e42e4e77315a4b9da2c7a007266f1fd149724f6b4bee79590cf6c13e3901165a9d05ffb1f1403e067967fc9f3278f63d461dff0f49aa085ceca47fdc8710a633a0b9362476e609b5b4aa252731cbf6949c0318ea7eef81e4de47c91d6a62bef1e9cc2866f46b70c3de77f3fdc27d8c77f4457a5c40ebf569cca4f10a58da581ec35554408462069302a9c5e4438ed077dee6499d543e764bdfdfaef742e901c7fa369f98ecc1ad5a36ab27ed877be9942677b2ac2b6d1b8ac60575ca7a7bd4699fc7e73ef779a0de336e42ad05343ef3970756eed22b9ccee032d2e15650f56b6760204673d569884a3deef94a2e176e591c6eeb5d35a007ee60878a19ee060bb0e7b40e16226cd3b70322b01a8e55b3a24e366991bf90600198d1858ee9cc6584e0c55eab1c0f91b17936699e30cbfb914a1658565f52a06ce8e002873e859a6f609e1b250fb5a1b325427dc0f18e221817ee5e47e7361ee65c6fec255844fdb9f9f1bbc923d10e2d429ff28d5c5849119447e0f2f82866788b069367a83724bc61fc0e281a11e51e2ee146c5476bd1708a241f75df11c1df0030a8d4e3406d7de2c213d8ecbb5b5c3af69d31ac58fe6e36e296501733ed3f89a0eaea05547f3770ff8ec355990fe670f81b51bfe89c67e7f305349286a9bc84cfc29063399eadd2beab27abeacf1a0ffad414b580d04d4237b4c6b1e981d90eb67a2b495e86519fe8c0127e6550cafd56c1bd00635e4282b3a2ec306bbb5d2ba88c8fa98ad1ca50ae0e7b43abe032155c8255dfd1d45f81e3d269974a3ad0ad52093fc5a07189ab801b5bbab3b3fbfa596109a80bd6bf278fbcab705a03345aa14ed8c6d8c810c9f807114f76643a43396fee088b06e81a441f4a530e647352b52cdc3732fe9ccc5de3156c2077b89c4519c80874ad8d38f054cc1f89eed093cd6855c5665fc1a2325456e1cf3cd87d89e4bbc195131715fd37cb9c3c89bd943a70c7805676eb92979433ddec6a0caf89501341277ff62cf549343893a3775e9a3a08cf7db18c726c5b24db4a7666d25efca1784f6171d1b073910062f77670bbe1a93190d30dcc3f028fdf8306618b82f58ff89c8f01705ad9c64ccfe09c3a175ac5562f46b5dc153db4e020ee52cdf9c378c7992df7830eff54b458be3cd7a27053c6c56e55cf17b4cdd4a26afeffbc5576c72bb72a42fa0bb31130289d5af273ffbd84a00cce20145aaad00147533bed8721b5d0427dfc5ab220f1aa9e4a5bb811e5f5400cc11d32037d273c959e5e295740a34d38b7d1ce3ec8943e704325b6ca0aa6003a842f8cb7eb561e4a33b4cdf69463bb9063d039546d49611bc71f66f5468fbcf9b063e7b13a2f2bdaf177be73419a16a49477d1c719b0f89b7ee61dd2a52ace66aeb5b733dee0d602d3adc0900f6befdd4d693fa04ab162b6655aa13840da36a561a415db59571dae49d29abf38f8153c2c3428da4eaa629ce2b0b3e4315260718109ab95989481435a6adaeaab6d87a1c72d3033b9e330c036949ced7b5b0d2c56f2dc1babec7e39746fb9a0c98d9b3ef309fdd4c74a6acf30c29a01376902ec35d52f13d2e29f770808e7535dadd91e667edd9faa46213caf39e1f9ee6e78ebbb2daffc8278bfade1379032933d7a2cbf64288674d29ed8543e4f38014dff5c8c89b261713d5fd86c6682b4dbe6f1db4a387dba577c48836c2776f8cc7ca1101572cb57984ffb6873515ab598c734260f5069126429fb50db8fb7113f938c17b66659d55b566ecd1bda575770a38e5141e79a257cf304ad61c12c157acf539f5d0d41c68b6a019a81ff2818273470a2eaa948853a5008397d0cd8a854ddece7e309a5dcaaaae2c7bfa069f01e35f0e5cc8c3a95a0f63f4cdca9e32ffe9f0b6b0142a9e8eb9af12508e1530d08b6b5eacbc268f2f613ecaceadf9308a85e126e851b6856e68202b0be80a6c3c3afadfaace38060591beaa233945fa79935bd6ae8af9c612dd50da73109d917cc1bc1650ed18dcb9377ee5ee7451ec504d8abe02361a5f574e4545eec70213b6b8a133ef719c3617d7e75414775c53bd35e7d3cb14ecabd6444fd83578cb2caa3f85018b8a8ebf4a7df013deaadc4f59cd269342e684e4894036b91487c25f4fa1254c68bedfab7e457abd2f8228bd6be2bb7ccaf791b0edfa9e46f1f5c8ff81b25a438c348cf5c3931eff52a634071793930e245383e28266185cdfb89da241b2bac2d78543b3855ecedcfe438a38f0431a2586b550ace47a8ce5c28b1f99f65d2a925bdaff716305e0d2e76c60e85c3c8c9cd619417617c1dd537a7862195c9731aa0de3e0a15d15bdca7363e683f651ce17e9a9eebc95d878694fc5a62172300dbeecc3a11be575e3a9d586637d8a9a6f5b4891a02baf8a750cdc1f1c9f1513dc98d09ba2f58c4672b8ad48592;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'haa2edbcf8e420fb59d2f1aa9ea30cb89e45e18c615875c39bfaa9ec4ade56e764fc09463e8bbddd986b284e1878090a1f65aae4991d32c5350cf8b61d9fe9ea4d58766de314bc400c921dabd237802e7738f4e76f7b768a4889652d5dbec1670c2fa64aa8d4fa6b386e200d2293ab5ffe18211ea80f6500519650fea68f8bd1d731067d9f672b4f97a912c420321e10c9ca29f4c0a03ee9217f02b670ad695f167c72560f4db18fb4129fbc3184b709594456329c5adf002e59df03b071b8d0c8fff669ede6a2bb30de720e79542be4e3e4639b3bc7ad9fd155fafa7eb210a221d05e6a2f8b7d9b91f42189a82c8678bdb4467bd47198add445b43eb26943f9c4ea96daa106002d2f593983e356aba85c8a37dd7fbf64b227b8ef09cdf54449461e074b388e3d6dcbd04dc4e3968c842523fc84402bdb343794ac4802e8c649204f774e4ea399a7c81a1d127fd3738242fa387f621e9e77e7a00231e73603da667eeb962e3dafabef0c7e951944633f5363c3c97c9b8c50f74ccdab07bc3b621bad83cf614aee836e4d226f69aae2d2f2f137c9cebc20eaf9690862b8c1c802d0ad2888d99d1a110c3a04f6627cc9c2eb40d2e3e8b42495197e3876f3988b20d38f5fe0c739393ce04797a29b4866cb4aa79af53fecf3cd94a930c6fdac7b46955e8241fb19a22fea882b741e211d6a22bde4e7fb6ccd657316943f26ae9236b03f0558b4df4b610db970c4e64c26b5574a5cb8d8438ecabff6db3ec5344d55e4ca9b1134f0b397f9fa4b507718d29ff1546ed821cd80060926a2b7749c413791f5e6524de38691d055c31f426d5628b05189163eab1a2b0c9d2483001f63f56d12e632c09df5fdf658997abf544c2930d5b71831aa4c499014253f3dc3d15d2e0053afc43c1e2c24ce98ecea13fd743076aa09cf482fffe56f43030c169c0d523960a159bfd9c87bf23377698595cc3d490bf1de08a2d97cd3af3ddb4fd8616cb20520bf55919dee01e5d077b1b959fa29f8c6ebf84637471a312b235b49f66007cb837d48dbfb3b1b7101dbad4531455ea438cd543cf3bfd7e83571954b36f1250f680ede182b6b200c85e1fc034a7b0944e8344132dce0f2e5751a2bf5e58e46fd8221e0d3f01d2e4128897b0e77caacb6c4023be0c717962b1ef3d10129d9c602ef532208b323766ebb3eeaf6c1dbbfb171b8912ca5789242a013c7b9fa2bcd80626978aebbd95050d54649994b6edac73d9c28d6ba5ec62c4013d357fa505e5c2913fb59b3dafb3237213a5bf997f8934a748b387a92877423c1cc1d81dde325936b467cfa43e992585a84a16543a58ae6818478fe7e53cc11f64a0bb89803247fdc37ad24caa149973eb797f7829f1f6357515b78d39c0ea7c2d215552ae305b53128c231b124dbe26a1fe5cc623bb3e577a2eb64e051b3bc80f120dde2f2098a5db3311193788991dfe52cdeed84d1deadbc499fca478c1b741660d0c727eb0e6cb0e989867a1542373e7e95187beebd172bbc46450d0cee683acaf9d2a4f73580ba4317daf666f9c49e13abcc146cf0782997f49e5a982d5bf9d9f74c509c5714135b440706b1d0d2fc01caa48166a04cfffb7e084c803c5f74e9eb89d3270d2dd07ee0398e57d3c5b3de8c849b50a2589c8a05baee5981202391662c0f195e806e792903a9a1b87ec2eea71b3fa0fb1710df9b2e1f244984fc80f83806bb3ff2201b53452b14a9c7f6a8417bced57af38a36ed05e9cb56d9192b9a231d111368bbb9a3898aa40e9dca3f11abee6ac4d769a53266a3c759828ce3b1d44e6e6a066d4362e7ff9024cc29055550e6100153121c4132bdb0aff57756d3c742197444a85eb0099dfd1ce58ec12ba810e87b330dbaca8dd233c213bacf3efa1f963de3a28a596e6185724a6d81db3b52df7287802f0862c211cfdf339cc776a3769bf516908968f8b28d93294722d51ec9df4ffc90c935c46f5588ea34ec3b1611324734376cb1cf03763230af1415ffb4d2191529043cd3b768aae651a00f17a4129d0dcb79abe891ec9c9c6c5bfb9c9a524f80224bcf9f2cd5d4defe1e9673c0450cb454906dd3de1ce7fbd26eb1a4de9cfc93c21e0c08a983627e34b9a7b3e4436b37682d448879e132e7f394c251870faa58ce796ed52c503092d4bb486b1f8372b2897d40e82ba94475d209b83808cd240b16ea17697441039a7f5f9c35e4e847d90e491cb60e714543d4026d8422513d677b25e6f5a09c14dc58cc3e4f463b74d330601226db06a5e0ef3686a78de7689361b51ae5c6bd53d7f9d682264e57fb14e8f57b0c3e96d7d90576ef2017fd0e74ab2c1f6bda9849d96e47f5d6e3da9ebca52f6abf18fe4b071f6d3210515b6824209760effcd5de9717547838de5617e1695bc9cf5766aa71842dd023a78998f1af36fd77fd5aa79bb7fbd627c5566e6b9f2bed41771c9fa33ae8ee7a071d26d9f7d319e3bc3b1e346cb7622b780a972c1e8671f8d5fca643dd68092e8a2f8241a76ffc4f2e4cf3e199565fa1482e5ff238493dbe63605d5a69dd20507cd948e8fab90ab4e32f00e1389e67ceeee8bc88b0c516a19f37a245426171b024063d07a3d4d919b8000da7b7599ce15fcdfe87897fcdc599aed87798128ec2062f959d4ea3082c23df7d597303e9642c495c9e681dc356334f6ddad19c51bf66722bc48d40e76f17da8bc95974f94d31f8e807f066bfb547f6415d920995cc140f1b31fcae5a80afffb9f3a1edc037dad146f9c16c217c5e54d92734429e1e7d6c63be7212ba3fca00a04787cb05b9fca8a052fab0c6bdd6b2e18b18fa68f2400c132ad1da644115396fc91e66d04d97784d0aacbfa04abca174ae0f0fd7252ca806e9af460e6adf7e5da6b073a603bd2fbad7f397e6dc95277f7615785c088fca571de93323738385dafd1beb47d3a03ed24627f370cd8ab9eca5ce2e0417e1e3f50bb7024a5ccc3a8f99a3ef868d2982f0f1bcb2491a3292141c90ea1e28931e55e65ca299fa66ac484886b390b444e489a8aca1ffdbd0ea3125b8185e7e7a6c00453983617374c834968ed926e52455e145b671070ec34b9d11883ba9cc1d71d3b1174a7ed144c56c0c800900c9ee19cb96c870ecbdd4f5829e9182d1913ff2cacd5a27173d58debb98a83e2c61e5d2414812f1c0627b5d07dd85ad50a3e85584cab50ddb29dd6e4a4bd27fb45fc50d139eb70e025d2aa381e5092960157af7b8179a86d8a83f82adcd66e358d01f3b0b2da02855746e74ed3f3fd8aa5a5bbe4ce9d5a857bc4bbe672871d40b386f02b1b3c19af423f99ec5463a0dffb76f9746eff9f3704e86e5be553dfe033f3aa27ea4dd5b3a09f7d77a14e9309e84b37388a06981e296b5085cbed1179d950a67a60065330792bea3714fadebb7aaa3faba125b70c35bd9b3664dcf8024515a7422ffd852e118d6ab44698d4c45a79c3e5bc13a6f4a9ccd1eccc691874bfcebb471531246a477cd2d12f0d304120bb5fcc8cfec577212b21edde069368c2253ddb4a6cc2c735af5f23a2e04e534b1c9f8229afdddf8480d778595253ed4e1e14143d006db725a80ac91e3d7c604da41ec5dca96fb93b4891092b34bfff4039802b9c43797973d5719f1c9615baff68e6f6a4cbac30a7fa449168e472e20115bf767257244a1a89b7dc9544fa7199fa52c7859a1f2bee2be7a0df57c69a3153d1ed78d62df0013efb95f77dc6bdb6832565d7a9fceb40c6cdbd4ccd38416c9ad4529e61e18cf624d7300b3ab9c02a00bad723b8566d50d2edb8867fb8c65b10482966bf735eea365a4e02d45f4599e6f3d92efb0cd6262813f17033c8ff5ed7399f52fbf31445dd73f82b000edd39c396fb317720a2d13db52444bb92a1c94bee4598b7f8d898ad3d5142b6318baa66621dee13f0ba6da8b7aaabce03034c0ef4c7c258e7ebc509bcbad7566db24b50dbc61407cade873da1def44ff13bb45c9c496397088b45e1793e0d2ef87abb538858686f580afdabea82fa30d85bdc740c65574ca181635698331ca635c4de17ad66a04de0235124fe1de2c385c1544c3ba1b298f9874bd16ffdd20412724bc69e458a64bcc593f7fdc8ee259ef97629af30f354f167a66cc7614abb575d3e96eee75d580fc12dbde7f531e8d780dbe455eacb6328ba860aedc380b4bac5b32bf7e8f636ba8381fc33aa6ec78e78857bbcf189f37efd3c74fc4260ff4b6b6a030b3185553a200a7c9b838d818a0954ce3bc57c34d9e742565ed7558e010a91f79758999fc0400cfb02f63cafb457ee3b13d9444f53361f80d08944c2e4b2671465570683b0c7b29ce9a6fd44fbbf3cb244a1184b2b19e2f194e81d756052a6cfcdf821760a55e1e8a4da9dc65c98f64d0629adf1f01734bc1f059bc27aa4225377505aaad1c33ea3517a7ca72a58b771f2cf5aba4ace250e1ea30d7f07e05511655e6ec1df40f613d7115cdee185cf26f9ad82d684dd20741b99a4976a206b915c08f8ee2c94fd2cc0fb0ea2406ab5c4eea2cc08933a62e6761de4eaaec6fa638f7ec956d0fab6b8d183c40c9054a5497ad2710d9104d64a0f9566f1da6485d799c63186cf6a5918148368ac109dff86ad80cc3af2ec9bdbec1d32850d49bfa6f66af7f7a33abee0c0f8a4bd1feabf19dcffef322d6e8c7e07d5cce3bfe86ce109e5bde7a624093942777a8e25ef65f265ee1eef3fc35f621a581179d2da99a875c54d31f172cd8ad05b9731f3f2ecff5116977662059ce3176c7afb6b9d51a2dbb7ae94e121dc86c7886e641e3f09a433e2ecf513673b759b7ba020aad4074e7838d49e8b02ffb360dc1ad03dc450a14695f6f60bdce6a329e8c3ab8e9964ac3c73c5694bacf74f1af5ccf65da123e0feac40e1df4dee418841cbafd2cfcf32ed56fc33da4dda572a6f1c192976db325902f9d69427b9314d05359b43c0ab25f5b673c2df0449b1c5a885c5cef43f84ffc93e25d0200ff12c68982068de5370d350d306144bbaefbc6929e438f296864c695e704a2f7dce3cc959f9e95efdce153d9e1ed7ad6e19cdd891ea666a7b4ca7eb28cee8221e75e2223db3bbc0e22cb3310adc61692df535320f233e373972736e38178226819b824ea52a9b08346519de8f5c907b9796f82a42102883869a4bade123d04999bc4254e636480fb408f905d85b3d9f2000579b235ba302daebc5a9064b2bd70f933634b6d75885fdd41aa1c552384b057d783c264321fc92005df47f0efb51bd8d6222ecc3363d2e8dd1f369aa75055225461c11d5e5565f42330ea6a0d4f835616ba0ff24ff30089e6832bf5aa475644882cb677c78942e6d06768393ddd4025ac7d367ecd424305eb9d784132bbcb24a6c8fccf8fb1b89b06a7fdeecb3c0ee0e682fdbff310caca4694053f487579e8a6c99fe63c30c616169dd18828d0b282ab79598e7bc57f332290e6c8d416f96f19045c55caea5775f9813b7f923eedcfe1ea90beba865ef968e55ded4b6d34238bcf4561ff312fe083f3c7db1378569c833dbc351df3a65b3f2c5ffa949b12f8b801605844312d5f7dee7170b0d04abd330aafca5657fc915a90a7e5dc5079130ca5aac01278a7af48ac60a0cc0bf8202bc366eec3b9586be443fad1e2f1eee3bcc31f195461c19067342a8619ce5f4affebe11f25ffc954026b4512c77c6339f092515ca45010fc5112894f5e727db5693e194db730f3ff4019cf4aedf0dab7fa2f0d9958fd45ee1dc17531cf34e11a114677354fa9326250dab87140d403d680d3c749c84e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf47f946b6758e3f8a1e86ba19ef7dab0548747341095eb84479762c038bdf0cae7354a0f0c63ae6007093334e222f68b011996cf625f1c31b6da1a8ef639a0b815e0111d18f3d16a771cd42308e13075cb5d54a4333ecc69e0c1accf8d0f63f6c2ecad07e267301c14cd3638c16cbfe9306b266b117ea93077ddd6d9e5025197874f1e88278889a3f31ce0675bf648b76187f8ecfee1f0a3c0536f5e199e9256710fba13aff8355d0bce2b5f99d73bce37cd971464b11888281a83e1f2af65d5ea8df7f048ce4cd5099deec9a9dc3c3ccf0a892dc06f1dac2fe5fa3aecc26b36b9a7afa2576b403f550f7ed0760fc62ef7f8e035766c58ec5b008f04831083acdc9bb28ed550a829c4efd39f07fa88d45ff1ad3b9fbdaa7800238d518670e198c4633b9f723493962a59afb7df1bda3ca721392aee44c71ca3e1a8a2b4cb8fc38585449a5ec455d5a9545a09980842c71570216dd5b28a7528f0d84d540c7e862d1a8887b16468b82e9cf567bfdea32e406c87c299a8904524e0381e6e69dd346a3979044e40431c0fa7f60dd426d5bfda0eb899d993e1c39d8352045fe2326ea78aa7222c34a5b7eccab059aacbb0d6ce6792b7bf0830065116adb5e0c74169c7255d1b83ae71bee424ea40d3aca97222bcc4e41b9a047788b0249fe0b162de66ef191ad3f898ad87244db91e8e80e4d699266af046d25cc69076b6af74ec9e1cff9c79430e56d7ed0f9f384a3fbf29223e06ce2ea156898c176c82b51d0460f60b6b68fd340a412fa4354dac81c991612256087270e14a1316974ad1df4652bf714e5c697436d22d3fa242a9200688c2be5381e95804887e42dd1cb0066e02f83721d21dddc5c813f18c489d955a079c59806a3ea64f104786ed420b48f8f98bbe8ab07b606a7abb781f83a3b9ba53a56af8f598ad94ad26b3d0c40881d3eeea8538b07bb9d91feabec209b4d67d9f013ad7f485fc39adba414e9ce32a934004da44687abdd63cc92decb829c04faab1bc1d54604908c8665ebfb68ecfa78a0e761b14d057fb4824d6895716b559623f804cc70e9fad23d6e5f6eb0bed5710a4687842de51347e3003faf7c4bc323673206fc906804b6145e1ae8d72e5a41085b9707a808f719ecc1464fe8acd9bbc9496cb7dba68f0355f4820520c930c29fc99d834aee6907f5fe0fc426ebfbf8f751b1d98f349ea7e18e31a6957db4a30da9c597e67b710a4a38a079ab598c09b88e4ec82caecc2e64c9c06c0d1c1456894ed40133c04952344c18873f063aa6d3c39882caaaa04e8f2a36340c5fa9d7bf5dba516bf1b7c7b4fe18505a0f9b167cb45f39457dc464f8e8f9cdb961de9a4700c3b7835390f1aa007d58f6e49e563d9054c1dc21766018999282a151ce4c43a0b5c9a9b4133ddc2f3ab416c682bd091dc58cebe198bc01d7f13c0b4632d351fbbc27b67818aeb70ed212118bec80d7967b640e11f982b1b8b383785e3511824bb3dcf37c5332fc8cf8b0e773b680ea19b181f4a677c8a2347677116fac2096997d3a9489c2d9fc65936872a8fe95515c525d00debd411054fb23de7c7b781c66f1d61586521085f68c79c42befb60f9e7418a1ed1720e6d542f3f9f0d64bf6dc4e887d1fe1cec28629eb266b112b59cde22e7a23f61b872597ac932fa0793217986dc9515bb409d323b997d256bcc640f396f37875dccdd619a0bb163d8fa0bf2c7407f56119b246a7ba924e1e322f56bb200d5b02608c1518e3f7bb73dd5e706ab6f2350dfea5dfad452fa8d595eafd2fdcae10ee8d31800bb208ea35ebe5a7e61a8d35bfa13b9ded62d4f415bb722911fef38fe45db68e908a96211e4495b3dc68c835b5cca5f15bf7458196b1dd80d935bdf541dfc8bed837392e34df335ab614cbf628395d724286fa3cb6fc8008fd508330c48329d6840e4576a2156aaede063c63db03b709419f0679b4f9865b4e6720ebd1226c6c3ff02367a9da663f7ea9bcbf53b26e3963b496dc0777b19ac1cc65776a81b48fa2adf6c65a78d184bb5e0d08f365de0fcf247a5e76536d450460d65924e1e883ca68f9ed144fff15d5b5af9fcc2b9333b89f8912068c6cf0b7688ebb72194057eed189f7dc6b22daf0b971d81bb865af73488f67e479dfbce2cc7266fe0da42579ba9b49db52f76dc3b03867bcbe3778ad3d9d2f5056c8d7581f3946748aadad54ae5b1d0a58e0629227f49c905697e92c1d89fe50e7b7060e443a35789357d5a5371c132826e879b84102cbc94cf536d875a8e4662a9f60a15c5bf0282b0ae9832db26c95eb2cddd5ea6dbb9eb920362b3d27267a8c1685ca911555fdb78f5c3c9441fbd8e77eda13cb26d4cc403b4ca5b5b7afe1007c1372453632b34a777bc35ed7080efc4f1fb826542029d2a21f88064ffc60488ca8ed73e8136ee2cffea193456342e677ac99e7129285f7d4a9b19403f97b546ad280a428f4593ddf0fd183a24a6515e3613973b305c3badc1157e61518a36c19cf13b3a0a543143ca5a1ddb34aaabdd1656134c996c7837ec78becbe4cae93d57ab563fcad31f845fe727e1eadc73d21f645695358214deef2a414664c3f7b6e90d2a17631e2cd3d590b6aec9f6d7c9678992527e760930f85649f72549d215b0cf541a6b766cd4970b8b3ef75e4c716226b9e5f799d477b64e640dc9b9139812d6d46ab6a55c830511b74aa53d432da1554075413940ebf89ac45d049640c76996d5a108803130baa1344f6c70d4fe36f18b7ed13c551ab6ca53a37ed836b241e72a495e118a6b246a4a042aebfa5a79ca3d061b6f29ba6a57bc8db42ee419243a7c83b123de5d864aceba7a04ae37e7673b074d020f104170beb287ba5d68880bc3144b2daa51763ad07a52303642ef43eb0ef7840384ae2411ccb7786acce621a93709c5ea70a0cf8fbcc0d5bd31af44f5c61ee802932d18dd353024cd9ba4835bd839cfc6c80a9e698a48f72a085f5639e2b87168931a55b39d1df63135d909014648036c4b70de0290d546b2e8064aee16f9e1a480ea3c669a13da34875394e147753aa54305bb163cb7264f3790cbbd8339adc5e293204a6d63d2774b8c3b74ed0e733286f35959b547a0d8812cde297c510d90d7de962430049d090898889d53ed4c45e2c4f31b83a2b0927dbb2afbb99c5f114d3bab9e2115d4ebd2d2d616a11284d9a8eca47cdc002cd2a49b43903c5c2e029ea833d564ac0f723a7f40d442a34c91d0ba6dc0d2ff31810b84593268b7493459e3d237ef92604b3b74a70499b568dc130f0d947d88de9d912a657498013eb47f12ef09b86cc35c6f294561726fc0b2092957339a7185a2f86ad424fa5484e540a20d5dec38b42465b5d08208d87d71a628e76e160968d23dc1aff28baaf858dd5ba97c587ebec1b8c609e7aba5c046ed54818f342d173b1be780bb2813f4e3ac953c273ce80d0152341d309d4763e3d590f07253244d0fa9650823a462f9b0e8cbab9de675568c3392db3f20288f6805df23a4f7527b888f031d91cc103cc6bcde59135c93dfc8567c28b188b7c397d36c63b03b8e67edaf4ea472528784a97d2f0371257de163bead0a3579bc594e5ce0e7225ab02369a10a30310adfb40abffe10ce86ff20a33bc475aee0bcf4bd4bafa5d5f8de2f1fe65e1ec7ff89c6a6794f4cef9a8c8b4c085f035fa6f88f4c7a94f1a4b544a869cb16b20d1c73d94e7d2644d32e56155d5fe12c562d0b1c51ef058a537a7a8e4a11504bf0b50198b41804ce7e84738d95d1b001d4513e50dbb832d138f82ce077f364174519bafb7ba690c3cf7a67306bf2443bb98706075ea4e7f21aee7ba5a973f49d18186793ef2418a6f9b469ca770f2ff567ffc2f8e2030d82ae655866596801767b956ab43d980c044ff8a28ec26499bfd2d73c87128aa001c0a2e9eac47e6891b74ba532a8c604cfcaf30c06e8923b3baebf12cc6b881941e4d448aa0ffbd5b2f6035f438a326ced04e6b8a1caa86c79106374cadcac19417e0220b09bc6a21435281100086153b76d8db786d06c2356f1f67326e39dfe1ab2efeeab6663d98399fdd1702bce068827fb4e6bc6a66108f70b11ac6e1a43deca2bc73eee6a0ec79566605f18931a3099d5d16e268267641c9cea3028770fec308603b0bfbd0c59716b74bee94c6e2b4cc4d0e8e526a93373def97ad043d2cc29fdb7c5b85c70339187a46dc87b39ed8f03aa70be67791fee02b1f59bfc385fecc99d706354292be92bc9d95b1fdb0ddf4d0d5737ff6a2394afb5e8cf09493d0ff117bf72373eeb7183f51234f80cde7e55111cd5511e85691739cb7a72106f793dfa886ebecd5ea1dd9dc6508a7f98fe7af155fb5293d87ab271ec8a2ef527ac363f6a9de1744ed416cd7be2268c48f63c4bac1c82d2bb1226f757a97ac94729e3ced98aaadb3392552e7458417ad6c97cf5e45c52626caaef9384281400d7ce4267225d6f413fa689a767ba468b3771c4e28f08801f5c3e8c5ed300ed30d79430b22e46c67c5f0e3ed01bb3133bd1f7a962106f732a927bb202322f3667fcc4187f3074fca45b69b38cca76a8efb472084842dffce703317c49f34b6b129ba2b1cd8f0f314a98cdcfdb4f19e72159a6730dc1633b1cdd34025d8fcb4f128856c49502189aa7c00222455bb8e3799b60e4fe4326f4be5afb4ec732c7a2adca49a4b66fc4ead683ca3cdb08332fd6a2f77032f6946e4fc57b457127438c7adedff217c18696ab46cbce2aa69974bf2279bbd207cf0a7951535cacc9d4b6627cdb16164eaf4fefddfb19ef93a002b9f18b27e71d6649f011ab8aa6a394966f8edc63f906310ca2a0c67a74b452ec5cb75299268231425350cfd7ccf45205c1d065e53b14ad2f79b77084ba9659392a482309900faae4b3ec48b9debda9158259e9ac1cbd69e07d29466fc3e8d5c6b1b7e164f1584a61b59fd7ab1d21d6ae0566c4e65a2a8ef60e539298588000b551abfce00cc4b7464801964fe67a069e09218c3823a531308d5ec08b4a8a890654c8a20f1e6d9f28272b131750d0d4b657f4fd22513ccf72bb2b68325c669e831977a673afa6fb55ebdda09db0162b6aa140f3ed1e01bc6b5d5b385863a611d02e059f658491414de311128d58d9ea3bbffe648d631d918e56c34d69f3038d856f6cb3657fe0bdc221e3063859e7c1868868a1b58959cf65c972f1347546bc9eb83eb95f2d3ce27cc588d7d706aa6d803bc544b67a790976dc276c0fb76daf38973096a5ca7f23cbdb264c1af8c6641756be42f5eca04604a7f4f4c527873db043d2da2be59d9066a21a1bc4f4159a4421841c0729f3d0fe098312ad4cfca2ac56444f1854d2e8e205499a9ea6f8e522526792a8811df81e54d811ffdf50f8c7c1c03f384cb225bfdbd7924156948b93a6a15aa8ed885cf2bbf1eb4e8268e95612004e1ec852bd9d2fc41559f562728f1b44120a97556396720fc9dcd230fc33420fd3ed58064d3010ed1147332a78ab7460e3cc580c0f1ba79d8122b3eacb23548cb0dbc3a892ef7842b90cb1ba075ec4a74107f10e9f8b372806f1b83f8b1ec3e338eb08487a80f49b3d5f2b33e19c67ec15325c064c8befe1459ff1e4d174d03e444d5d0f941960fdb20d45fe6ea5a080070c385ebb5398aeb8b51d36349ce99de84ba73b64882ac5b73146fe20e4353aa12a08813b78591bda0977e4579568970c4ad2e20f833f0a7068674fb35ebc80904d701d6aa03abc1eb5b6e66c1eb3d6031d665c9b82533a1e9992c9a91bc5cff4a3c1ed12c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3684ba1e59b3c4488cdcbdec22443387b2517900c68bb58ae100bc44c9ae442a6a1376f3a46e0c534aa00b385f62e2b2f9d7099c30f8e0df15b067b9615a730dbf6dc8ab6fd78a0f0637e578b44d29a86d9e1ede98aeaecf9db115ec25239989efd043925ad9c8534f96b08eec273b8e1587a68567a03a05546f3d37f3073dfbd08533786c968a802c5adfc2e8d304aca04fcb666eecfe24300250bb991c5f2a26b9388c4077dbfc8ab9fac42d1a7a96056c597b20282c34c680fae4760eeab1d88329e209de2e75ba5483eef916309652665c986a193f86086c25f591c6af40d7eb08f6b5b0b47f7de0ef6180d6e16cd39e05a20e8c579dc2e556d78c65bd4ef6fdc9ca1b12fa419e05120ac133bc30ecd694099672a720b0012a5ec9d39465420b79795ce1453b3ae8d8c09378f4dd128e9a909a5cb1e6ee94bb5dde84a80cf04b5ae49dc5e185b841f0c40bf82ae14354f8cd61fb570089e8d23c642c2c34b68d23bdba72fee2c1a1a7e8d8b3fd42458ef32a2da6ad180ddeaabac93a20f84f1f60bf985041efdacc32e14832ac7b847d969097048c9478e90ae7184b27efcc3c0d492096302d92fe2b33a8400bc325b385a385ea7bb46a66ee09ae45cb4e341b930aa4db1406efb7ace1a3cf60f60bc89e3028ca463350b0ce423b9bf9fcd20c8c5ea12fa26afdad1a1f5013a5fff51d35d1cf2b937e94cd27d5f95797d7b673ec4959b3f5e86e91ea064e6635850e581dde689a1fa162b40c12783d8239773ee7c19f46ce95feb49302db7d28d4d1fbb5edb55db78fa314341329ae17cb3ea1dabf9b79accf10fcc904fb326cd19ee673843b361582a3c487978e9d65bc1fd70f519dee455caa2fb53937910489ad25a7900e3546de32150cfd144cd98468991654552839e2ef6a0aad666e6ba06fb00ebd2b429903b303540837564588beb310c4bcd94fc69a5500f4ecfaeb063c4c3fe927f9423c8e0a1553048ba715250a393d8ee59cf1333ec6d226654ac0a6703ab672998bd7fc3462ee1a2df2dee3d6d916e8a1a99466999abfe6e06015bdbde78796508d0256506a7e20ef9279ecdac7fef91bddf08a2c9bce4170ac13c012721f1b7d29f70023adc44411953db378dd8d223f16a05afaa127bf8a237aae991db2dc8dff0ab3736debd91249e139384b5bc80597bcd56c034ef7989805eeabb276ccf7fcf0ba33b9ccc202b78046c477a5875b2cd7b3919f5e98795506cd783880569fda5037005070ac8494a426282599f7e92b59dae84db58588a4667e309038f778627e0f1aa6ded0555f1d3c359806e9b07d3e890599c38c606f895e206b674b640d84b237d70e17e39c564848fe73f2298289899d8e35bbfea76785b04e819355dc1ca16024a731500a35b24b65fa5ce51f0355c114d69dd59cb55a00d9fd93b7a0e89de3b891efe11fb109dd213d96611462e458877c59b1dc746b596d1c54cabd425ea2646b3e0da4e83bddd3da0b64f15acb72560a29ef2c5e7f28311c496f9a9e777174cbebec6941c2c096fc296c591361781b5542550aea03d49ef497fcf27d2bffbffd701d33cb49d97e47f9db3e3ef30b10adb377aac2d64fefe46a9f8ecc9b5e02d97e7b9993d1d63e72a90b50cb56210fd888143c85e1770ddec966806c03196a9efd5a37717f82bb5b5a791c705dc7767f461c6aff47920a15f1a4f94d2c610cf79c9b1284d6e47f74b7421076ac824145f4cda56a73ba7074f1f3da6c5439e45b60e0ac87ee25f5ab2cb5f3368530e4de3251c53fd9a033303e05ceed9e4d9895756b713d0916a2f63f319b8508b31bca0708c2217e554e0b24c91ea3699b77bb20af568b33b2a192561d6cec36c6b25817bb21f0c3d9540a62eb43954bd2de444377584f3361eba347c19d673b4ab6358388632f8aa79a4a2bd68dc9934ecfd5257550617826c9f279ad0a21c650c817c4eff11cf533522ed5f2c913b5e002b3640a617b3ef0ed19859026f22691ea90ce684b22541af32c3bde36a438207bfd954f676c67cdfdae5840739ae83264b631741b98eb6bd18146bfb325510c04767ae820165669fbbed53948a7b56bbcb2a62267d65831b425419340888a0178551fefa60f946370ae15b0173fef95e4d262fbdc94f88687fcf5ebad969edc64621a5fe9796419771503ddb933044d94ea65d5ee639f4bd317a9dc519f4f12ed8c6a86c361c056da2fb2648aaf0c165eaa8acc21b321c3d0efbedc1158e74e21078791336d3e59f73782bf879032fb51a85256b805d7db365e55eeac2822b676272fad15e0fdfdc6f819eab401975052d1e498b488a98f0d12e63d72738700ea3d9733bd0567f64498162358c247908ef1024caa3ffb2b65672138780bb4828684f0ad977e91a7004437028215ad0f5fea441bba25e49b9be179a5a4b4fccf79d86fa3a0e1c5e07440d5f102fa38ec35fdf6cafb7f18eeed65b87868540e3078d48d7a6446fab54cbc333fc9bbda51aab7a88b7c406950e3a2a4ba0cb41a095e42282a73a112074a61bbb04aeb06607e3ccd45874413b95d8d2cf7b50369fe52f73a7fccab30c657482e13f23c28bea3d7f0cc91c6c43ad2b7de3db54fab8cc2a9341abeb4b438c55bd6e6f382f71988a9c71ca15d67ed84bc455c1f34cd2583d706c27339559b82bb5c08c3a303b2c7c0e2ae5b65f71c32db736dcb69708cab00cbbcb57de4e5a212ddd7753d6b903d63c48e77114be237e6be71e7e133fc77fed70cedcc5772156a902329d5365884ac1b5faf0e718529b6e5d7e693b2c2e1c000d8c9efb642b306e0db51b7f8823053f4e17bc45e604e01ac6489f182923c260e24fbce13aed5f0d9e70bd9cff33713da16c528c4a323961ff18b6896cf790c87169aa0c97c63da4bcd54399c8b1983ba6cc119ad1dec1e89d8f4b44c456c436f2571b24803f45451a7f3a18ffe04c7b22cdf54aa2f2d330d9626000712ad1bb50f70be191b4933e8f4537a5f33bb1757e65d79e33cf07ff9bf7d90c8e0db0118eae6171efaf10bc422be316c9e24e5cc503802ad72e29cb0b0b9c5258d83a4f56559798216e982fc0c4b22fdc5245ae19c3539e4379f5692354f190be35d401f9ad5b1c311667e418bb1f8029ec4b94c28d2005826df40491478e7c5db872dae778ff551673f2213dd1eb9105a4197ccf99b18357770e2875a7e16ecaf746976bd49fd8224f613bf6de63327e4b0a5217e8337eaff3db22a9a9332a94854da2d17cec2567fa9817ef10515b0b2c97a187c65fe1e8c53da97de3092a5d478abac99e3eae3b421ece7cf2cdba5a8a33d5f2389403e3c4ebf03698183253706d6e1b28a79d13faf21383dbef80aee15fee2ead3fc0dbd4227a31b6a80debde12f9c12c398c75a3056833f7f78a7291822ea6fd7d0b1cf847f4d9a852f22f485e7e353bb26273b2f07ba3f6b7066303a6c07ac0e1525c5d7899656656b4ca47fcfaa3167eb7f9b063e4885ebb7b06dda11edff8d4b614db42b62f8b948b0681f77d14109b49ae56e0b302016edc3b706f19e30c2352809ec573a63da342f81d3e704c4a2fdcfa9c036a7e70e707362680a9d28db56b930af4cb93545609607229344e947f906ce0d8e168c055aa3ed1be17f80c05032c707a95171b83b1857c7dba8ae6c74f259e4b5926800c7d2640356501532de72383e41d7f9b7c0b58b0343d2ad6f2941d254b98df319a628784b299b7dcff05e10d4e07602186295a1468c636ab5d41a597f79326286c62af31ba0b04ea127c4d34751e77262d7f8156ff63b935f8dcfb7d46a4fac9f9812d44185c55eb7cd81a760180f48ee1fc95645fa1a3c803be049bdc9222fd1fdf4a724066ef33dade03c3d7dccad0af65b5f9dd9f8d4f9ccfc3ecc10ec2aed65a461c5d1e6a3ec1f3046c39e1253ce666d146d681c1b421372431ee6a196545807cc25383f3c2afee59e598d20604bb7b8c26eb39a00934cfe26624645f3c3e7238df077d4eeaff4bba174d18926ebf35e62bcd125cad40bf444d64ea1506d0d9163c79b49264787aa8186b69e5dbf0d26424f3026c1730733be8125c26f370eb9ea403da6ec337706a6a2ff9c692d65c4e87e8086a52e8b352d2731d4ecbf7d82347ad9a9f618d4d8e37cd303ac736411528c24f0a3c6aad13f6ce9b1823c8121a1cdef136175a5da3098eaf97f8217fea9588b5bb81d1a6d9f12600271292b764472e29c37cec02a917c9507be7b8e74395971073cf906d3bff6a0abf8ab8ef210f2564c0f3b7fd2264eaf29af3a9367f4777729d8f972a473d5b01765db803ab82853029dc55832f77ed722e471c798c376a0669be634aaec424ab2194428878d9be1395ccf57df62d3ab1e5dcc7cdc4d2dca991335d9179f48139665023693d609042db11d9076df68a53dfdc4072e0cf35faa5edfcd491b4b9c0645ec3db198a41200e9889966848373d0721072ad2191bf5bd606a4c78baa3c375cb6cb5d256e911358b3b1eaf3bf7a6f25d29432b6387d55634786e019a147768eb13f9f000fe7f8d9e66775be3283a1956f551feb51db4cd361bd3c524c1c2bc9fa38d3c140d1092b601b761ce6f3e131be1f2238d1a14928de8279dff5c0f629af0bf86e7a4ceba6c1e7f924a9c28d599df626ba1b9dd361932b5fc6e532e7ba63e7ecff3fcac6adb291734f977057e0c99a8e9d2b727db9c05f8f10dd8385961a5a6c3cfe6a20a7552018eda502a408bdeb4c93e5f048ec00d76ca181c695432910409c9f1690e352c1e014cab90682414fb3be6e3f6c9929aba4b4762c214c50a3b2125c0ec3ca2b738b4311f09f463e103ac77bd0cf8cbc9ed8ef14ed91f5776b68c46b151a5a22bee036bd8f962d856967100146af52a9a32de80df2da84a051db2325d71ab05c640de8cd52c728b8e4ad1960dcc90fa61c7743528f5b5daa7e749304708201b9ccf3be28b398fdbcfceaacf7b6b9ce9c02e0b592f6645305290bc09ad1731f02ccc053a3980338e673f55aa87599203f21d4308a36cc3b75ef574c71ebbeac09270a9cfd806e0688ad9444d78327941b17c6d8751497db05302ef11c559a21cb96889b55070b94d2331c2ef24dd697921c0355b42a720b2674372118092a90da018d6a2114eaf15c27bbddf72e7d66b6c1f0bef49c51527c63c8d02390e04b1cf1ddb91dbf65cef1c106b2c49225afa431c31d1bf94acf1276bfcba3bcca22b611b2efe9196ab50cee738dd790c83f9c8615cbfddfca44fb24efddda24d9771cb24582112a17f9f2b4f286b0c9cbff881695201d7f18393e6aa313a50ffe01e663b40fb5c688a674740564a7c15f5a461f012e766f88c9d7446f5df8616c035513067e2848bd10175890dac8d8d9b7fd960e154140046f608d5ce691a0bdaa5dd0d9688673cc5564e9e6ccb01491f863c4d1e69dbb99702880fe842d3e7ed1f7d622a609641838a953a6f4eaef05d1c841f5d1bb6832913c994902278c184e514b607d0aee04a36a7e76ab8cf469fe3be429a6c6b73f8c51d3f44a0d5f9f87fb3e1bf616d8b885d509c293c8f5ebcbfd4b2992f9104296af709e2f2ea503acf877d3d7c4af9241a7146017414549b7193b034b3b02dfef3aa72b86824e8375ff251c39aec5952a4d8eef766077e412526c12a6c8854410f9f8835ec2b66d54c40bfdf29125612b5d8c7222ed87c231f9c44e18e57f7cf136b32554ada69d97f621a3bedc0e41c3a65e7bec8b6fcfafe2e4a2bb152125c24b502913e00caaff1b49b97d7877681caf6584e87910759a3fd7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1138b7bf2bce870e9424d0ac5b2592f1fba97915e32ea989672aa372208fa4080b890934e976a655092f210b2db9076b906f84e17b43787cafce7a149af8ee4a794dbf3e698c8929f355850b2f78243b3c0ece66f33d17adfa539d8b2657dbb84a1bff479628ab74656334d0782c0787cd7065ff2d5700d61f67bc6f4108ad9cedb901c6cab0093ae3e9d51889ab58efd9014e3c6285686c124f39b02901e8d0858dd89222eaf2bf0b6eece3e6c5767bbc249c87fbf34774636d561e48be3e9883d4ad0d36dbd970cd71277f09ac1e2609258ac98c0e49940ba4d646cc421a18d983dbefbbd95f064fa75de78fecaa76e7f30dead07193d6a0c364f19826ae272865d4c77f9892b65dfd9e3ec374685fa57c799d278ca0e10d77041567789f07f1b1c9be59cd8dacc91316e7d5ee77e019b0f1facd8e02117d82c4caf54bad95282fb2f1b6af86ffbe32bd8a8a78261106a488499c74596e2f808c4c606de031d146704012858754d2ed9cf8eef13f31fad282afae3dc1c5fd6554a5349a446f439a7f932a8fa79ecfeb11ee6cca6a71da25aba0ec2a3494e950c712f4d113fd793df4cd59a02c04b51aeb113861116a543ed28e986e649500790ced2dc26843569e1c9519b7f5c7f60696d848dab020ccfb0ff67aa277b0b79bc3d613a566f1984108d44c98884baa178a95da7384df8d1893ebb926cf47c94e4f15a3cffa76718de30663c66f315dc2a02ae227ed99f4109d71ef00b812b679469cb3b1b8f23848c960bf78064afed55dae7d5cb5c2ad5891c70df3023004a5e479ee70e8d0593e80a9179f9e08a2367f2a269d864aad195ffab5d57c6bce53ffe0be6504b367c38b79884af8977b65336ad933676b42fa806f81078e760b997b4f8ad2bbb93c368d847ff864011455e52e415e27e61938951b0e30074f79a2411295c29b5b7a89045c2e21d7fdf5f4ff1615eb934adeb2953e24b3af6fd26bf975d794f73d77a741a295ccdccb6279cf727dbbda70b8abe089d24f9f16f3e5bf9dde92c568fbe343b36d3f5155d561439aeafa8481b2ba47bc18cd67c261615568f28226c10911540aee36294670468f3952ec9d7192b79e2c13770ddd8804bbb0a03aa544db21b0fca3ba7941160451d3891365e3d89683debddc9b58fa6edac679ad5db62e73e46a592e9b9f599fa57b23d28cfbd26f39fff3f5adbaa777a080c67359ba5bdb70b0c178ff0aafe13a0dba1d15f7fe0b24337c5918fde9169fe4c6f4c6963748cb692e87d6526432fff461b502147d7a168ab6d0824edb5fe87fa21579e8b9372b8768bc145c8ae5d3fa8defc359de1adb390bd5ecf712dba503f3162616a1cc70208db4cd340fea20c718858ebde6f6c56ad4e444116bfd0b05d3070face515b14a83792f746be512057b3a891384a46d38a0bfdde1995bbc483c705920125766e979bee9e2596a06fd44555d7a0f416fd5ee36ab76da927bc4932094af664c59a04d023f8c52eba1cc21c68f9ca8b52c7aa731c8e6bcef54ba1d023803f9e29ee554c3b5a914d226d236ab870518e2fe9c309ac43069e4fe0b1a435ac36abe4464610f725186d54fe1d4b557675dc58d07bbfcbbfce4887e4a715160f926964d0d28556fb341f5ddb1e6237c853d1f934b08ca5f42a19fb6a98f924235fc1c45dc96a2b72e293c46b1d73d34ee158217c889d8e3884c47255bc5b5e74d09fe26bc0062ab6366b34fe6b4d6ff167b98ec1b7845aef6f72f6188a18fedec39b11cdb349e89440b97614ed052a54c80789ef8acdbd6ccf431a3b155ac7389cbbbb43682199f51e14269a4c78e9af2adf7922ab07dc9a2a628faf2fa63152e5cf3deeda3a8082736dc30f7396bf2d73dbb105a49f178f1f7875fa89ada9786cfdbfb5ed5542d2525af97444a6a6e1cb01afb97cced5562de69c15ce7fbaa81ba63e8f5ff33e26b5f4fe77654c49e28a25ab5c5bd30f86c9913aa9164b6888e8b4a165dadd3375ab5481a4687d1575ca8e172110c6c241b7f4430b3f48af5f4b97eb6e7796a8029e8725564ff98e119c63b3d6b9bdb25cb2aeb611bcb22195a59a7e9efad3ce6ea8e5cdd26f9f9b665a6bc9f00cd3b07f8325079345d1efa7e8474633f393df88097bdaa4d4c85c554fd947da53ad5c6f79bb376a2193f260741ecaa69a008f010e2332bb6779756629424f23e7ec88363ec5a433555bfffb6a3f3b033a90dab35382e792077cba242febf54bb7ed38f113d5e5e4b1539cc626ebb18ae964436afe1c00cf916ac3769e1c544b5b44fa7768919569a36142c708551dc96a09393e057e6386d52a11dd7d1b11d55806d724e210a1ec11069ee868b9afadc0c41386f3e537e1cb67d1e531ff0047f0842b71a5e2fc80992d6aff0051614e0d1bf44b1713c7999c6b5077eb7927fd7389e3303a16c55c1d97f702389ded744eaf36d5d327a0577a5586508dba1ee28ea669d2b6d629b07d4f517fee2a59f6620366ed15a614231000a11822b91f637fc0dff75c8407c796a912dd771e707b5f1a33b48971c9e5d4a5bd22e4862b3a6b14edcac20fa85bf25a644b18295e025ed376318ad1f269d2606488d162c5e72107a09d8e585ffbbf3c4dff6b925c382c1d0827757b2338bab86b7e449cd5290444b9d19c90c5874aebd9cc163d21ca5c08ebe1a50abfaef8d012e9b5c265add082ed01926ef4e21ffa071091da2be11ac78e1c83d7acdba3c7d84f54fe61c5b726011b98a97a3c8bd1cb20b5e2b6713c4bed89ce90a0d405f88dcfc66628fd97bd735de5dfa4693593430981af41636498ea46f5b28436010aaf3def5343a21e4b04967e5b29685eb3439c3eca2adac50363a3704a993d5cafd19caf538b6baf9c43f748a46bafe5014c71817ef544fd9c7a97d628377404815bff40d26f866b17d4a28ab5b5f9f16295a3d9cceced1167c1011e6276c2df2c60bc39ffeb25ee894eb581ae2ddc725d5c491433639ea9d441a8d96a05e28f3958e30fe4c230310ac1f9ddebfab55e88bcb4936a7c823f58a7f378031a928c75f551da467842e475971da07b3649d9bb754c0747a14ff7a2b66226cc00f443b33984f2df4c682a35163cb0cdcdd19fbc4a94461e66ef975d7c63a86ad42541a80da0ebe33775b020a6c6574f46a9f5320795e7fdb9b401c593f96773d8534612fb41f92302278aecdd2bfe34bfcef936e29f0e44bd88b971468643c7892d33ef2ddf49b8459028605e22ce8f6acd2646eb8b7861fc191ad8d6ffe7d433ea650161e024ac88a946d2fc8f25501dbb3949dcd7cc50e1b27d0b51619dfe18e8c0b7bae881f013e41947c498b081dd3a532912f2472272d3dd7dbf01d0ff9a10d66b6190601f62f51e2101d937d1c6fae19e6141609bb418655fbb453c72081cae2c5599c43b256eb3b2196ac68f90768a258bc629719f74109354407957169dd533e9a5c5c2f044cc8a45c973b667c22c0459696f5b33d48c5e4ca256a73bd5cab5bd2afc4ebde28a3cd312d8d3229e52ac0b2b369b1bb3e9e364833f4137bb6e67e863ac78cf36100c722a76accc8636ced3c52d92ae4242014b31390f1cfddb1f892be2f536e393328aaa58c89bdb045d75084b0bb890783d6208bd907b2ed437feccf66bdb6f4fc463468af42ac615d7efbe62a97e47b1a4c978d861ad7b1eb69437659aebe95038f408674caddd34c3ebd001b64ba7e62a118899d8629abfa6a56bff3bca7130ab329e0a6926468570992682c2ec2bc5ae81a1fe549f9d742c540aadbb315c6e775bd65daab9a9a0e28dea5f2b3657b8ce4494035c8259e910bde6577582defc0af74d01076d2249aa978202dbc3d70b7dc717f7eaa80f2a2da8241ebfd9e3bfa69ecc659a07f2d25f80ecbbab53787d74c4fa264dfddafa099ba13250a94e3e9e1db65570b228c78af84cd52ea96c642c8601b2011d334749f8fd9bad357c5e9c7e9c0a539ad54b6b9c28e81f2baafab5e0e948bb25bf5086b125688ae3b2293b268f36b924f74f4563d94d55cdcf06003e96123366fbe6431d57f206a43bf899442a137db661e0e3deb4797ea67af5302d100f4cca1d77f900ac983796740083bb218136149587f81db6c435e0267355aedf1c6811344216cd4b8852917879c6b6e0faba3c8d0656b212135179d20fac3a431f4952796fb5031286627b66302b2740323fe77961c5476bcdc8e015f197ad8bffb51b26ad6727d80f04d969066b1d06f22ebd298c6256b9237515894b41357b02642ec678421b0dcb7a2713ccd9328070952f50a9bdb7f7e9385fc10c599b2b82a2fb8e39590e7717364485edcc217da68475b79fae11951c5222bc8311d38767090422cf98f0c69584e086b7d62512e192ea4c938731cf7b1dabe6e0122d9384d8cf8b18267582ad842bfdbf56a26be1db6c3101bfafd7037d19ce507f7713a91e94accead5223f4428420132a0dba3d389a6e2115867d9d53ed99e42107f185494d06efb685327fda7b6ef393c817f32ba529ec5bee5fccb5b402eb6a49fbb3267ad1d17beead1dbaa59e5d48ce46320468db2c2f0e8d4941923530dee59d47b7a9434adf9a262b4111513234d4cdf36a9d06b33ee45ffd7373ccf5fc91a248879a51cd3f297741b461e9bd7890c3cca617b2124db0bf86a4c852a7046bc7c2952c7afb931ca424858882e7cf0a357b409eaf87fdc9335b05a963eb5b8ae329d347fed2a6515457298f9370377dedf0f3912c36d84366cc7205547b0acef3e1ba516c846028a04404de8cf3c9b4ba5a5f3e28c98e0a93e3e723e87fd6e90d4d5c7e2001517e6cf48e0b64dee594fed2175e1207c245485242a281ea4cbd1389aec934b3303c822652c57d9d604a06c3b7cc7361583ddcce62ebdec99754a3123ede6ad3dedc21a926354f8c2962f3073111f151c8abf993ab0f050313e3001c7ce316e3248f9f3d8fc9c51b3ad2668d05dc526913765e091e81cb6a1e5f266bac3b6b4391725564449b35711bf1ec9162689d113f2d8b5caca2dbba256ae3ceecaf4202187a8f7e49c98f7e51bab5c02b8bcfda8ef0efa6e1b256c704892c9241401081cd35ae14d763c797f1ea044533a420430bc5d53444d305eb931427ce0176dce7f3c6698f8e184566bdfcabeff28d05092ab2f99f52f09d844ff7dc820d0283d5344cb35ffc8a7c5e2700d8e8639dbf6398bdfa27fd9d1abb6c715b703a1ee5479e7e8609721adfbc614b428ef4fc09346764ca2c140571407c1011bf95afae446348420657c1a04bdfb6241c0a6827f896437220c7562279ea960f77c8c3de3b7f29cf8e1a94bddfcc1629b2f0d1f7d3a29962f62e6d468b00f11476f0e4abd60a7c47f52eb8bc06d8bdb1f91a71e69fedb8d5ba7efa0dc5c2e97c47156c2182db32f3b23af6f1c4520eddaf92026de3bc03f89de7be9045d627a1e4c4a3a773fe7008d3709c2c3c849a7dc5bf7da8af841d4496c4f1f1a88f84caf87858b9f3fd20d8be8df0548e99681e666eccb026c378d8f452f115b9537c517d2a8fc0fcdcb211716907f6cd9b47ec10e03215698d7c67b8c16fd733ea783622e75afb5ada09423cdf33c7dddec427d44d08164019b573c51cebb72838b35ae79f91d1b9626cf1a38cdd91dd69f95bdcfb6321aad6b85d68a338b1c8499afb9ab8c7c37037affa5e9484ed8b15800df3a749e8e1de70ce9bb780ae6aeed33212e9e015ffb150e3781840b983ea3f2d735b76d4c509504dbd3a888a33222a0e38c0bd030de9a611a1dd17408b941928685a8c745a0c813ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h604b711837cd06037192c524c42b6545cbf8655ae023c47863da38ab79096d96090b5c6815242b5bd464218ee9fdaada28b75fc19e4218aca14b3ed01689c2e0ae6216d5c2746768c7d385cd94717aaa1fdc63e05c13d4a169c11cfc97974aa5b7ae0b59b2638d6fe0ed12604d51c41d8ae1c8ce68a5b33ed7ba8d1ac4e441142447b56a99d41e0382c7f5b6d47d9fb477515822baf0cdf15424a45ae908b3313eb33a932fe02994672eef3b06ac2dcb177b43afe8e029b52bc0ad8981a71a5ed1a816e3c7ba6b8935b97e7b7c1c54c90dbd57c4975cf4a397b1073d2de90203602559b9dfa456f4f2efcaf733d9339a89cd137ecd06983940f5cc5de6a1ece0ff15023188aae61fd0a40af0213433402ca130d7e7f23e3b50e5347c5874776ae6e7e7c9f918cbab188f5411c8652fb324d1f0f2c5c7ea6a6f1760406bdd487b3b783035e56485fc0332d5c75f7e15a51f981725b45ca464bd57e68439198e4bbe3abdc6f991a09b78bf9f1d415569150ddc49601e121f968c37eb64016979458842e87450bbef44f01ce81780750aed834f9843b6e8dbb6c4b33ed04982271680590faea9424444c8fa30a304ef04667aec81b0725daacbe1c6d573b088a68b170ab201279a2e5851bf835110d6aef0e68ec2e23590d28f26d443673cf2e531a12c58199c2040f62857c0ebdd509cbcc62184c11830208ca7a293f2e7d4ac776df420f146d64e7be0be2eafec3b04d0a7ca2bbbccd4045b782073cf53be5cde364ed863bf286db728184ad24b7ab1b05d3331e1c800789eb36fc8d21d61af7bdd8242f4cb7b32448f8ff71716176cf0e4cf3bcf610cd912a8fef2dca9edb657f3f960bb584dfc5b3f86d9faf0b895fee775ed45c639710145c5eb687f5fe82810ce86cb059dfd03cca41ab6e316007655e8f59a2c90d6d13cdc758303e067d45914f44a4edfb069d0e0e49f644262c82f991806e95dee74f1c3ad384dc27ecbc4857b2496945c0324fecc11c8556502f13019315bc916f1bfc4cd6750824b7ad56fc8ccf3224cbd994e6739f620b3d2bcdab591dc9727807a2d6bcafd026234b66350c4d88b01792906a601154a503bbaea45f4e44731bf3a80136e38da8d7b9bb6309500e573a6cf9bd72d00e936270a1ec7228283642c05454ffb861985f1784988fed53df26c7107d966d8cd67a316fa031c8efcdfc8fd1dde8498f1cf40f83451fc60a826ec6457be69479dbfeee7d6192a1271620193abe043905d108d85719d1e8700578acc5a85ead8a271840938cdaaa4c6d58fa41b5d1b8bd65f0482d6aa42d17f2894a1531c358b4b31f88453b54839f22c3effd937a08fe923c8d43d370cddb77c9a2744bdaec624217b4986c7255770c6fdc99fdf00dc341db9ef79cf89c4c3c3ae96ae497006c1f7224c2b21c604de53769bf22c21e8cf1e3127c0c7526602eeb09a72edf3d0983ee734772ebf4c84530fcd54377b1ddd5d5989cd7108b527481de3c6ceb1b05f0418350970b8f3ad038b7ffc0e4192d94dc1b8cfad8d72f52425218eed2ba345942ba07483fae9155fa4196d3c340145d54adced0c4ef4f10d1d593130e012b9eea4b3abb96d5119016f6bf00e6589b6ad8569393566fd13f82de4514dcc90d6aa8e3cc9db0272709e0cfec4f5dc767fb12d9d8180f619f1714ecc17b9fd6ca33c454dc896efd27c9f7741616118083aa1088e63c6534cd102b2f72544717ce8a8013f30e27f66b07b93987818c6f52b7cb5826562ee2f8617e864f4823eedca8aa771a8692a2acd592ea6a151c4ee65631b53fb4fbc9db39b0a117fa947b64a9421ada4561a84c9459d37f49a0f7a4d3a0bb6e31e553ec3fdac7a471c9f7d1c05a00cd9ef2e4b0473dd153b3a0eb023c42e99b9e3c96eeb2b086ff3411a425ab0cf0238ef6e05b4b10d5339a87a5f36c3ab4d88086b0cca5b03380ed0653172cf6ef5c9f57f756e68bc37d94cc608f0d3a623dd86a4f7f36b43f422efd9dee3fa7ab3f202ca72678c4c17e58720093e7b3792313aa8e5fea15fdcab4c06e3ead29135e907982f9ced8ee9450d0eb1dcbd1356b2e5c238bc13c89a753a621765810ece295041e98b83c1ba07a75b27598fa9992715e4c22e60d9175c14af495719ca8aaf2b07c4d3d6f5582cbeed45769d4688dfac0faad2ca242070a4c63ef9fe45e30e8e99904adc60340196b60dc565dd3e8e23e60d222fc204d1a18b98a0eed9944780f1457c02514655b195be33a65735321fe5f73d8221f57970e08c0d0dd31e2d7c06ef7525ba9653c476baff8b1c22cb8cf2785670a6857605c7829453dc25ea78fb9aee3e44972a1d27ad5baa883bd5c7153e822bce67c446856ff7ab69036ab46b2f486bfa445ed9edcd6ab66440be74cf778dcb81726ec8c8b4b841c3020947eeb108371f0073453edcdf07877c01e932162c3b2333c05174e42f33e7aa81276ba43a5f1581eb5911133508f6dff100e017840b68a431cb6bcd94fe75e82e837a2586087941773a75b1b6cf7eb4841fdc2d17d6f22530e48ddfb3225470dd6afb4c0d314faadfab08f890f28245cbe5da5121597b76811c488e24b555783c2061839b6a29f3b7c36a646c27e9b8adf00887cd358b50a05fe00f55f3530025d16b2b458bdc61412f70f51e06ba42fddd3f57273bd6ac555b22a8dd3a9a67c945955fafef9cdcd0913c1587b677b106f331665008015dcb73dd0f3be8325204421363c9ebe703f9ed2dc43fb43df265a8b5d44f1c38aa1b5b264773bbfb3cb70a662b2bfc416121983cc579a8b125c6eaa54b9b7d68faea066ffd46fda997f9b9961265279c5c41cd2e217572c19c118b1936bc8548932e8c8c7e045514ec050541bcf0bb74fa9389d2aca6e844027a12960291149ea875773d9af523cc4e4ab18696f0aa20abf7983e20a9af39e6b10becaa313459d4cc35fcf402a9cf5903f3d729b6310cea3349aef25c923611aaa6ce4a0c30b1c677f869ac8c9ab7cd8037d712ef00248b6e8ae48f6c4ae5b7683091c4394f77b8d11b39a4f1c6be08e4cb583c32f4e08d81fbc62086028636d4664fc611a663bdfb8c78d2bd0b45f012092a205854da6575b6b7e7b1fa11865e5d74667ddbdc24b1162f86aa6b5be8e32536655e943659e695a457360c4f5f7e7f19ceed0bea6d8af65e50453ea4d4b28815f90351051e542c63f901ecdcfd6eddf014d9c77d5517ea47b980aa2c0f1a7804d52eb3f0aa8107eabf150e4726885227c57e7c5dbca31f35cfe5d44bf920a3231a52fc54dd52af8d2d4ce9c283ab9025686c5a817b01eb284855a078be3cb130aa161bda17c519f2017591e79d8088b03797b8a2cedc119ab97e8272218381ee726f0d7ed30f79bcc1f5446f5863596c752ada96ec383006a47244653b8bcc2acacb1166fa4b1920dd00805d186ea95db02d9c67f43cd846581199350c743112c34d638d21d719ad23fa327aeeb9693973b5577771ff6dbd484b1e70c4d8304a22deca6367425e701ff4f8307aff8616cf65e1b7e9422875424bf62bf9ebb3e69ddbafc890709a76a263d18b9a81183ccd2f6c7335cb4f153bf67f416eb3b9c1298b229b94667ae2f1265c37bd351bae823ef6bf8fda74c600e1ddec35a2900d43d489c2a85b5533fd8fbf238d4fbe25f4ffb49958433d3866be96d5b96ed0b0ad2474c1ae5f1f133795da102656ee3de5b8d9aebde7737307f785dff2ae0d5590766c816e7a5679af6b42a9c1737e6364a0791b0ddaa24b0cc53c2efe9dacc1a918179716c940cd950dea24b9ad4d6b45bbaf147b02dc8251a1a7085024229916d0d0d5e71437eeaee0a5dfa6255abd21fa4c269555602d3513118ecd8c08d0a14097c3e591ea44ad9ee5ea3916af4fb7f6fffd27d18b346bd29efcbf47be736f0925be06debe3bee755026d367c7ab612e52ec537227080471170ec72c9ceaa6891db7bd372ab749d6b24783aa90477b714035dfcd8fa4cc6aa9e36184ed7a5cfb648e89c41e6d27fb34d7becdc34cb7ccc03feb53739ff6156a3d3865bbaa5ca27436fdeb14f54ff2a7d31f00f16057454f2e59d20de2e6ba6aad0b93e8260222785bf05549f68c609227ca7b3e07a90cec4173e392d1e2911ced4091ef406de87309ec8e33aedbaa835f6cbcb201207c1ca3781ac3659cd6dafa91274f0c63fe5e39dc52b4c2b47a48cdfd827095cd3cb76e92884a80bd14b5e3df7935f92f47f39be29d0612da45908c16241e79ee37e6272e5bf298050846a19f035c470e1b8b48c371acf5b0152ba1b9ebc757a3163fac914cdea366773f8ee1e2de8bc93e4801fae6ec93e1da7a624af3660d05096b7e5bdffca9024c6907038c7e085931362e7080359b28e11c1ec5f516340833d8abd62a05e6f823ef9c9eecea47cf556c55c5294592883b249a63dfd5980501cb1b6b8fdd683de42873d8ba065d76a68bd58442dea44816bd78b49d78488552ec1535840143fcdbb0c156851234667d85419096e52f3913f5fdd34bf8166a3c068f2a1e75ff5b91cd58b183e7e66bf1a3b6d97f624d494a869d6fd0e89d9180864afbf36013f43991ef3a557d1fff775590b12b4b59d3616748d79dd8b20c62905a395845e24335bc2d456fe0d4594729880222b4b4cebcd704b83e34e981514df9f26d02775cc00f88246bd66616a0e7ac55f6f6090ad93ab6b735501dbfe0129311a22e9e08420ea3c8322c487beee9fd9ef9c99b43e134bb1cdb3bd988870e68cde6f9a9e69d763ff8aef66a466639a5b0a2268dd81cfce081a8a3e7f55cc724006d1f3de0f51f2bc818302a7f5a478a81164177cc89c36773367887b2ba7bf2d9b6a5242af69673d90b2f0169956b2a528c79d60c31e706ad026c790a9379d282acbd8e7d99fb95b87951ce9d3dd93ef4108b0260d44853c0fd14cd691b9b9f646c22aedcb08d0a8f7588bfed1845d64e73d8d5f36b4ff4ad98a9b04d1819b286f5fd18a8f5f71d65c5b3f47fc2c4faa455971a0fb6cac7727924329d046dd7eba4f28daa4573bbd1d33d1cd95d99a5aa342b4803e7a3e72e3db26fa4f80f36b82c2302703a266a880549788c78ad1d31feaec734f20e7d5b8b88b2b254cacf6efbba5548f736faed429493f2101e43b09b41378583cfc1255a3aac78c4cbaa4b6a12ab63953e3158e3a7195604676300cfa1c9a8ba959c33826b3858480f33fefa5c2055547bac2fb051f5a87f9de8d64f71649be336d471d1e4053662545775ef40e1663119969d94a98d13a5c739609203c0cd2a7a32fccdfde31432afd20e64227f33ba90a1c6c0a2ff6e3cac8ad70d42cbee0339c3de0f6d13176f36f253518275c4b6a5a33e8514ab12c69ed32ef1049977fef7c78bd0894270f9e961fc4c5474eb0228664d0db96551788b7c19af75cdb87881a878290e1c3ee124edb3747311c14a322be89db7a29addc35ab1d5792fb432b1950e523772e63bb2a63268cb7994f09e31061d5c50c5ef780ce805fa8ed677e44c70e75b913ab7ac9cf7a80c5dbe4cf64f4ef649081d7623c8af7ba27f7ed6ed34b61e3bb925e86e1d77679909538219c2ce43faf1bd5e50f50ebdac3da61e5280cf4091115f3e17fbe6d902e623607e6a7037a22216ebf824f005d56e01be6d462f55b460e652f4cc26279b4134fb415c391fff5aa45c9203cf51d0e24f4098c2d0d38a8b17e819e1f1bf5fa8e2f3fb005857225e19658e806bd93db82b38e901de829ecd08074e459101eb63e2ea25e079324911891eac1a50add956d7c7cd50;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8ea341f76698c32fa34a53c8c5efe1f0a2fdd9db06615b4c471ebb55fe670d8535a8e4ea8d07e9b0a29580b131c0b9ab1d05469a2ad7e81fa3705dd4463e1622d6da0cb98b7542c16ad36bb4006c7994fa398503020678328ad88c7664f5eb7425cc33076e26a3a4815629c6bf8597d8ebd84f606e3070137dd32f877730a512e85ee2c9a250fc68f36738c699f65b61a8a66f94ef3f7f415c127fda90d7f8f0308b0eb05a168517f2063aa3f280c209b54d53267800213b8abf9ec31d980689d91a45e65a9fb191370753956d7bd8fd66119b349346013e09c6ea9a74ab757b2ac66b99e2aa81a7161b9f980c848fb06a268008446a03a4fd5d76f6f2b8f30df22ab0fec2208f76f178d3bda8b24445f43252c5ab57ea1a1b1235c38b8436bef2868b9783b0ab3d5a9ddb5e91ea8d0295040ea4d9bd3917cff1eb9437c408004f46b95236a6fb65a57a0433529c948cb19b7565390fe1c21152e4c5e594a17674b3c517994a8c8961c8956fca79721eb9ad95aec5e3c4597c2a42caf9f1195a0dc068a63efb70a9ec52715069bb7ffbb57560e50433b6ffdd51b04e511a2b0a58b882e6341a603c65c6654e7b1c89c7590cc9d56f64eaa61fad31038c7035dc48cd07fe92e8a18f55acce4966a1fd3e0c88dad2e9ca66ed5c85cc9edb56ae844ae85b69de026fbdcf55cdb2c375a0a64868878593348f8bdfa4c5686a6e6781603dfcb3f3ad4282834a8a162f19ca1d53751f55863e27249a440c8a08dee69033b6cd843484d16ea612c9300a733372e667482ae1f00b95e1cbce641a05e17696e8752fe524cf8b145f8b50de76fe9e52105ff839152047c3b14d70cfd9a8ba1c59c6bcbb25059921141441a4caddb106517cd1efdd0422fdc6e5f5f12eeb358cd913f3f286e1d5f352ebe8195871a82aaf796ab5dc4d851f256e955d5821d1b767f05851eb86d4cf70ff95738be270612fc8938661016a557fb01fd3ad1aac33bbcbd3e94882b1dc434721baf22339d6d727bd18c3da9b913dfe520f9d4c549ad16eb7f2a17dd6886978fcb5ece85ef57efb534d9ecde10ac938f8b43b52869e1028e3c9d989517b4e3edfdc96f8e6da5b1908ead386e42ab9a5d86ad7c60198abcfd996546fdb1e43bddc1366af2b96f136f612009dc07e27f25410f518c4d07aaae6dee5635553e317ebd73701243bbd7aa1cbfbb9074aa7c4757e8167cac7af25db6b977175f7bda5906cade4b296967bfbc69422d0baacca3bfff96de684c20003f5f8559e9134882e80447c9902312e06fa9a774896c3c9de79714a3747b70bf94e1275e114747ae767b88f9113b1c7cd5d92e83c2e8b4ac1cda36b6822a67a6211ff73358df32a3f3e81b4a865e573d5176fffbc6d123ab289c699779e4ddd55e35ace1d6d6a77790ef576c9fe34f9e11a27ed4887015089dc2309c945d77b28ea545f9f3c6c77738ced44489cb34339291eb7cc9ebf414988d73ab1c948cc1514a8d5b582f582b0137f5d274eefc301d49c334d6fcc357ceeb7f35406a84773472cb0e040d51e0882024dd2172efdd3c70ecc96efea2a4fe2f43b087ebb5d96f82fb3ac3699e252f96bde01eed684fe2664a1dbd6b554d6261e7bbc0072a5fb737acdcd8d333c1e6e58a68e68b07d7020532a5d76aca30c4966755f77e4e2e17fe10d2ad658fce683d0b195dbedba2150b413d9b272fa437ac7ae388cb95b67a6a2a0cefef14e6dc1939e5f0b2f62d8c61a67887f27275290534ea1a860a546c8652053fb14fe23302e8fa45ceace9c78518a6bb953965593ca2f60fdfbdb09103a5474e0519bd8cfb9184c0fd420312541c41b1faf9f8e691b667d7a573c4e3a5925f128c1ecdfc54e26f705e01653a6fa8fc9dd28a6a76a562c523aa5f23939cf8566c56d510b615920b13c1310c24515d70e043420cfbc421c6687398cf76383a52f2e5a251f57afa828697dad7f9c7f4480a4733e3a5ca2304fdd00b521794177c79398275ed36aef175c0a2c3144c4f1ae7a0505bab4ecefa663cd88145d29d0f66f1fe0880ec376cc68c360e9916a5acf1abe84f554c1e16bb0865343bbf8de243324b10edc063e51f6399c57174144be7c393d8c79d0cb7c76cc03e091e440f0d6034bee6b9a77ff30d9225c2f6477317ad2a7dbd7caff8206eea4c9c341907814032cf9024ff1e9947c8c44af9d73b896659e0d6773e09c38b41cd61d62bfbce9b52de8b3be4d5d3526fc003bcd60bd285e3ea56d170b410fdd8d1cf1390e1e039d917cf1ce14359a2ec539d7c7472db893e0d987182bac2799f6b8f58cd20959422e4dd5d54287ce71d9158c223a6f2ede25393d077976fb4313a6f8fcceedb7de05fafb2ad9fa84e22ded0df09a3860fe1aa16a814f074a59fb9a8057e6be9a34cb3e5736dd77372ac8b846cfeddbdaa7fc7482f6ae8369efc317278c7e4f7df0dae41b63085ab7a98027d550c91c955dead16b4f27de5b78ba7af2e92669cdce1dee3430c35e138910438e0a67513b60dc0f92edf4684a035a9949eb3a5fe5a6eefb4bf3a3029f844b83041a82f07464e2ca83567cd89bd57f62f0e1a032a79777e0a509bdaab33f382a98b9c90e12abaf03cce2d49c8c138400680f6a1973a9c7037943b920fa18a7de7b05bebaed15122ebb813bb088f2569335307408325daf03926fac462add414f4e7f4b0069898bc7aa7f0bff1f92bff0cedc76bfef36da84c81741bdebf1b94cd230a08908b90e87192b446e36ba66157a1306baa52746220ace34e8c0b83b850e04a960f5aaab33fd3b6b31a4e01ddac9cc133294e14e0970fe4b81864b86422ccdaed32f21d01eb73d289b1d9d7ca43b30e04b8445f249aace2917cbd9f1a32a6e8e94dbb7210c979a712432b5b41f5aab4d47925b0a4bc73525d3093ffbf038aa55357d6c70a45864f8c24e683b35f3ac5447aea6879288e2fd00b3f115f23142abda20d7af12d82624cfac54af7134976c321dad148f86716de57a191fdad028780513425eca11c4116c436551bf37d446aa7b7a96e8c768180478c22cea3130b276c5e661f76423f2bceb49781ff71039cff0776d9deb9c7a793b0830dfea0ff3903bd1ac8259cf6d25ed95ac780a923a1531960bcb3297754303ce5fbb8bb31c8caa65eaab364ccbb22bbbfc1e04f696949335118cdbd30cdeacc44cfe4fc9d3c01bb203aa51ffd386a9ee129160f9269a57940cad43a531057dfc1449068953d179b1b29f1e417eeb5902b63c08c0d1011c7f04817d593cefc1ce71886300dd904d2b362e94151308dad30360b130eeaadde47f946d47772ada02c168ef7c90786912ff2d013d251eeed90c8c990e1a1aa99e5ea22ca842a2566a0c08c15da409de51c8096f3179ac8265299b27a6b4266c6154a27b8af28b41f171194e2eed57b0394e06a8f07ddcd573c0763d30b52017bedfb525212c65c5feafe5e3c5a658f4b10903cc948f3630e9fb0290fb07f29a030e1fec01e33833aba42a29df9b3e4f02cfdba53807e093522cc14b67e4a394bc3de5f2149e09edfc7aff198fec8d303075411bca828ddf7cf47fe346dec8cf0801a1ba924612ebd498244b4c545757678197b292c838b9208ba99a4cb04e08204bfacbc75bf4fbf0a88404da3aa1a1757e89d1d1c9e6fc276119b6d1bb107959fc3721d32e48bb7b8c4930c6de42d9ab0506dc8f61f8463b195c49249272582bb8ed379d6d077db440ec4562c3c9527c218e76a6c1fc28eea4ea658f32610f3ce211cf9dd6ff0062115d45078bdcf82b90bdeb36f5298d28b7162314ac553721bb65c4bcd1365fabe8d6e0fabaa6265644cc417e82aa1fbe49635d822bd850592543d54f5e27fa7eeabf44aaf15d6670aaec023f6944828450f6cc1d02d2439418ebd3910de887376e706af16b8460230956071a9e685430909bf96840535271abc1ea8b64fbdefc685c62f8b0a22df9a0ac78a2afd949d964c83362199f2ea0a9db1a15b07ba487d00d2626d4ad2977a925d08d7018f1ac23918f60731cd0a5c42b0adad20bc9c521cebd2a8ebf58ec96fc25559aae5a2f9fbf72ad9934340d0662a73e4948c09132f52a5ec8ff4f82e0343d16028ebfa329583c929026c047375920450bb307ef1236f06d3e6065f907cc70b50f6a4b6554be565da556ca2fe8230ca754258f220116da8fe9501cd6d117275c92e4a7176e7ed04df7e302c5d78a5ba98b1af52daf167799394b20ca57769fadcb1a7144cce5ec8274175269415a80b323065aff72a62c6df3d4986d92598fe8b9427cf9c012b265b15af40c89f90355e305a126ba5fd56ef0c34da5f41a2d5cf9ddf8076824c60265c1c73fe74c633237b66642a8b35f3ab46530c3e47443d619013aa23e5df42b77c1d278474672c3c3dae6a52f66ec62e740725a810a3254d7f81c1e44d8f9aea0be3cc69ef6932930c8c0db3e3753d30f05e5a879efd7f29d8965dfde2b8789e6ec9c0cf0d1509a2e8d7126ba685c6e4aa97cfedb94e6e67fdd3efb0b8eb3332384258ff7129b6b170d7e54297f1b949f8ad994733906ac0fc87653397aa9b1cffc19cbfaa5604dc3e4327c786c8fc04dd3105eaa9c2d606b6440118d6155b64cee3e494ca99dff099fd3fba5d4d787dcc91924e7477021f48960125dee174ca99bf17c55801bbc2f9572c2b469c4c7f4d32bcb5930248a3044a88e1a72fbcd1bc4739c622ae4c10b244a49e6ba33b07ce1f208e26cffca8aa482c86f518a373354af57585a2d3f1fd40a85bf6a45ecda025aa5973c05af69f119ee8dfea05f052e21af955c363ceb819fb59d0cdc64b7d13c9271f8a575cca5273a6c4fc585cad51610ac2815f52ee53c1ee7bff1a4a79b543e184f231198b2f75e9061e7d15384f85c9a434447757bfe73ea8d45b1719a0134a3e843fa6fc8c9e9fb1c93b5960748aae91a29bfccf634fafb94ee1e92053d845b622fe73a20cd9627831651344ec1863d5449738c2d2b5d9636316029694aedf5762f4183e89c96c2df7409874866c8c4e3c38a1bfa1e73891e89ed947512818b30b17eed1006e314dcde8d3998a363c551f55f8f4e5fc6ebce3c64a06e7eafd7f04541697bae1d2770b9a7e10d3a3438eafa65e08b7a55ace7410ef7ee903b1c5011231e3b3fe6f6a100ea41a0134ca10ee89c493ab864d9d5d12c704e094d2da8da9b35f5fcbbd385814e07a7da28188798286121399199445a54d21686398ed5adf4739c9dde6e1023c8a9cf54475cd28f1ba0c91741209268c63d387ea1d9ae9e75ea9d0499b315ecd77d1fb9b64a3cc9a0444c7dd0638222ad7abf5d8fd2540b77228ebb82112eb7a5c04406d1c21c7a343da9804da52defecc940201d8dbfcf4c3c280f9440bbdb6b8c4524e6570670e0d7bea0008a8f151f2a5d328489ad25a73e9cec6d38af3acc4fe5e27262dea847216f6e53c757f93b0110f46530f7abad62c001f0771c07dc0203488b6351a7f36ecb2e69ef5c39f1155286f5725ca99fb1d7783226550169658a2b8cbd231824267540421295a5a7c352fe415b70693d7b7735c15e4ad93d1c8cbe84fd19a3037c42fbf886217860828c9456dd3ae5c1ddb777bee46ce14e72613157a84e107ad97f0ab399e66c508f1cf586d9168f549eb2edc5bb3b7c09ac667275f02d6c7c620bbcda9d20cea1d5bd3f5166938b11f97a95ff0808f1b9024f2b8e325a29d86867fd1f82083d96044743988bca835e9542ce9233ece0ddfdaf6326290939abd2a417c412470d882de115bfbd611d24bc87;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9a8b396f7ca18ae62e0780d44e8efd4365bc33382d9ec2cc04efc108f85df271bbe72dae1f26e899eeb5a24d227fa5005ebcda7a33f4040f611a6a83998cd7244717fbdadce4258782e744f33cef06b2630de753fbe77dc172ab922f4db047b441bfa5e6b98ccf2c217a54fde7e91b430b0583ce1ecbac8a99884f4f6ef15cb919c8ebbbae7431e355198e00f03c379e41a86e466c08e3203d4f97bfe89d0d3530e3c43307e69f0f44017abb2ca2b76cf2bc688f7720b9f41cebd23555d76dfff129b7756862986eeaf359456f0ef8cd3aa864146642525a7ca8f08832a82d539ebbcd6dc38fefc538b065a8cb249f5c87cab2bed97732aedbe08a87aee40b07246d48d175be6cd41915491867529fdac5c47f387cf4affd921eba6b9f1bcc97cdc69bcfaf2efb97bc36a6678a44f62d3df3be2850699b744a20b0f704b183d5dece3678760ee6e93b3effea83b85af78e84bade83e17ff0e2ce18bfa84aa4e7aa289419b4063921c8832a5f65780ff436a9d0d89cc9bff36d2a811b9f7cd1498e5a0106757179e6bee5b85a1ad7e66cf3b8dde5cf8c0f88c864e48302befdea07e6f85572ada102b781238186d0f43e4dede6d6d53c3049e196ac900188d781429b6a3cb7609df07051dc506ec0e25e6ced643ed0d27efacddd8f75271a4cdc40a9e0f8284c5cc6c26bfa76882070f336d95daa187c1d2609947de4957927e6b532f20ae00533911b50c3933e0d6e4ca83e0aee44da63c67944edf50e93e047c77d36ef7101b29fe0271ab5cb2c3cff6365b2bef1fdd928b1e4efc18b71195135992da9585daa24a60e670e486a90fbf6c62e8c400dd7610373da93c10d609d31f441825e7a1eaa2ffc4662e684fbf56661178fe8e5f235f5686d3fa93163e2f61abff41f3cbf6e3603898a0aeec592ce1dfab54e40e20b8fae1a85d021ce4d7c07ea1e62fa2c9b7ac33e8d80748c043ffaee006adb0ee5d86dcaef2bffe47623d2c43983a043fbad17db987058b03309b26f303686a6b161c70deb8f43167e2873d68d0ef949d94d28d8f9adf2cce16ed3d4af720efb26801872640889d6d2e7af06f49a1d7e6bfada6cf12184f05abbcecb82c284d8b3329306d2e657b0cff64b0ea07bfe7d6752e2a9128f2f8d43be7601a9b3b88b5f68eb3f58935656f5a19f905ce2574e829d4233978365726bf62d22b7d1f37a83c69b28b12e036ea4d6ec3bfc9e731fc9e194d13fdf93fc70c87f26a3b56299ecf9c3863828ddd656eaef82b1cdd52e0724a7f4094b9c6b0c18ff5c9fdfa1ac3958b302a9b69b235efb80766e635a1ed0cd45351552be2683ede77f6fd510d85f831595ca0f7354c035695e119dbbaae6b5736692040192c8e9bd7c01ce74f5cb3aac4ff3aa7f924b9f8b976776430b243474ad561e163a7ffb215cff25c8b7bd497ec47cdc6f43df55d2041ddf358b494b38d2b46647f2f998389a28a174b42ae78c696b25bc8082a80ac37cf6e19e6661d823ba3301d2d5ec67b63b5b72cf5abf12ad82bba376e667e311f41cf537f9ef37257e31c2daf3c79551c5602c7b68c856cb44dce4797ef8eedc0ed6a75fc6951ea0521075c2fcb4b2760d3d3afacabe79865d0056cec27707ce98be988a0da99ad9a39a4281dd755e97124d60d3a34db090ba2995d71c827d2eb0e6287945aac5e453905fea7685f8ab57fa2003ed1534bd59fb2d439439736f5c40d642f28c0477edbd67c0ca6b0b2143e6ee5bc8531bbe4f9500bfba5489aecb8fce31c065eedd305cac1a754bb049d7f54218d38b9be29e7f54af7682bacfc712648ed03bb7f9c61b24450c74a7a7d5a85b2e58da1012e20af81d8973d73694ce5cab939159a22ffb3325440f5cb48636182a41417d7397c1c1aa931c5885d86af8857cd468719e54f85de4cd8a7448a3ae1e778da4b09053bc7913d67225368a2feaec494f2dd26320362598ea2beb80cf0d71e1426bff073a3bdb5422210c8369a0f863dc69ad7763c42973dadc80779aa97683ded4105b03cba79c88e30c403ecd0f04558388f74c62ba06d0e7798cffabe5266278c5c6e157b191b519787416cffc7ead5ec4cdd6d411f1a41e0c9ea126b1426f87f4feb8e142f0787ce17abff39baeb03da1e1ef18b64e6755db6a06f2283f2a8f6f2384206b912d070128c68277a2ecae829e6452232217419d385eeecac0fbfac4d231011304ed03a61ce16ceb65a0ee5f5f1a0130fc69d765d485127854b5b68803710d21c972547aeb7453638fe9d55601523980fb5b6b029a8cd56013c421dce4f5b4b1acf45c238d3353882c1eb8c7cfbe50f33062c0f3c1f4e66d05746099cd186106927a0fe3106aeb7199dfdff8e37ae2b35d95b1b94b14ff815e6bca9182dc134041992d6ac938648d2a62f1f5c27488e65d4328b75a367925653d6e5b2b9fda19085bf40e1c007ec864ebd0ae7e26e909f0c7001ca7ee5bdaa669926032c376544fcb3e256313c9262233f9c026c67b9c3dd9989c1806e6b14fc19cf2203cfda98e83afa3de97cc727c51034e9805d4b0db7c284c13692ae772965b70c5222ba9935d52d290ceb8dbdf74566cf480bd2e987aba7710d82cf205c918e83d6a068591adf42f5c8d3b3afebf1456d776da86a220991d438cbe3f3056e055b9e5ab62a6fb7b6efd4779cd619aee4bf7e41cd2c3fe0cd476016976163f4f2fd61db091214d0afa48f87b5612aa3ed0fbe982f2d49456d7bc9ecb0da9debd5a8aaa1e428fdf0087c8127b1caa54a058d3d650e8b64365b777acf5b96920196ec8dc52a876fb6a094206c60d971e1f31a1858bc8140fec0754f5fd080ae827120f7650e20b2289487cd21d3719861a6f3da2f00084f6a6693310a65f0ef9ccad632f4c511db10a8c52c4c0d6da53391c586f2ea9fd04206f87f40e8894292a6c10d13540175beb64684f656b788e354312f9881bc55b4302f0beb96ac14af3164f470e90b01760944abbcf35eac41df811e711eab21e09094ecc8a1eb1487a52beb9c1e370b47d6075caa9aff634dde043a33d32ff17a315e74884f230dfe926c533dc2efbd7035c4353d2f752ebb6f4db6743f31ff458e4fa6d036baaa5c154f054464d989c15331b33b5b928b6f6d1437fa0a2046b7fa3f0f59cab2dc5f110a5816ab48d5e54128c45b1a9b144f7e9e1f70b24b945700dbbe89ee204467ce2fb594aaa9c494555d57501b8db38753e04abd23191e7131007dc30a8ac10841b524de9a8cceee39505995012554e3d42ad17b0c6139184c69ab16317369a143b052c0836cf3b96f8507cf134a51df1969ab6bc9cf0e6a82836b23e7b2f66c2e16ca016e54999ed17829da9bb94b38a46ec1334a57ff02bc19536e861d60be3100b171ee860a27d76ad2330b3019311861ea4241cd751c9127810f34598b1b123c5af11ab074ca2877845531f85419249e5dc5e385c1d959fd96086062a7a998ad9e2a0374aef37aa0df8ff5e2aa22dde0e47f03eec9994358aed96e8cde6eefa2e48e5de4b40859ebf0c8ecbd56c430328030bcc4a0ad25a20ff3555c7338709a0abd2cf6bf10e70ebe0a80e9633e7bf1003781334f6834f8efb14a5c8e42d38b569ee669bb65fcc304b50ab0346c0f23007a11bfe65e1625d0196226cd8820353c1f71688075cf18bbeeda529a21a4f3fc8cc776174de6d1204e5c08959d72978ca32f1ea464d32aff9f70edbec19c9f62af01b32bf15858c3e67ead0d0f709be9e191a8ef5b787cdfc8d97b0f1312b1a3434d18ef34b5d2d60e85c352878b9748e1edad3cda25ff957c672112eebf5c2c7635016a72d57f1d77eef8b55830d36fa777b224ae00e9fe6786b4e0b2abcbeb28f1b25bb0cbb34e0ee905b842804d24e990f7eaf1257685ac4c8b57b9dfdcb1447b66bf90c209beb39bc444a69f599c8b04dafcb0d0bd997d5fa7a986f774e37009bf74f8b8ec966083aeeff069548dcf594b685c77708e37694d0a0669abb3f4bd6ae2583ca83499cbf70563369f912734c1cb6029a064de1f907917e40120e8ea0ed291f8868d02285c85a08edc65c22bc1aabf82693464998a5059bbeeca9ffd36aac3cbf633a1f731ee2c9417e9bfb6f14198b64cd10c2893b2d204f11c5f3fefc769b9e55b9d313d843f3de95416242c6e3dd3dd27062be053a46e145892e02bb40fa187da775b0c454df2399992118f90c884bc2335551586327222c7a560c52a39040afea942e13df62a18e741d7247ed6437e066883668af187bbc5d561bc9df854a16c0f87938b2b6d0b7092763cbb0b049d6d30378806437cb42e481f75dd3e571fbd3be65b06d58ccde159352cf023e7f904a2b3ae2109919b89e8717cf2325738e72b6ebf90b8376a4f7a24aa88ba5dd09761b2695dcd195042255b3d654c28bc228405eb56da175aed50ca4c35c8937ba0cb42db4bc650880069348a18eaf7c1b529aaecda3381ee120f58929ca8b547088726b4e8ab45b9ff17c7bbe5559ed5e79770a3a0bfc5ab5a95e5841003ece65df66d94dc26af295ef34db2318d9c9d6c2a50cea563f5afe842aa8142f80920ad979629d629178194de7648a4600b35e0de4914346b1ae273ad23911d2ab07b87bd3187a5d07e423732751b8219eb5e065d3e1c688664d0104bc411fe04487a61cec110ade4a1d57f922ebec5ab1c5978c363696bc81d4bbb888988ad9efd1922e0b47e892c3a7e7f42acc145cebc6c766b2a10869424bf77eaf0bc01837ea3e8d95646b45626fd05e8f30639739196bd1e5d964c722c6e25a9661a4d24f77bb51116fc72e77b75cdd35a6f13a54f57990842c3866190ad0b6463e099fdd38f24ee193cc2bb575a0d2fa27d3c0954ea2846b9e539bef3ffdec34c9a28ec918496ea9ed1121104b4a616572affee3e06682d6a93e52eb660676eb536b6337f59b23b6b2886896ae16dd6af59b2d3c86fa40e894579032981134dc1d2905c62ccb9f495448862b2ae42bf29629e1f7f7ad3c88eeb537689f3c9895f38fb98d9d5be72bc54a6278ed662898e31c5089658f7240483c1632f50c3d75c4454201420c440f8f2f4c259663cf865f7dffad38d86b923fd8185b94daf7b6954abe10ca8d36f6d0744afc772fb02f9a7ec0ecea00e9386158222c24533fa898372e1ad2247e636c7a69e54d18afc1c8f179cadf9b957538519f61554c579c01d4484b24b8349a43cb49ea8b0a6744c86be96a80bbb4ee723590ab48ccdec9113d7828cce3b200fc0abd6208736d7fc2a5ea15877801113aff3dbaf2ff64c32dcd354d0a76a2047e36be75226eefae888fc35a36d00eebb5cc151ccce9deae63019299d7842befbcccd838d4e8b71be47d5348f3d266ea2d6b23965edf4d1bebbb30b9a566455cdd2301a293c0e8bb23233948d9025192748f2319ece50a2afec9752b6125397876d533950dfdc40bdd4be3835d103c31243997396e0694d455220c9f0d516cd366ff63ce3ce99652a26f6b0883eb2864fd92b80027726a23870b076153c5995ab7220883c804d47b30a9b7c8325f08fcdb9bddfc887701596ca78749d0dba11e7cc826ac39fa368b9eb536e91b30f85e2e41d002a18f3cf6a7f3a9316299a1fdeec36fc2a5ca4e0682bca02427b67ac7a57a1d8a9b708690b52679bb69318ad1688f3ced587c413386de18d97c0ea2d0ed57be52da0a660b9325b8c6d28a09ce5f0d07641daf9a255ba66b6a83e2dbec9042aa5cf9a4809a57a21202175b6d9381e5de3d0f6663c56ce139cbe1fe5970df3f9ad92d22d82de3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha7ded39401681620aba5edea992e96d3f19824a6074425d45d43895238085991cfe0bc0397260317f0bd73beac59042e3c54a765e037210fb26ad1ce8e23f14983b7af222d73e38fe64dc10deda29db83ddc6b1678688d11499a811760d4db4eef14117808fa523539ae4dd85554891ea5df844a4f8adf7ec5cc4aa70094f3148d9047bb4fed55837c7cec56ecff1c39cda799e28ac0ab7ab59865a29d5183e3e1456a81f264c240645d6a971cf7c2d478e055064acf927f1bc674169abe93c7012f8dcbae1a2c42b4479357b5b846d024d73c6c319cb9b0d94d27b4ab0fadadbc81b3a99aecf12f144d2b2c3f0bb87c72a08c378aceeb14fb203bc5b5f47c3f515912aac98a0fc45154dcc25b3f596525d62172b41396667c2a0125e4d28a61da34faa8bf4bd5b2a114ff2a177d389b6a4f126fc0a94e2fa23be9b033068aeb67b4e39d99738bfa3465fe6bfb73d0c94f097f009d7a66958729b234aa25c58c89f9d77f71771750088ace59589c3faf4d690c80b1124f03322cdde983653db5a0b8dc31a08ea640837f53df3d0ce7aea2d94030b990008378dc5fa325e5254fae1356ef55f5df04e2665d031562c2f52f6703ecdafac4a63c421864b5a48759003bddf349c6dff6461d4d0bd99abe7796e5777186e9c0b2134c407d894e465b45236863602004b29cf27984bfa19aeabc0a1ad85fe4c48430d33714618bd11b75b16a82e2ebc08ee5105a3cb9d7cb0624e9495eb972a3b75af86304d4921bb2c4adb70f2b3d40ce21369781883e37fe9d21f00d2c40b4e28396e7bcf9104b41d88b258a28cf7b446fb80b6e67ff696c398e0b1c17cda5131f41025bf7c8686ecd4a2ea44f643cd3d5e1fd34da35820917edef94d571ca8d0c63d1a36130896e19c9dd346dfb838a041d026a071d8f2e63b7f18a619e3ea07c7fff72ce931c34ccb885de1a1ad6f96cc4bab30f322c99059fc49e202a1e70c3f27e4d0be35838611860e81ac47edeede597eaf120c4be20a02f5d681a06d96d57de76290c7f79e024e13ab24494955e5996dae367506d16b06769a69d990af77295071fee36064c48e37d8b40a03612f2f8e996ae7aba1f48446293095f8c0694b08eb10f4218a7d2fcc1a885cd2246fe75eb9d174c7802b17539c9c34e8ee6ad9c799d01ff84e308502c6204a4752790817f7c5d3dfd9bc5242d875380796c3214bd65e1980d37a28a07d93a4e4e7c9328beeaff680ca6ea73b82a8507f77e2230002c1730cb65c6107c93499e0e789c55858b664c68116a4e6669f66be524aff1c830a3f191802a95fb461f4d2c2eca1f9b300ff8cf81f0748d78623260688b3ae5609112c365ddaa81e2c4c50295337dbc602fd99eebe211a346649521b98c7ebb9439e1deb258a313624793d3c88d04fb6829d791694f959e441dfb9cf48e593f572ebbb085f6e43ff47d49cfc95fee6fff958af1d88c712daeaf56e6de9ca1e3af2260ba237fdd585e8771abfdd49689c2556ad42b077915d341e41433a4fb1edf422a9c71ec60c4c0ec71c8cc831586b7434cf0e02c42a5abdb8f6e31e242ed9596fc379d2639abbcc833e2a096eae9e7153626104ba3fcd8034ffe665816c3e7f8d226e7f67fe4fb381fd4cd43fd4f985b8f9cf2e95fdbc3eada36089d8513389ddeaca02b828a3b0fbd5403922ae02cb435fd084f3d60b73b742a4931ac5b05ef22c67c8f076e41f44149ea1ff950aa7b5c478e5b46427642fffc754c903acfaacc42bec10540faadb2e2dd17e984ef736e4c7a31577f689808a9c264b8df245a61ba650f17a75c5894ec487a6210a33fb0a932457a7519ffec0354cf092c6983ebc436829b4b8cad27922a9462906a6bd108b4533f6bc5c1f3e7710bfc922925f0034fd23d670002f64fc7c662b961532cd9a7dae620c4d7345520da6200e043095d404873c21a063cb6d515f73032f83418791e197eed5a63bad38ddecd2f60f7e736f11e769bd24862bb23ff3ddc2f9d30d820c6c60e3790dd7ce3ad701e9b372e68c5dcd560406f4ca5d7cda26c26d5a4a21f8783be3258785ce6155e7d4c6d90c163b823f49b9fcc389e84769c10a933554870785ab56343e8a24edfbc82c6f78a1d349bdf438a731cfb64d9b4bda916fd44a14baffdc1a5f464aef2de467e1689326661500230e801044d1a13add9a5b66f28d3182bc8e8534625c2ddf133ab707484ed49b070631c191204b137c23d6ff37dc2dcc50a4462b65fc4c304188dc4676a2e6db51c1c9d1c80fa555c468cd298c1a33d206cf4808bae1b61e485db9415dce1b117150d86e0b79c1d0354424f8d0235f638c203c51d6e7af13635eda8a011fac0025f369f4c74fba042c48919cefe41a0f091346d6499d2b5af361037a95aac6edd19afd421b18482a94004757db04be297009d713017d86f2ea2521adf82809f28f700c0ba81970702a37b757f37044f1f770fa419ccd1b39690931fa9f9b0d10c83bf82972493ab3103709ea311afaa9443094cc7bf8e39bbb0a7ab1a91847a13b062b5884f400d3fa3783c757bbd8ce9ea5b1f9492ab17f2fc946a54304a31e486aa7371940921549cb564ff0283e9ad61b420fe39f41b3c251086ebee950e65ff820b6d31ce8472b622aadb0f20b308a2abd55d82fe4e9ecdf34164f1ad06e867d1846aa7193cd88063df79cef092c3e219662c1a47c3fa73a345e3e41ade8487eb1979ecce0281304779b3e9c6e4485f231ea318add96550c091c61f40b36e8ea7da8ee6402b8bb036a4c7da2fc8f1e36697b008e50868a64c322b06b572b23afe8a14570555a880b138f45c36f37fbfb65423740da941d84c6bea295b4a77af6991909d0cc4cd9b8cd48c4ba068c0c55695477bc49ce403746445eb328c34ae1ee9302421a9401a760cecad4a3eb58807cf5107e4c00567f778c93279184fb1e214c3057d5ed0454e4c80f0b538fcd0760385b077b6b2efdddcff942e4270a0de018f0cc54fc0c4a9d9a4de0b278ea3ceb7c2cdb0aa98f1e1e5f183302e80a711c8c1d08769dec02a892b0870f3c012985799ef122435e62f8ec75f3dee5a7269b7dcf48184a4f25c8502aa91a8b4b7e656ec27492581741d6b59df3a51dfd329e5b87df7005b08ff58f612312fe19f386f47fc4de13b3b2eae54510668801898b82415749b9a230978588e809957e39173cd48df319f0d5b56586f8296c6d95a81185ad3b7ab1dc3aa9430909ec793734f292bebdafa4dda197a55d0167fe0fe2ea60c4afdec63c6a52e021486c6699c83584921557eb70d9d4c9dc7124279ab47697e1bb154f1453ce85b95668fdfcc6d637df532ae741e37f3a54975402de314312aa485da32ae230e03841b9e519587369cfebcf6013d9c36fa66da401e2f9b54d43493d95ac017f9a348c49fa3afd4152438d77e7e2eba00853e7e8637973ba8472c576221072546481d9f22bd9e3e79f53604b02c98106c0c5497d3a2cfc187bb1760a45c40aa59d495303f683d0e4481db2837f128bd02d5ccbe1d59b11d2b0f2e69cf29007acdcd5b1265a8cbeeca06472f2c4e24dae51a753602a3522c6e6fe5158e305ec542f7ab24ce6b7c5ab1b34fc0cd9515cec85f30fcc386ee9e25c399dc9c24d7c33a83d227288a2d4845da5722fa8760192d7bc776ec04f81657263be7e07df57fb6d6d0cc762d15d699812672329709a4d05959aa54550f5ee537bcea10e3650851101c3e44988c0b77b0d948077130fdb8cf6760491e9a647f04b1f402e3650a066a74a4933c9e5882982e2e4a11c185f1d2bb6681970fcb0ed314048e31263585ea0b2b6bc0a7df741e1882276cdc0197f9030caf8ebaa6ae50effd420ade9f9ce188c161886588f7c58795846a1fc8a7af356025e42dc0fc5810c7fb48675162d59c6733fabc1251e7b7dd56c02d2bdf13508422548c73fcaacb13f0937e7cc3f8b351c13ee5b1fade059017145701e4818eb2e7779693a5f9839b196a1281d84d00e2695766b4e3eda365122a757b926199369623dffe8fb6bec0b7cf5328ccf2752a4354b33408b5c6ce5171753935fcc20b0d48ba0b067ab78b005197a249500b818d60abf674369bb0593865521fa68b2800ae0989ddf69edf9c4b8b3f8bbdf4917f5da8780ef761c456f0e618e8d319733f248591334302cb0b97db66a8a788869ba606d14f8128466a9b80830977566bb325574a1084dc8245d25bfe1eee7b8c443afceb5c834e4ba9f8403398e712e163f08975056ba58c982afe4bf00fe21e72e05009fc34ee7c6de41a5af15db63675e5ed5851c82b245aa3884b19174662ece0ddb98ee3d81f1a44ebaec6da8acec7f0ff39ae6622e23149dcc1c9a50b3e79574f8e6bd77f6b216256fe962e17db1a60eabcffe9735a9cdae545ab9e92c0350fab98e1674bba37490f4796f10f31b79c73547af3781ee96c5bde73f873cdcd55b7f091b892a2b97abd3880c0305c223e745174fc2508d3e85e29f53af4bd691fc9dc47346a0a68a5f1bb543d12e3110d9a714bd9df9bdc634a9c12356167dc6932f8e7e284b338eabf1d46e567cf81ecf0de0c51108d5b778f7c12916846ce947a01f494d787b58912757c38f7067b313722384aa96da7826d479f22650831d7ebc3ffb651d2aa270e543212a37d7dac94fd55b495f227ac1096859d336622eb39d68a1e582cc54e9b1c9a62ea93a92fcdf4a66940042ab5cc8422ed67a29191bf2b8ca0f75f91984249f40df21effeac0f0beab2494fec43bbe4b533b8a3d4a534095286f577a1eb9fc71dbe4eece1ea7bc1ba37917413378dac643be31b6d88cb56bcc10aebb9b9f2e4616bfce885e4e436519d72015afcbb7f1385215c564488c7dc1e80476808dc318429f5508c263502ba3619fa4256524788b07e9d90703a0d39d005ff7a5cfe4a7d66360ca6ac3742a3136bc6f263b1bd32394c513cbe89a74c4ca31fca5a73483715509d3ff66209dcd058387135d55cae18ac99c62965b993045f2b9521b6ed5211cb29f1c79bc55ea96b0c90136750bd335bc1acedee8274003604ec949283cd5ff5853160b0ea7c1f05299b7c2531ce2a6287c6ece8dc5ba166a6fab219fcd534663a6893c7de6cf143f8d2b24d0017a3bd17c114105d2b80dca310660acd4bd71672cbba1d90fb7b670d9050bfed1b13b39442edba5ff4af3613ef1295babd77c88d2603c582548854dcdebf66fcefc8b5906dbeb6f9dbdc2cd7cde64afd30b585dab5d0c081c55a77dc612c538369e4dd913cee75a1cb7b93164a710820cfc764253d8c655a12ba0b20a53b2264856155c56cef5d284ee0654d3bf97d7cdedb6e39ec17e2687cc08274407620778ce7ffef1483ee19feb1df9e500fca12618239bb8cd96812272d5f95e87e866bc0ab4183baadee8910b4aac1b666cda5ca2a44c9cd5ad293b899e4e76075a1e9dea5c504603b82dba445f5ebdaacf4a1650818652fffaf3975df8bfd76ddde5424d1564d9afbb5bb139d5f61b33fad160f6ca8a87c990790432cacc576dbf6961eac391954983e7db2df666d5bdcf1a5551e1447b8f7d23ab58eab250d16466176686076cb4738a6073cf35a119af8cd759ee91605e8c2a2c6c025872aac9a0b77827596b85d956ae11c73841975745b4b647cf373a1379f25767e5589a936e4d1bc9a12906f0a7eb8b6b6f756b2a0cfc68f6c89515be3e39c1518c828ad8bd078b9a3ea428ea12693ad89d3987fdf89b0ebf6c9baa55509cf6537ca4dd8dcc57c56669b8a35131d50736dfd7c46e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hce63ed2cb88c7bfda1056e952543e132496e82bb606a453895b8045bb9afed5919a0a7b561dd234f13b4929655b6b730baa4a0dc05f3588cceec23bed54b78e906d5deabfd6a4ef7c0dc91f2c99f966b495cd59218f36c423eea0fd65012627ce69d7149bc5b65d3be4e311aa28097c1174d43b29a8ec3dad4c0dcb72d4b60d587dbfd2aa1ef864a9e76070dae60c2c4ea06340e41f7e247726d7b9d9c6b9a28ff2a267bdd222dae9282bac35e0b67394ce2ec73e32ac1a8b9e51743c57c7a49b3fdbd21b50ac28fade7abf5be4e13c99ae77c9eed4a078c03f42079d11c4e893e9f21ad491619e2acf117a30538709e9f759221f2a2951522c4ecc11644903faba6e4e644f815d7b96e7bf8374e76cc3ac929f8f631d3c35693c873f338d48f844f23e498eeab0044191a03412ff7b67109a15af8a93bafd58547079180439cc22cbdb63b473c4641692a7a5be39cbac96649fecae73da5a99d19ea9b583c3fcd216d8bfbe29b1cc36a917f51803ca8a51e9677dff60c93571f4a74ecc2da927166036c06083afbfefee918cd7d57e28c18b09a7f894a9635d09f81a2d87207788841d24e7fa378645f863a2b9249e03605ae4512a1d6325af2a117d8d070fd3ad51ef6e90fdcbb3f1c70856292ecacccdb0326f1eb624f07bc878041c1903575f3988bff8ee848b6c9056db6b76aa535b73ea9116efdccc32bcc8e5f4b7fa7ae0e548637c68ffa071bedb3dc5d2ef73a9163359bd73f0e6892f47993e8e0378c2f6ffdbd121165407fee6431354aafd1a3159275cb4b1d329d7664a377454f2a8caf54f0be87af47eb7b025fdb7753114c8f782b438e70638348030cc1cac34e8f0075d8967ade3dee9a8c723b8e7a45720ac98df67107633f097c0a8f1b7bfecae1516bb6099f724fa37810a18e616e395fd1c0432b25620c916b154e4aec4faefc011c9fb759279fe9bf2e53a4143ec8c6cfa12c8bbcedcecb77295dc43c3f60761c9717a327d9111b0c32a5a41b4151acc66ed2f1cc4b44ed77ba6a02cbef56076331a2d5e34fd39b3de6faf9919dd963f1e0830e3ae25b6c738b68df3a65aece0620c862ce28de348a2d64e673302be828d12321202c3e5ad7863cbc1a4426c75f2c77cf0520b466fa6dcd32a08b633264d9e8e48191fcd1f9be20eeb7c43e4f2f9efb06bfafbf6916b76bd61dffe3ce2bf8fbbfac8e6ad3a4465c4f28bf3ddbfc48eeb0550c142ec07aea29738da716f6bcaa24b063cd8d8b33a69764f7d9c9e9dac6f1d7176b42440bd75d288e570d7230a659fcbd97347e4257b14350d3fda8924f82a64d35c8f5b576d7fe8321e7c2d48b062033215cd026787f39ffe2da42b0f6399b16838161197559d85b450c9ee4312886ce32e9bc964f9b2d8c04cf80b535bb3df28cac53092c2b884a241366fe23846e42ba7c8a21f8e7f5e8a20b77db688bd1dac7fe5844b08fcfd5bf49273032d21d8573f96f833018f0157cbc01e7c0ecaf8fd4faa26eab6444cea9a88cb5517d268a4f468e15ccd8566438d4fdf344af14d260a758b47adc9d24d89c01cc19e2de118d59fb997e6717e8e47865c22e53226abdb03f9ff31ce646d1c103f60619e31688d614c0e46ccf590751389c2755cfa0427d3e6ac4b944b51376154d1dfdd358b4db7df8b9e066d5007cd648e3bd94ba8009019f4e3ac8546f8f62f8fb949a5b1894d96339b3a1c8ac6fceee575d3af93ba88bc3efb8693dffadc572b3779a31161040ddfbbfd79587f6432e4a207f103530919069799e674b41703b27f34ac2e0abf0383af4fbc2fba94582ee7c9154cdf6c50ffeb7b86c047b4688cd03038560658b3a39f7a7097b7b7ee8bbafbc0a0737fd395c81fdb6be40104e4308e20668b046a457ae1bc1767be9ae16e1768ae37c229e175b1988a87feb656187e5b29ba2b9a2b53fb77db76ae0a67b07b86f94845d237421e68e92906ceced33ee752cca19d1309a5ff94e475ae9efdb1a6ad9a0a2ec14278fbd80fb9a6272d9ab6f9e70ae4e9f219047d0aa9feddb357e9e326dbc906ad85bdef4e976a475dbdd79cb0c9aeefc116e37eebd801ca489c9459800f0c89c771c1fffc40989e1b44b9c4a7876cad88fe83417f8c5e91194057c3092469f907b5d8479ad415d32201f97d0a421df05f00f3017c07eaef19fc354aa115d40a73f94b4968a16d4c34173b479d1d8a30aafc3d389bdd0562d3f9eaf2152350a402a94741a52d9455e6503080f75e27333c33df4f8e8eb75da782dc379ae667d0d66a3169f9f539afc264c6039979c82643651db27b9ff9639781336f35d55a566320bf2977341ca56dc4c5939f569506cc92bd61a175b6243f4dc4820655eacc5ed9b0e286456f03232f81597aecb5da15926195c3ca0e9fecedc7d32f3822d9a2ffe9d7b75399dc5b2bd97aab77f0dd2c9e4e53b99982db73db5b312b6589def64c43d49721b15d1a22cc1ed3d14cc6b597a02c53b0f8a0533e3d88ce6a6f55735d501b4c09672f67c352164f1fd7e0aef60373125e8bd2231ebb7c2c7f85a3e4b19ba1cda04183cf8f1c462f41d2567432c0e0ddfedcfeed75759abf1d9d47e3ad50ca72ed9cae6354d7eb7f45ffffbb573dd3a12d62251d0dc2030ca974c1b1b955bb7a03f27c6c9b28b9aa0af1f747e61e368c162f929a1f23a4d2153d6cc8bf19568c23a66ef3cd15c0ea88ad0d5266b9f0205d0b2f0e555a395cc54ce6497fbf82ce8672d13d759688d659d57dc34881a75ceb3349acfce2eba8f5ca8462c25645f041db43ad5b6ae94f92ecccb8c456dc4cf2a3521d256ebae5d222e44816806b8b4c0cdd96938a9ccdad59a02a3d90295c67a33ebecaf509413f347b7fe7e6d16ac24fb540ef943bed483cee6fcd24585d607f0bf5f0e7a2ee1ee75fd1f9560f5657148523a08643cca7fa3e23700285669ed2be7760977a831e6792c1a4729257351791f3bb771c2bfd0b71a96799e1e8cc9b554600868451c850faf960b05b53ebfd1a491c42b6444d4ba62f1aa0460ea13906ea96a2d0de904bf7e5216a5151eba1543d185e9d9c7ca5167dc6a487c4d50747172c5818e2828d32722d35b9f9e3088bc09354f045c3e544f1932309d1b4f229efaea022025a3986861c0ced91dbe6a399d86355f2b3847033fe45d5bfbbf4ee7b427ac9fcaed0b4d08649e4f6f7164fccd0091ab8901534747b0be8720dce2390502a3246bc70d121247bcb03fa4feef14ef6f63c593162a1fe5925a013acd04fbf42caae10a52a4856762b8656e4991f7524cb474bec228d3eeb0e2a686377e11cd34063698629ae249ee717c6fe6474fc228eae01815b5d973265e75630f7eb484cf2ec34b20f42aea94e9f796081a9eb15bd5361bc51a5f3607d278314d1bdd70837a98ab98b4977053cae5bc80df6b6af714288c9ba4350f4e1e64c1edcaba48f2fbc86357a650e7d2c508812c5a7648be9bc8d3c96a0b5f11e3e9d2958565e7d7096343b5a826296d596b4081f7357411d75827efb5d0be98ed0adbfa21fa99e51526368eb710531309d7be28eb043a1e6abc8ec8b2fed0f668946c41c7a38318df23bde26c782c684928867d455485029fe85394685c3f267c3cda1735aed23c22cb70e89833512fc21e9c8aa7169129a22c6b9cde4c6d6ee0a76dce71924210e563322fb2d1aaf1f8d5a0ed081adbe8271654665826e8928a1ac2c46dcd192e988278cf6d0eaeac46dd58f6a7809a4a9a3b6c635f6c7a66f0b9ae80632dbbdfcebcbf97220b143677162db10a61afdd7b54f24ab20b97fc8a3057fd4baee995f424f951bcc9b152dd08a0c1cf7cbbcd1dc97a76dc2797ac8f8d82a695024c0ee446e7335dd4c3b68853392f76f7232a0d0b83e7497bb41629616816a2a3d50e4fa40dbb24bddeed6c4e7b47a96d0fd7254a09e14aef0babb325fa7b357c0e5a083f465fa6c886fbfd8dadc57c51cd8adb79c4031c2099dd5add9e5c01c4bea98aa67e3de28077299b881abcee7ffbd799fb9e7bf5b8e1a592f27a486beb455c0693129e2b8e929dab7340826e3ea95ff920457af4594ae746b5addcc1cb9f1e142dd8cba2d682c9903acc5a00fbcf72f1e9b49400bca7ecdbd9071954b6792b3e546ccfdeb0e23d56749bf357fd76daf4d51be6c9d89eb8e3e1cb3a05b6fe56b072825bb6527858d4f9452833939ee5c51c98c6d0c3bea529611eb166664db539577bf19954499b4fbd6eadfbd3279b4200018f6d8cd608afbddae6a4212df6cd92f23bfd70217f3fca6ec96323f2b76d4921062953e4a8a301fc4f9e31918c11e2031470b84a21d8b7cc0e722bc97ceae7b30e1d0a9e68f0985123ffbae81a8638a2498c8f89886fc349e0e404efe28debc242e465675e2855500789e42b9ab1c2fde4c23914ae57961677e59ee08690317b6812c12a66a5b0aa85551e84d8adb3a73229d0b75e17b00a49084fabcab81c2acec756ecc0efee79569b35beb4697cd8c019f60d3ecec1f7eff3cac3636d896ea38a082b9ee16e060730613b0bfb0f2c261507316dc09becd645ca66e41a7876de0498c8f246985c866efdbbd65d1815a1a92885dfa45de6367a365e6193bf8900e30324f1c406316783d3e018f20b345f292b931ab321006a6babed2b0550e526a04527b5c3fa0fa65d44a1465a4688127f9846005a4dcdf23e83208f01d4958fbf20c2f3dbaf755a79fc5d9335619df28338c66c4147488714d8efb0bb0a5aa9d483811204d02ab94c7d48dfd5422fa8c3594b5f48eaaeb7116172be38cd84d0736e0e5be373210778700dee27d6b81f465cf5dbd91e8058f2b9c07b9b103f0f2d9de6b1e619611048971844e58109dc72af12c99fe6402c462823bc0e1c68a8bc3aef5f54422e26cc0236fcd74c2c00d0b4d20281e245af994be5e3ac0385aef5aea9df2da679d01aa621bbf82bf886955455b6f68f42eaca5b3b267346fbb915bdbe87dd772a330bb639b797365f7050157a28049dfeff0c5175267fba82cd5f270264483bab50855fec418bab29c497cb1554b3b4ff053ff44920b995771315e3c2e4b53ce9d3ca4efd7d1bdf1f460d38cde869f407f4750f06f02948a450fa67b30e69628b7668f3708aadae4763c19c5bee37fd04588d648c5c90201150d5ef819c09d184c7f19a8bada7a870268dcae26fcf692bbf308f1e2ff4cce7b3b54e4b1fc91a1b4a59a4a6eca37d5e88d8a3ba2323828ed58fe9e7bde46c1dc920405103184b3c44b57c6ff32ac966f4b52d2e8eccf9dada5607ef00923ff8f1490a0584f80b9be411309679fa051dd8990685853ccfc47cc7e713ac47746d032d7e88017bd0a475080789dfd97886de17ee5a68d82e86b020b827ced2eaa35eebf3dc3bebe34ffefa48c49f405649eff4a74abf8bdb55adbf26795ba41be074137f90093397efdf08609ba8ebfad4fe7de14dc37ab04dbab75a0a32c1d78baf30685169accdb67178fe9525acf498be935f6bb6d68e47e531069132455465d277a613056b19997bc682b51dfc684d868db78c81ecbe6942cd4697936c9d8788334217288ae255a2abd0fe2896c5e3bfe51840a3f46786e37a23abbfd229455e799ac601659353fdd184368d36b9e75d5aadc8f2b67252185615a2588eb775589e861dab9b7ceb9fee5bc631486fb2ac844e40c08821895dba7d3126a99f9f2a448a681110bc482d5c5005be921527ca485fed1e8d5d71f12a67d9b3070fc1a5d3dc96073a364995980c0f8b18986ad090962fcc9151de38dafac5c31f334290822065;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd3607594484407311a7eb3ce815d745a45b6ae9ea5c8d8f25e729ea492a73779bde13ef9e05e88daa2a3231d9ea6ad521c4fe43c0ae7a0ab3599288fdef2de78d1717c882fd8388be82efd877efd4cb376c56e6d6fb894bf5e36e8f3aef277df32fcf28844c3a765c3a621bb6d543a6348319703a07eec5f3472e6713b325322afc08c5b71e9689dfbc816a7844074f4481414651794ef7a16acce5757da44f0c8f09a4ec27630f6f43a29bae98fce75c734bbc1ecdb913a3f0b15eb092b56bc817567af23fd40925c10ef054d8737cd6b2c2ff58a214426ac62e1b81cf7a77a1cac5a17017fe84d8bda9c4ded4d190ad824ee3f61a0dd35f32b8eb573cce40a65c07ba2873b9b5466098b888ae9189ca83aa9a4d8253fd3de13ee6a7efec45c16ff2f50114b2b5a45ae5d9bc81ff730d451321832957f98040e7831040e7263d161ddc23615e142b0d3b1eefc1fa6b657c50ab660529bf1953c09e2e4b371fea939c59a5a398132eb174362ec21c477c6cc55b22fa49220e7951ec62945e47ac2072e75c3a6185ee97183951a4cc5914c8deb91824d94fa376877dd2ed074c0170c0234bef2301d772575d6981ded8a18a7e57b423a1c7f442724fcb204fc5c1331c445d8978293f0b960f18c59b4eabaf8332f548c8eed4bf58db288cb0a9b973504e33d504adf833a9a34da3010a478f5acc1e35ac95768ce9d8e9c51adfe0c4fd76c8236943615e54175a8ea502055b4066d35e5faa2619325ce7248d7588b12096de388776f479a06cf6b2113dc94521509a1827155ce367fb71516fabd5364bf08b216fcdafec1b3c27cd9a93fdc76abe298c8543da6091b2bc4cf3e6bc15ad7ed413b0a8a0b24feb41c53766dcee0e67a8355dea6d7ab7dd9e5f67c0bcdfd12bdd9e62cf25be1a4c03e5923d12d046ff49d74a61a6400ff9ea33d0dce5b431456c43b1c2cfdfd5349ec5dfb94b819521bc755ecb8d659d476e7fa47f81307fc45026c9db07aa44ccb432edc3f82df843e0ceb2422d7584a813faeae9dd2303f5610bda1d7a178354de661c55f9381ab6731c57ccba916ae8abdd445e70ab939a528ba928ea70d37f85affbd4d5f463d6a469daf9aae9295602f10adbc6c5e273d8892908ad94c0826b3f6e7edead621389a19406530c6d2ece2c9383952c5f0561e4b6332f81c89b414a662194a6d7cf3cd83d11cc9450fbd5a4ea05173cc32b5eef357fea795d8a07fae85b526c2a97012814ab12ccc87dc4f0eb98d5d8c02049abdc07bd4715207ef45a0bc3b0a2bedce50a9361cc803a3669f99fbaad6ec63b07b04ff89e7d82b5211dcaa257e67a96a8fd57534e7ea200319ccaf3a8310de25ab91906a50aa19072b09f31a9ad794cad3749ccaf5e013874d2dfad6e7b21b9f63ed2d13cb2ad8beb162d97fd5493f9796428f9bc202c5af6da4e70e1ddae0a1dcff422c48069eb8f9c154002af7bb0eed122f55216abbfbc61cdc9330df2dc7d18a4466dc2e3643de87a08d6120fa43d3b36341d85c0897153ea71df4b9c7d5dc7ef607b4bf856782fcc08560a7ff57be0bec30deff23c2cbf22ffe9148394e5e481acb1915e53d42564169860c3ae83ceee2b3a6cf42d48c9e34e06b09ef40b5b1f63c2d1f89b62a69d39ca387f2347d73755abb19e0d28bdc2101b274cd760ece870af800f1663b241b26867c55a1385aded140e6709195d51cfd2862454d48b751ba088310fc48541767a17cdcd064cf23a4d9eee2968726044bd3f1444506f3f2a7c0801d09921b07ea899bf21f424b831e4e2c5dccbe8dba790403f69065a68ca574fd5c134a0468cef32c8e8a8846c43e8c942a7be9e366fb3fb9d0acf2a71513c88154d9f0cf84b9e080e327a6011ec5373507128b2a1b2ef5d041ed7fdfbe8964d2328e02461d46b4493fbaee3b336bde19170e2fa3fa9fe769ca5c41b2f059c427200963f1b4b2a6d5c70269b67ef7ab1822c2fae50e25c01a2a30b838d8ee43c2bc27b89b8aed3b6de501c32feedb1155fa26e6439311d29bd9a7bea4b57d3bd90ccb872335e508dbc0d95108cdeee08aac6b3205bb82a6b9b4464f76af240739313d63a6cec422a8095a1a1e04bacfdd71957f71e0435656112ac1711f981a129e456b04b4eacf5e850ec02818676c04949d7e0589eee4e00bb5328a6f8bfd5677bb7c71cfb14a0e8028befda5ae186ba242dd292951297fe9c0a14673b55dabb8887888d1dd1a6a777ebda21a63c0fd1f5a96008540d629fca84b0f5498c3a722f6c85d71b1d1ebb450d43362f878166b4483eb415f6346545eecf8fbd88e5c31b59533a4fe987ad039889f075ad0f32eed37e6d5153e5e5953c759dfccd8129fe16f0681d3619a2e1f32ecbaf26a2e80037c61be52159ac29b7da7ad8a9f261d33726ec70524c79e84694a6bd367175b8fabfc49e9b8d058cdcf7c91337a3dccdd4de21b67b7e085c6ab083c32dcc0fcc7ee01db7f018d440f95e0629bb2a5ca212941e02f20ff4c157f835d83ba71f24efe39e434fded6e58ad8bead088717b378312ae977b63766d0a38a551a8580494f60a7fe230666141e761f9365763fbf7e467c8dee717c35a9d6dfade0710ad58dce8ce615c28dc237543066923bce4030dbf251b47fb8cbca1da8a034973cf426d932215552198c1624d85edeacc851a0b2df411903a23f60e1691bda4fb1782e16c96f622f9064c12ad93e5ad4a65b10daa93215bf2c15320e16529f66ceaef0650d8d8d140a8dcb7b2546f8e52986250c1d0da26ab86bf5de2717ee3759f3df1e5ce8a7300de4770cc7e1063578e9b94f7f560dd036598a2302f205b4eda7738a3e8a12b81f12187d7131a43fd891ecf83bfcf7c04937f245fc6d385d170defe312321ad941d0f7df9e1897618959e310cd03661a280f62fb3c45efab3a0170bc71db36b4026380137807c0d6981802c3d5247aafb75d58198507e6edd07e771faadd861cb92c1d1b1b58e6d9ac906c10839aefeac7faa5414d2c81fe4640abc32ee8a0f944682ffd4b9e70b1a7299ea343392e73e67b1a11b36f0dae469b9514dc81798de54fbedf1bf6e353533f1956c6a7675979a74318e3c6919dcbf646820265f311ed64e49e7b7bafdd6889fad1629b79c88cef987e55355b97d57fac922a400432ca53609751572596efa0c38ebec085fc1e0e0bf0e84e2f9bfe120397a3dec639a1428f4e4336c227fc6c3f1838aad74cdfa05106744ffdc8d395e8ba75fbad3c926132bd7745bd6e01103badf33aa3af13e29c92764de5dcfe617ae3c945883cff2a4668216c0b76c550d7b983c50b55fd3411f747ec7b7a36d2a0027ad442aea4d776275e91f39c4990b624141cfbeb382c3a590273086a9b1a627668eeb4b2341ac81809b78c799bc529a53cfa9f23296c457747d26d4e27ed8687aa585f8b71bc74a79131dbeda00cc63493e95dcd0f5ed98ea7aaec5bb54d4a5723458f6dfeac0388e11689ce82c6c18a59845bc3f387d913b67490f8872819b35a539d58678891d6db26c6622a0d0b860f1830a1cef55bf0f5cd1040656cac8c97e7d3c7bab5f381f1b90b41d68bf8a33ef5046675b55649fedb7885670ae8fa06a2b2b05d502aba3e203b4c23bddb4b987d07c56f934b70e28839e0d758e4e6404f17485701abfb1cc8aeaabbc2d9dcf93005099db1bd345d61df6c5b90bf2d27e417227e3595d47474697b5980f5c82cc16065d7d3d96a77ceffaf5f06c4fa7cbb1b2627f1f75ca1ac934490fba1d665bbcffd7c108556ad7f55172e98bddb553afd61f723acca325211c7c2467ceb627b0a2bd4e9ae5ad62213e05940db3c125244b3c01c6feb7137fd56e90c307141178af5f7b119be0bc733d3739ac2e6d9c0b70765ca49d9166badc2c67b0de5365e9c43b8712839867384115c9de65007e1c864a5859af6939cccfed0edf9a499e9f5c49b3c0593bf505ac2d1d70dd0209a85c296324bd47fccbbf0cb75f35af1a9e455528ad3fad734e596ae8fb568329b1efcab01529fdb1f9fcc58f6a125c3e24fc185184d7d8d886fb1cf992673116254e67d85b8ee5aefc5e8501c99212b9c3d624982ca8aee427432e744ca407a53d5b57a3623a31df9783f9ef3dd3ffa20417261fea06eb3b95a2d604b1e415421973fe95f6db1f0b50b04707182cfed82df8ba97367130d1f102f7b0c14834c5af0933080c0b622d1866e1585bc1f3faac2cd6ae6713b4d337f14b6331341bfa598ca1d1e32e7d6e5aa6046051ea8c2e42fbd141d17ba5be5319e4c57821f0e1c01c828b70019cf2bc143c16d14d6315c8e2f9fa1e80532d85cc15f098cce13ccd91984a081498f60be6c2ee1f43d7d12261491db682bd2d40caa73373d329dfac2947fd37ba90d6de48dd7f3359f2fe729616274047de31269ff3483134236809a4ab5aa25f7261ec24004e0328119c53db213ed8743505efbf96b2698b83716ab0690b3f03af47905206cc2e45057964c413eb356326954147fef891fab462d7b4ebba04f3394572eeb7aafcf06aecd7d32b4e460cc1bee041ced81b80b7d698c20e3f36a767450419892e02555cb8a4dad6eff073ce5fa3d60502739f25d76f8025cd85c7026a200793d1773a507a382e147e994f88adafdacfe0c6dc3cd5e7634bb82ff9c2642fa62bde4616d0cae230133500dd994930ca76002e59205a095692d634ebb0f1830b8db58ef9b4bcbf2836bb786b49ccd73bdd944845565b5552854a14222886796bca5f734071f56e3a641d5acc1eefdc5c19ab3d75d11c1d065c2b39491c380bea4cef3534f01619ec2677ef5d23e62e4086e725143098dce63d8eef6bb24599ec996c287cc29348f85697c803a9845a63e1013d71d46c58c99deecd9f71abbe039adb25d7c4f1914be30a7d99b280256d2c7653bd9dc6c566092e4c25426af6f584ab8868f7d287fee524d014c0d308e7c85dc1e6bc17c9cfa82420863af189242b21060190d08000e610e05347818555c66b68207ec3b5b33880cf1607986b0f90a2e7b6985f9b6617e175aa8540ceec52d2c9ba47bbf867af2dd7838e3e649fb6ffd2a727b8b2a4984bae3372d26f30e8455caa829a8e17d895cf02d598844cbb00f7d53ce93d4be677ec361927289c118a62680449c6990cb228cd7ea91243071ed5b070e7f989eadc16e9c135256ed74a4ba75a8bf0413735fafef852490365529e4b4b98f40e5a2430e2ca7b50d94c738dd40879e0ce3c349e695130723e67d1af0913ba92fba7531b6eb37fa5a8f8c1b58fb710582f0fd1985528735a6acff1cf0a1dc8ab21648b813d63dab57ec51ad42a167aa385c8576f5e2434948609357fab3ae52c5aa9ee0805164a07b221ba537a4377b4bc7fae8f6d6d61a94348d21dff6b65ebac306f76d4bd0f5d30ffe6794301fec9766e71b8a36329b162484ee4ba4d6cf27fd597e9d86838ea81885f6899212d264f2f8f4f8b0fd2619bdb31509894004ad1a14bf890c3db9c783137c163aad71023988436b8fc483a8d281bbe0e20aa825ee79d1f884512f61320b233c84eedaf4306193710d1a0926172b1b19b98b9f05a0e3867850aab57438d904989276a7a070123be1bf4fb337b75c178ead3251185d4d1dca71d494884e5562544238ae7c63efa675d6924147c3b46e6e261aaa26e7993b7b16f629539e3bd8298901c5f0c938123efd3528cb7cd46cf74b3439e6882a1830c0427f9a4dbd10b1c722fb1769445fd12f18fdc27cf67dfe7370efc0f8f607f72327aebbf1f4f034dab6d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc79bea23a6b8697e550d0fcd97f6d5a3be3f8fdf83c9918bf9047896347a28b9d4ca2a85f7e94b000255f1f2fd16a228e745d870d7be46dc9b6658845264d8351b4eb68efcaeb7b658517d2b00b1f5a2467276940688d4900fbe9dfd57b32a9086230d565249a0a7a7f53eebce4475a78941529af97058d29fcec7c1be395ab189527d9de2dde5258911b33ac21505d3d94977f036a3c0d7bb5b6e504ed6ceccba3d68d6a1c9766a655bf99702d83b0a18cef894bf1ad7ceb5d96d12a797fde08d4c018d0001ec7a3a14fb380f1907f7ccfbc014da91710b02e1ce2b423ff044cb4a58a6045d460062ce62e7d1abbc8810e15e28358034247524fa70c375086bfb828e0c7c59ab5f7282f78c652ad324a4ddf44ca6d76cc0602575dd1f69f9f679840a311923f543bfc7b93b98ce85ab7e75a4b39aa0cfab0b180689110740b7f7867e0ecbf08a88ef83d976008de3311f4579f4ad62e15f3468065635c4ec5913b5c9f03a4083ccd1fce5e9ac33554dcc5871c469658d7e1efa79736adf2871bce68c921debc7b7b6282ffac2eac9aefc9119b9fe2e45fd16d771620e2feb80c67029dde1a605be384e7a56d55d69e783c9b3a29aa26674209b254786f9265e2457c09306d8dd57357224d13dc01c09f3a93d31b960cee7c5875607c99a8decbf4eb2abb07b8847b19333a61f31ea7f112e56491410af44273d466a05e5483aa8d38f4bcf7a9c2df21791793c04cb68fbe76ca99d368115eff222ea15457af06ff9437769024e85222a3da8e732a92451c8f14274fedc33e8f84e554647467340d0b9a0a40edc10c10ed6ec04606ef3d7cc7e27296bb0c8d951cef9b1a172946e5c27c4eeb5875ef5fd2b1d31100a857b8c1470afb37cf15e59fdd4491a7b2f6dae541e27900e4a439ce7abd7a9a2391cb9ea220498325cafbb7c24b36c2b4f9de4245e3d6f7805f3d48ccf74fc45f88c04aa4050a17e55083a0bb80f7e7600e6bf1029d4020927b05ef20a78698de7f7670126e7e6f64f6fa9d78af80b7fb06892c230a75ba7022dec0fb1356530bfafac6a5d127b17023550a13692cecf8c4971007307b7c1fce73515ef061f7eff6083cf28f8ba92c30cbf3726c8faa5b1bfbc201584be4bf88a8a09a7c359581aeee33c800f314a8369bc0225a40c7a8f4fcadd88734f83b63afde79fb02649680d1ffc6248d353b6d2a9f3316913648b5f1a3d604f17834208c74813f0b2f45d0a37da6dd53eaed83cc1fb4587ad86c776c7f158fab63d6468dc1f6eadd6cc3f8cf3e694a67847a5488e557d0a6d30ae1cfc81b92392284e9c896bff797e90407ff03b68e70e55d77d501ff8bc8085c3d086dfbc571e16725653b26cbc8b85700477d2dd7478b66a89f00608fc5b424d8bdcb02a246946f05fe37df0ec621890de3d2bd18007eeb228585e41a1e6e29b69ad96a50d363e70bf3b89990188469cca730bf07b8878cfb06953c5e4a03108089acd4baa1324aa49fe6b530feeda69c5a68c779f2f71c71a6225d5b25db0218eb4e9deaec800cab3217b6cec5e2b45eea34835f557cbbbafab8d6f1c6cfc1e110d6f47df82540e97a36fa5e9a794774e4010ef53b6b22b64a35d8dab044468e349fbcf592a3f1858b413d95776f112f9f0675e0d2babb274ab8cdaeeae7c5738614056451ee55f0a30e5f1124abdb4c95bbac35850bca9b32bebd96a1e34bdbc8ee2a60c83006fa29f77f0af840148f5f5ebb53f2f92c6c96b510c96f7cedc5c1d87b769be88e7f426c57b399c3b226c108392716862d904bcd6859b1740601c20e84c943f3d99253fa437d6246fe8f623520d293b33ad6e28b415357b14faae59fe6e1e0954d2db8d529728090a9961f17314103c2d906659c1c302622ca04ff691e5b4ac2be2e2bb752e3541fd7147a33a997989e17ca3d79c6f92d70e680abd8db1ac604f556897d542bbe0ca42c28e79776bc93fcff431914d235f18cbfa49e573fcda916ad79d3837ae3c0aa9967a37356dd1763601266f53dfe3b5f02dc66092d47ed14820d041c382990d126edfb167c7ac1f5782faf4c5f8ddcd0ff6c1bcff80d1801e09a20195a654abeb3c3a7e2ad3c704992f9ad23da3534e61e1630fc664679586c20fba766fc02d41b4e0e0e9e2d2f77ddcec3f99ac0fdd7f00a846525b4e4168ab676dcebac66f0e25b12c7b2d1cb27ad191ad9e4e98b6651063efef4a1f72df25c601b4ba245b9dd3bc691e1da5cd68e763dc7a514636cd508dc4c6403714800bfa93eb7682411f3dfeaa468e8b6638fabb213854ed77f822e8b730930797bd24286481876f3b1c6d82dabeee34d842b4ec9de9c43a0ba8a18b6663f91f0ab363046480aefaf6bb542aedbb3258e91d9ed51a02c21ac62daaafe29e6e402f3a39adb866ac6a68b3628ea6764107ab6e04dc290d47c349191585cd5b254a4880e0b7c3211cbfe8fe01aee3cd9ea4b057a3ec74c3df49b164dedf7a6b03ae40c58c50a595fc4e212582673f92aba189adcec514cac1db111818e71833006530fdcc0e2c93ce79ac2cd644e8161d38ea130c8b1c0af7c64a73d7a19e11e51a96853601cc81ed5a90c9affa10360bf4f5d5f0a0dfd3002eef11e6c23e8954b5bbf553bfea1f22391260a678ab65635e826be66d2d7a2c54396e50aed867a0c7d68dc2e6b28f8b28801fb107a63438e85243f104cfb8460d501dcf67fc010babe534413bc550fff306b10db0a76a4deca7bfea54bd86792988f56b0a6b7303d783daee54cdda2ca29ed02be370a45d39e0b2624d0de636e601d08321c9a2adcaf4f2c551acb2417c3f733e0e68122e420a346b49c82d512cfd6756a8a962b0860b133fb1ae06bc1f9cd6f5fc9fed0c410dff3679750332a5ef9f9228b7bdff49bcbed5c878a1b4af8763786d22ebe9325ea81b584221ac476692085d949709c55ca611f8671afa96705df7148d8a4ac64806c0a4efaa88e2090478603d7f1861edc163d0971ba6d34104f6fb7b196eec4f9d75379ae2bcd8ac67c311e281b1b2cc54ce84b1ed4adff1d496fc2ef697ff8ad32a0eba50602066a182d864a0b7043c250049b84c6af4b388a06c05e7817378ced79a9d9d75b499fed16e54035ea0645c368e861693e6bee6d3d0c30d2843b29e2a0b1e93f35cfc26768f4f65136d75217d476186aa2e8b3ebe25703b491f7d21554c062c6fefd241b75cc379bed3869f5f6775fe792b16860523e920bdb1518b2f95c7b6f2618d70629777bf204eeee8022c3bf1d1d245091b6be1cddc0f9bff18354ecb0131286075d707e5c7adfdf937ebdf3a54b559777acf76755e6129fa2bfc8075f69467e6adc2189115feb35cca22ed0aa34b8d0756e2fd42a2f69d1bebaf4ab00331817ee8e1d96a0ff2dc3944aa4f9c010074de6c6a847fc0cec8af4c18783c505c141432f2963583d137842f770bcca7836a3f9b9ec8de6b66f2594f438dab274e52ea794e36e378cc67e89670bb9c10d06b6c1a41049ee0f72054d64885fa6e306992ffcf4d03d94eeeb82c62060bb075e956826757f5f1c4098b5d3fdc298775aa0c8a2cec571431ccea3a0974813d7fb849597f8d82e66f49d9095e84ff37e3d1f5063e6eb4922a0c0f603a22680a67862c9d72c3032a0432e388039bfb78233136d3a0ecacd192c53d98f8e37d48d42d760a6cf589522b25151abeab6c6e91f95834773e60bf2271fce6d3c63497803465543003a966882cf2cca5aa02d7ca2277e4adfd2748e6553125432a20be867a833605f1e5b94ee06b87ad07289258c98e40934cea56e3a38ca915df2d41f0ab2236827ff675d8dd9f681bcd8be366b91e1bd585b795506d63872019d4e88509c1fa987086b3d75b232113535226d961e36d4e4917b4527a3df54c10eea0351e82fc45f1f5373bf6d77f72fcff541c5e797d691175bd3fc7b27b30dcda93647de2a16ae3d70c720d9df9074b109d76b7501595030e10b2e01a9fdd67fe8b214840fa3cb8e1e95aaa4c9e3d2c28c398fbc47dfafe6b817a8c67d9166d01c2288b64ba683d5cdbc742544a3cf4e0080c5805594e63d00a2305bd60a9ddae652cde39c895e739beed002746dff24928bce11a3e83fa4c05490374423a1bd6bec85af044f954b6cb52cd0546c4e5f09129171759c3695089d6ffc1328920e5439e446aee5ec5d51d40aa87fda6b7b3f0d96e20c603e39a210a063d3f527e306c4be6bcc502f3833023b67bafd1d240e257e9272cde4a947ac3254d3f40c9255415edb5e68cfac6ad1a73567d0c216e028f304bf44f50b838e5c016e8e1c30dcf2217d8c84b12060b30085d63b74841ac3696d97fffa4103db282f147662eaa8a8a99609e09359acffd8a09118525f2c26ac7df222fab5d3666f65db099b072194af71e0541a10893604539eec01dcd416da4dc85ee5d09333302bc4a0fc4c20a9cd8b836dcd63f3cc991844137bc7db666727e7bff03330afb2edbdc2ccfd2348e600b7ac29012f237fe69cc63308c75824e93625053bb6d9e4c7ac27fc3c8f9bbd9841e60dfe0c124d6715d099523fb69e87cb31fdb416d4554da84570bfc47ab94587b9fdfcee08d9b8e506823f563bacf28fe0aee4329e0d3b8b01ae29865807926ebe5485a632c3a0c248cc8a6443a5a2957c0dc6689e24bbee94849beec33b63c595e86ae69475272e607e881aa4442c7fb83e7f49ed8000a5928bdf8b70ecd648f42616c2fdb351d740ec48c1adcff975ca980322f6f3a945432a20bc6402b9f903b36347ddd87d4e27bf16784357fa8ee58ae19c1b9e066707eed49e0e2157f83b569e8d3629ff1c6b9e7c60313a0e505c2553597fc4087db980dafbef33221ebd3263c70af30c3a0e8131c997a542a6783517c739945fc2e6b45fc72e9e44dcf84c51089235fd8846455511dc46f612f079bffb5b2b08e644d4870e69321377db9952a545b7b049af2e1c59b4b4e55f074d6787b3c28e9d382bd29610314675bbbc2449fbe4d1ce6432ecfdeb093869a86bcc4e02c96b8f781c7af97d4d789ab9c55b9735ecf5ec8ef0388d6dc471aa354d886a365e74ba3e384a26e287cfb4fbca5a3922e77775d24c997cee5d392f8a1c451d6757dca086bac1c96904f259f3f5ebf155dc3c57a1141e24ddb734eb66fc7cce79b88541cd61c561e4d6cc232636bfa1b4b3b9cb2239e2a49bca1030f353bf15860c49f8978ce9580682d5b253fc07a3359fcd01dda76cffb4fc5b9be5f2fd57776fa3f39515658879293d6d0c381b3d10a3b0c77fd05b69e6693bec2e2212955f8e143c4d4cb0a539b631979907acfc47bf7822d77cd2a8b8b3c9272dc1c639f54451236f4901b0f0dc76e48649a6f94db76e0508cc212590f891fb0bc2f6e9660057ffda9ffec2e5026b5382d42aae1c7402f4094de7ae94c54886b3b30aa907a83d2e482c68f7790f061e0aaabcba06b41eade2e5c7faa8c941435f4d7245e9a97b509163a97da549d7fdb3e01814af03dc8e4736e4298fc8814011b3ac3bdee26b121723b9c1a247087ef3a06ebae7b650fa2ab22a8791e68b4f0e7341b4c618ea05606026fa092b9902c44e8ab0083ff838f84c095e82ee9be69d13846a1e4fc5d48b034f48e3550a163f4e71be38a2e5f39a79e7c438696e14404ccf5d42e3858f89deda30a88281512b38dbecc9bbd107459184dec6770445e24851f2ee5471612a818b0b594fb393879248535ac0f3a8462151f2b0a4b0e0769f4e4d96ebf8274668cf278e22ae6fa753efe2755d9547b05294d92baa5f2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7c73f79b991f38b490b9891b3382df69beb12ca55a4d4c4396e26b5fd0857adaf6bf839d5dad68947c4e7eb7755f5cff60e9552e98cfaa6b7061d32d96e6750f843ef5dfa681a6420a07b145b81f1fc1a2b755ecd1f1754563972b99f95ff8671c8724d0bdc24dd4e02459dab48a7445868b042a93763525347fb0d066cfa765701d81b431134b48dc9e4a9c8b36c878433b6ca0905207973405bb6dbc98810c4a5bd6e35cef9a448e5981da937f6164cd215a42749fdbbf737d06f66c7007bb90a6e0935074d78f92684106a45c3ec175a9052d5f6ebda3b18a4f049f66a00aa86fc168225a764965276cbea19dfee61741d3d33025a839c29458df55d01a0c69c4c8bf829f1bf141de3f6d6e525b00057526fc5d18478438292cc68a24e9a9a15b6d5c3163e1f6d7ed861d55852424429273666f4c6e3e9db17b915e82ca8822d3d1de7cf7b82e93476b5b3932f028dd8a655ca9fff75342b56a5aa1c6864ac05cb69f4805608a5cfc70cb8e3df24b3f4ec7c5bcd411d421c6edf948c7106c52bdc459f74dbc87456ed1b163701117084d1485f6e76c85e5afe0a04c095a8c33f988f3b32310211688a6aa1c59e3c734b56639e9f91660cd44f3b53eabb4f4044c9bf9bf882a16a0d324d80278dd7d6ae7ffda2d3d8e5b0db4c8ca1f69f0152fee67add91bd9e14c900b53b11e3adc1f6ac69ab03c23b121d2067eadab3e0287c5ecdb1584e7121d50df79db671eb98060d4c6c827da2875de39290e5f61305431a8cb732f1246af3b493a7d518f1732a450df772c80039c2fc68b81df1a391269dd98842c9c4e9a35fc661841ba5da77dedb49c8d9b04429bc00243e8a2f2540e61c550202db3a33b7a32e52d1d004abaae8f2741cc475bc411eec57280b2c9047fe5ef51093cbdd8203525a2f29e753f3efcab2f20c06d533098f7d079aea11f0aa3981e5014c76c0b165abd8a75b724a0beda5eda3c6c8e02bc58bb6eb1753845a6ffd4d11510e1f6c140b4f57fd75f3c743734758a6ed2c0e7f49508dd9c6a6b367edf0f8418cda92072af20db5f4ec5eaeca8d4f9c434285e1c99e3795b63ee2ffa3f2d05ab008e5d8bf0b3f4821c91245f1a4e624a901c00dd29a23d222add481b3a22d1cedc8c49a134fdbdba956a95e14a028a0760d272b09a49bd742fc912f9565b3009422b641be7f590fe7e4f7c3aad72fa8be115f17eb16febebfe15e52898b7e746b0b01551dfb7049a30f8e73727be71911b089fa17ca813b50fcab7b40d5f088103372414fb8f5fab32176549038ccbc51f1a02b6333696b0793f477f4331cb3d32bb2ddb2ccb81bf59cb40834028c166a63f915e41d8b75ed3fc8cddec8714049cf466bac0e7a2d3752fcc6a5250067aa883209327a49ce6ada8ac5f64c49a5b22f71318eff303fa3f89ea4f1842c1023bcdf3111c4976a624ceac78efd4fc93a692913626156fe2f2740f9ebcb0be6431c8424acef961dfef1ed3ce97bd59b5f939e509fcf4916910c75b045a59b92826d202c01ea0376d89784d2dbe4e9409502a7e8fb9a642b45d759e4b9dc2b682da605e46294fc2b161935f236bd0f2190552bbf1b5c5c24393a4081e5428a4a1640e8637a33923792c821746a4ef5eb3fa1e08137288fc58b32a06d5c992aaa8137267f276985b1e92dfc4e41b09ccaa6f88490d95527641ca32dd9fb6e37c2c7793a4168e2eeaf80e1e3024e60d6d2d74fb6d77bf0c6a5fc8b939c9739a66acce53a2052928ca57d277adcefcb46d90830b2e650cba49df1f703867a3c9c9700a3b8c93910e1d50691ac7531aa776b1d3ba2ba6ff230403ef44879af26fa011ad4fdcb085191bc514aadfe3c6db2a56ca18a6e60829e0c67ace7490433ef95e2d0d198019c0382fb884e0ae564d935568345041af06c6129b4526359cc7a2f2eb1d6244d4b7f9c4d894f2ebac3445bcb4956b93d6353f020de1383a68240b2a9d5e34d1bf0570b2d2342ad3af9834c3df61c29e5bcafb82702b4be65743abaf12a0cb5c0d85415aba72253b317c8a202a06df4afbd6a1917f59e66168ab7ffa6e1ccef27872918637fdea5e81957852e80efbca964891694aec6a6d97ea77d30864f9c4cb52e72d78ccae1cff116ca75d02f1d3fccfd64fab7194dae08715ed2a968d0f21e5500e0af7d75a66d17b23b1f19e69b504663fbbe511c50dbd93ef33e529290e3ba47c21ed0d8a69f893bdf92b2fd3e854b752774bd698370d4c5c846b6f633f5859491c31146d0a74b9e5afa95c08ef53e8c237ffff53e24c6161f460fec178ce7a9215792889a0d70b6911c0e473022d9d2594c36b555f456a84b6468475a280cdac8c898fced7df127c349ed3a0dbe9475281fbd30df9d5498f75030dbf2dbb9a26619290ce68777e284fd9f5529c659766aa409af3c0abe714a629f040ae2e8c7a036c70e7f0f83d36fb961f55863fc9aba88d3bda74c9c64d722b2e00a701dcce9755e945e324c82ec977ef66371f390fb015a57b95e9db9115d0764a7b2109a615dae34b14f80ad241b2029534afdbe68d7c710b402cffe119458eaa27783f8cebe20bbdebbf85ce4cdeb4dbca6412a0fd3be44d8d68b35933f18d644edd5afe2e479f2c02bd6f955194b0a2b48c823f9c1ce8a3b7ada1412634769f003f70912f9a00a94004f64e9bc4a774a67d244d8095971275785cec16a6118d414f904e0a3892c225b0b8526e32dfb98bc510a12072587cac7ad4d768229068b989f8ac9498bcbf2f6a05127fd44dc14d8665751a7f63f374f027ce4c34d7e6b460630b6aeddec4b14e7bb6b17dd589a57c270774f818b1598dea8433a5efc3a00d12aaa42b5d85570f1bb06099bee2643a9cd76ac45faf19bea73d666646baae671d393d52de0c4954b1ded5955d6e450e71efbd6cedea3edab66533f812ef1df0f50acbb32e00c1e4c0ffc2de7eff4152a41d171069b1062a130786f6745506e6e656250f4e35f9737a18b805fbbdd4607df4b4003931143d30fae743bd9076a147856b6650e05d6c57ff5bd40ac903c2456981abee7dd166a69082f0d087848e56b9fa4b2b89ba85a3f32e2a553b0e791a5d485c47d584a1561781716fc508c4397c1c4a2b15ccd4b2d89d90c0308e70b95e8e4877001f88ca0a1e25d15bcaf0f7b3fbb58be87317e8953a13aa6bd9bd8d1d0ba7220f73edd5b122d793583d5e627f9f07d43614d3e84f831331963c4434341da1ff743dce7abc5463bb389dd6c0c85b74eeb7777bcfdba70d2999396d332da861b9aa777d4b3ef67e377201750354a386025c57e9616202b8586d1b77e0ce16ab60053c2afab5914048c1d5b1034019c0ef1780a0d585f800e4a8d84b4d8a1d5d2a1a8cb717226161873a4b3b3c177e82dc1c9f554b699ff412085aefddfd3c32499b1682a0208c1106e5c7d02b7e9842cce890ba717c61817952e570796387034d0dd56df0b69b673a5e98e3a474e1279cdc711e42da9cdbc2595ad54b2fab9f0df87fcff8aa8fcdcc1262235440240cbdc8fd8cd13ca055226421d9bc5643ec10383e37f703f60cda503aeafeb525f21afebcdd446c71272fb624f9fc280ca4c3eb709ee98fa478140c0d9915fc9806d37ad9be9b24471908f545d77951f78e013bee1696e2e77ffd3aee893a323fe68c8afff0045d2925ff2cc2e342da4d82a803af8569accc90ee6714a1fd8bfb6d934b6b6d8e46077ee54ca38450b55370112b14eb648594069519f0784ade599445aaf5bcfa0140e8232ae6a15f156c1ea749271c7fd8b856b51a2c96269e7ae93a8453030ffab1c9422e3d6f8288c4f34e13bd3873ff4b30806ba8e7520da6471ca0533c0a9b8d9cdea3a9257a0f8978a8b00e6b8bb399bee9aed11ffab0f73957e0da882038f72fc0a6c5ccfe6007abc4012626c406f42059a704987284d73e37c0002d6fbd3ee72501e69a6f5fce664f4162880a65945bd40117fa1a2785a1c3f2ea20c92d3d77a567df3798afafa480edd003ac07acd11303d6c9f1b61037ede9ac67536245be05ffa6f224cce10853d307c3236f6f315e9c195a1deb1d98977edc9dc9680185eb314b80198112749a99b242cdff8c2cd75969d584a0864e3418d077e5f7b8617bc0570c4127043cf22fa4c73ee0603fa36f01c0cfd985ad9a6fa05da91d2a272fdcf89be11c4df5a00e1e6386ec85caa1a6084a3bbc83480b3ed2887896edcab8c9a26a4433d802b6cb5b26fd90c71619d479d5026f3e0b15ba0a9a36a4a2e7647fa24a51c521829d8831f52f563bdcf8e91f72655c27a2f305d090449a1d502a5d34cabfc85ff95a0187fd434877ba91bf2a383410b708c4c1b81e9c30b5a6c1aa17dff9f3effb46931fdaa871d2673b08d8157a28619f00b85739b7f3e4c4f234fa814ca243ea86a93eb12700ca098bdbfcba20d6b07510fd292b6c55d4cc5329c51d4b3773f7c05ec5b53bf67b559be8c5f5f139be04df4feab8e24713406d2d04929040cd77c3b78bc23992455d401bc7cc941303b6f78177149dfcb2361c98f9cab188dfe0f048c07e5099d6c3572234036fe9fc54978e0ff75e73099163b7802a5949751031e614417e6e49b2020ab590b2cbd5b2079f7b0b997690c5073a04b7e4195c481cadf0fffc6c5887b52cbcd359049a5078782345481f6e3f1b423395b11169df1998bee9f9ba1e8be07440b2e04b0a443879503a18e5e534cee527aaf7b4e880811c6f58fb8dba21dbd5fccc23226dd70ae4cc97bc9127a9dae5ff1a876b2a417612eef9840060d7a44e10abc1bf5f7a76e09fe2a2d92df019e8807f1ef43d5be98a608c7ead177ebede5dee7767bfc1fde84cf7e316e03b2fb8275725249b0bbe687c8aa2a131f5d99aff4882ecc11d71955d2f5eb7355e16b52a0b89e9e4e9d8b5fd63270d3cfd663cde8430596b6e21820263a74c6988d0f62dabc17f9678cb02d3b1be6a543dfe5f88dccd85fa30c3e530fed02023dcc26ba426b18c28e21a4aded8a42c027d818aa865045444f6317e7c2d4ede4f7ec71b9d5e458f8b6735d6e040132a9343361a1bfed6e8bf785314a6e797543dbf820b1c3b21d9a3b422ed6c44962aad37f6167d7d1a4d590a9e4b40e9f56000eaf2e0f6fb9a15052193c536ab34856bae9de368f030ddc3159a26b08421cae892c75125e27904a70e33ee5351333dc7aef2706405a39d3e8a8357f7dc7c5441da1c1dc5ad618721cf6437b5f916fc50f6ade6a93fcf36d43f3570f63c259644fd931d8c41c016e288cb9e922f8754b9c9170eaf7f9273654bf3a05b3ebdb47638e99e0bbf12ad20523212e3c73e133ffc9367beebe70805d2ca65051603587fb9e5f93ddf41ffc837929c760263e2bd4694e951f4542f8c9b6f82c41110ec5865ff2e09304f0fdaff5c718a102ff84d4926c7729036ea1ab75970566281419adb991d807dba64554ef93aeca34359a0a0c068f40a519ff652c375b07c0a49a7abb2e1ab71408179721e110400c23bbe40d06554dd9353b0f366da965863592a2f97ebc2ae584f89d1cab0d75ed020c794162269d252420a85d7cc1819479b90a49134efbfa5a18e27fbdd8959a2e34395e9ce10322e7b8d15883a7928f50f708e0be4112c28a476543f53ecc3d4bafd95ff275d85331646e2ba34a6b3bc4cdddfaef42e68d14f1789caec42f2b5d88bddc306a85212c77ea050c30f6c2da3ca925d55793236ddbd2b877798aa0232d454235b7d0ffc24691dd57cdc25c954d939721a88f42da33555b5c3147617ccd5fd1edcc993fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8aca33818f0d1d52df0263786519ce8ffebcd924de0a2f3ac2380e130bb39de814f18fa400b6cad507d2d38794423b13aa919349ab1afc26f0c510e8ea28049bbaba13500f6f5b56db2b58f8097c86320c4b26c2a5a5114e226e96d90d99e2bbea60f1e065ff6551bf7dd557c6c336ce4a5253ec420f081ef3572d9d7281926faf6701247d4bbb92039de61c2e39f075e6bd60a5adee240900b34b3eb3443db0de23dc5467d0315404f8703e5940c9fbf5863d8a5e9f16ae97967f92a0f7481aea870d9978b11bb753973caf941a070a4e0d3b4216f02643d7dfccc80cc32f6b44f82c0c04b23bf0c23be8944028c93bf41b2e0fcfa941a60164c30c416ace8526c76a50267eb9060d177f074ec42495d48eb4ba23451483f5d7fd189025062db255fd3ffc90478ac3e5252ecf34c607845ea0747256b6cb87064ba4ed790dafd8016e75430860952047c12a0f4af2b327ccc3e5666d1093a540d02e7d641a7730d6aaaea91b865fc0873cb91a8ba85fd82f721c13007ff7cadca0f1218eeea04efe8fb5512ff8909eb18c3e31b547faec761dc40f51ca85f96a3cea0df1277a678a29c020fc8d19d5fb188bad7ec434849681f7ef7b3febf14c0232d2cdd4732e8f3338de211f6098f880d451567f8f6b10ada63fc26134454677a6d4b907d5a857ba10c86034d262e91da2a428d2c87d893b6f2e337582671ffb333265d992da1085ab5496e5403a66d913adcdcd60b8ea8e87c85ee5bd90483d78524d0b67ce711d1bf682387dc528d319b08675df75567ab729b4d0d128cfcb6545fb000fce5828619c2ec0600da12ff70ed0ae4a0a2bbebe6157dbaca46931024218c8ca6b6e63e83e2f523b1c81d567b1251a445d0dcdc559aa81c52621330e8ead8e7ca5e4e666dda452d12735b742bc62d26db4083d0ae7202e0e5bcfac09a1bf0061681d325272c3fc6575ef1dd160737e993be51f141ac834105d9e5cee9361bbe4d4836e57d94c32b34f88db070817b97886e480675594c0cbbedef3c93987528fb4187d3b82b2d50665bb5e877bf2ca775be06d46f8ad917073f9bd85cff7b6aa90f41e8e22ee5d9f7927869f34f2c96d61629335370e3fa9e45b333de089f342fc02125bc02730c837f08fefb90eeec5af95324533eef668e8d87ef210c203babfb81a74fae90353ad12ea88f48101704d5ab1b0cf19729d47928f6ac6b95f8c077cb82e741941d0f1a33cee455040686c2bfb18535110dc29224ea3cc183f3fb3562dfbd4b01a62c23d5663777578de6a2ecbea85c145a8a0537c011570247822696f1b41ab7aab8dea8f9908168d567de0fc92c8e16310e90a79fa87359afeb498cd8cb8e999c1cc49d617407daa504116f9b10936096d19a964966c672ef071c2e98e0971dce2e4aeab38b9d395d66d9833d1cf91ed87997dfaf7b60e0fa3608a86f9b251b4db2041d624373a1f09e94ff1b22eaecff22f775f8732238a37cafb65c10e714b324cb4a3fa1e1cca5fb4ea3d6e1957f1b5eac23a1f2dbce9c4e996d8fea3578dd98d41e10fa4a5dc10b36e7340eaa8105a67cc248987fc8677c20de064d41706295e9b53e072af655aeb069d72833bc0b99224557a995e5104b2f3c7054bf488f2a72c2797530d34f2b1da51732d83be9935c0abf8d9c173b24fc94b8d6607a501bcd32912c49ed5bc800b4abe22020a80f0f6aee2e71405ae658942ac4a411baf8e3b36e9fdd2c79ff243aa18b8ed7cc16aed11432e7715b1e72d46b4cbac89a6fa544433c61b478e8227e18421e43d52b88aa44233b8b08b577b82f50570f7fc1027b9138c1b5040520e60168de893ca7120c5d368869c5b55a942119c95792fce174c4e930232f77972d8ec9fb3cb81e1180f9aaad7643bc0b5b89738d148f92fa0b6ec8791282c20afc77293b04ab266eb835d7d7c6b3262510f3091c9b853dd4526f8d1eb735dfeb93a3cc0a4c3d05ff6a78ff9b9e482ae6397c3365dc7e229e0aee955a86527af868c0316c10569f06de7819960d9701a02e122a1e1bfa65905cbfc32a49f379e4d8a50166e5faaa836e27e71726f2065ef7693f51e999730e3247374081a5ed6faec3b7039c8ab9e021142ef2db5aa8ce8aa9836a0b22541f7b6c864a6d1a62918a6cb3c63b0cf281083aadfb7287fbaab1eaac66ea4a9250e87a9b6603927067eb262a4977170269bc1d1c4381151c96a16059f4cd6b0b42aa34f9db16db51f0c36e0db7b03783d946d64407dd21e0ba5994e2662ab8fbb3b486770ae5e151827fdc4a3cf415372d9961f4c2abccfe62bbb173962252ba28a59a4640aeb4f35cd6a4205af31dfb52716e7b98e206d7f54d9b5997e82258826d051c61aa36bdfa212e4506f98036fa3f75f6383b1114bc248feac363c42dac70995f456ffb1d3aa1a36ad7a01ee7e7edf56c5c1585ce61538c85476703705a08a53f3344c343ed387fb89cf0ec811d29bcbc7b068bfead11f112698d65e1ee1dd3454b924fbdc0727ed63ddf431de9aca0c18513b6f2e40ac1f29239079f40ba1b05f9d3806162998c25f0fdb65cf3b17f7bfc596db56e4efbf1e32e4154868a69e74d5951d561dc60f5a609d3261377bfa1d6b521a3879c34f47d108017d4cb4fc096a362f234b80bd081752788c1d5170070b93c1451f16781f9fef0d33fdc41453438b638f6658967939b4da524495a987eb7bb671ea8b6ab05ac0a40b3ee20edd38948553d7b45ecfe14a2aaf244fb1de41a32ff0f7cbaadca23a97d8b71db632533831dbb8ee8cc23265a82b4f1c0f0680491aa2df3ba77ceade92a99f4a3381b3fd87533cf20327c448f89796909fa27e9a2654de9b71d4cf8179ae93913b5e2a3f7f4f05d07119f9a86eca4b363992db8f5076fc49d341d4bc41c029d40965b4a7fbc632d7767ad076b4e50b5ce28a17826f469374bda4a460fe97045668b8ad3cc491d392584f9db06412b4fff14a666946f3f39553af3ef2f9ccdf30cb9724f06a5c1f64ab887f87816a2d24b3bbe3bba10508038baf751f3db2183f614d426bf94c2a3b7cce025c3c5d6a58cff77d0dc2234b9b638e2b8388e239ca247243b780f73ac64a174764841299f6602ae0a12d9a95cb0420558315d6256758d6134f2b99be70180bdf7b438e9842c3f2b626eb22cabe402d1054802873cbfcf3ee798b7255f3a51ad35723ea6b859be09f146b2b1717200db75090cb6e06dca94902795703e2f56137b57b8e829bd0b109e1fe4b9e6a05c36a2269a52f5aa406ba4bd5811947c0c1e04b74519defcc7f9e6dcf72f08bfc370234103ec3c8b797a3e42f862c4d3721a29749a6d18ff5ffe219c6e20dfe40f8f9ffc2f9f0850fb7d9b97231d6ff0468e5024fe4f15b6bebbfd7319a18025ea7e76677b1d729133696c7418420bf793afd67d0c343b7a78e85f3db17d5c2ca394b4ba3dfc5bf8ab4a1a507930a2e03127d279e3cd162cdb1a36d2c4232db08cb072a6578782aa73928ff34499f7b766002d37584616879cc4aebf327944516aef62b7d403eaca4f00398dfaf3e6c3c9cd9b41c9e50235a3f444fc6d99e7643760ea3a745bdf28bb6a1918626c94c35abac5d3dd134f176724b2271cfa8cb8aa04cf037ac4ff7319cd4bec601e0a1d93b2277b1ae00061cd7af6d4c870691f3cc72114b6e7f7eb2dc84a99169ba37706128ead6b41ef7f180c46ac4c8fc4dfc3814e941a2ce356319e988109f517d5c777fc1b41e2495f687fd0ee4fa54bf7ddc0bda43d9e6eb62b0f2cbaf0e2156ac356908ac7fa6400a769518262609de103ec7d357dc0d187d7e7bc80c1e709a3e420317a640eb3a92e238f2082654bb587cbc86f5c7dcc1e17ef08d8944d230cd002ee8bf730fbe448373146fcfb6534768f7b24b8855a94d76f22d199537670493efd7b3547d3c083e62d4fae9936f53df184b689f70787770ad6e3b522804b9be17d0220fa6d64483c9fbce4a7d84a0ad723e4cf8e3d28b8b9ad381d1362b2232ad585fd8bf22ad5109a6e5fc5cf5bed43475ea6d0d286a6d4d99362f28a8e17a89567d5c299a2a86e3b72012ba1d21b0175b529cc068ba8ab42379021c754133136c223da79261a9439469fe1e2aabd4cd2e82810fa22d714cfb7954a06425605641cc298e71ebaf69f9ee795e8326d091154cba6016f1cb573fcb06f1f0ee73ca584d3eda1b93e67fb55a44be4f1e7398f337bdac080b1c859b62e0d60e8c8424710bc364496c3cc488e645f6bd738d2e3dfe250f18c3f7d093de92632f1aac4786f8761d50942803e9b3f346157f3f587e01015a495f55b5c5428b347bf751d45df8dde91c9c638d69a6eed2ace964f8b059b5f923873c4bd92a9b070a640e775d36146681ebcdede803f3c3678a0d472b622add56f187c6d84b661e1eca835cacac3efaf045ff19288645861f79647f0e2aadd44371b975fee06e78652d2eda85844576f5592d7446452fcd5a1f6b1078dcf6dab43f879a0dacc39c80fe34c7440d4415f3ae3196f776573f42143d6f8c5001fcb356f4a1d98c1b5f78a2d19153ffd5c5e53320e25fcb52c649941ed0300e764f625892e87fda41eb1a1fb06dc40afd185a588ca3299466e4d1e989dac16bd277e4c3ec4985b8594fc509039e5a2f40a9b8a2bb538aab64a2dc931ab774eb6799b1ea286300925f993a5ab695e7eb8c410b72fc8e56647bf4b4238b1d0ba8c2091cdda125ee2308fa31c249e181066b8bd93fae2c78d07b26bc3cae89b3a3faf3f5903cda3f765881522ef4495aa662f93229d7cb407fbf1149c8951b3bd257d2ad80c5282adcdef6b31207abe6f248d2fa670736948cf5818673cdfcb46cb790773f998a82a4b74e8fb3229d16afad49f1f8c27fc22149d79ecf16d517451e6acc78347fea63d698b698af984e582053f01008197c0e813c793f893b33530ff78fdace08adf5b0c32e44c6c72896585691c467f710cebb7cbf961427a8442d96dd9af746d9ecc69c9c3bf46aef517f4d651a102e19bff09fd5bfbaab964c5500c0da333d3400373534accf93326b8a2e3f66692e14ab23d64ff47b494a7e26432984a5f0b22b9b6cbe25e91718250258a939009a81114e596a2f0bf78451e245fb363a99a41fbd25dcfe1a809dbc2dff7d5e78a37c652b388224bdc0bbc84ad8889467f6aab1a4c60be24173156369609d0f0c3f65bd0df4be25ca795855b19250ea6058d9d0a7fa36b3331cf21569c715cd06c3f46a370eeb6498353e7e0b8ebfd79bc070d385af519fb5af2848b8f31d38322fb2b5f8d3a342f5116e63a95e406d7085ee80e9928e434160261d276fbcd7353dad2a62674143595b65495f0594406bd9a477d76e1ef9bcd3f290653af80bc300bbe9678af099c85ac56902a5df1eee2813f466cbd41e96db8e958ce434770a4a30159d126e2c46e6b80d6bea5dfac03604b54fe0cf0ff540d6776f3af11aa99a5e7881b4e6c4efa83a46c8351fa3187fbcc251eb99cdbdd92bf4f8288c9ec2709fcfe73f11a86c3edea7e8deace853cc167471bb2add0206ed87315fb49b5201dad87d5ee8011c421a2894f7761140341de41c36af7ba3f753715e7c6f13bc11b15d31448213ece0e242e9087bd50670b2ab251873afea01e38a7280eabdd1fef0f30f3cb83793e8025d06d266c5f59cb789a5003090c66d7225926d62c849fbc920bb1f6221cafa61fa01f7d3e27a47c2e3d27c21af46ebe39d2b86c12d32410753995207a322e3d14ad3ec8b8bef584941087e2134ac74af9ffc1b0b414574172c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbb83ab552b5d5d8d51a3171f78b94462ca67a6fa1a051d446710139edbc365026e6b8a155a8ba7c68f39cce0ae1ce8054cdfda20f762ed0df9f389958bd15aa61b7ca31d70b8947cfaa68396eda42ee22355068d2113755a83654a74549f083718938fa1481cdd89d29533d63a7bbae6049d87da3a5a08699ea1dc307b87a0e5a5ed0be7148f0e86daf059c281186bdbbff777054a32bc4155f81658b5ac3eebcc289f6cf772b1f718f57e237320dee0c6d2125737efcd72b14e258ede41f444a30c99d96859b8400a580ab32712795bd5c19cb46d2221eb6da75e6a579c6301dbfabeb7671c7350180b3e20d44e51e8c1a367a6aa125c02dbb3d3e9783fef541bc51e8948e31d87853c9871298669d045df50468dd00c79754a85a83907a6cbebb8ba0607710ae83a4443818b30462d527807bb609ed4e9757e3f69d76bc99a49ca42817593ac4c57f026bb6bd4f7fcea9cec5c9acbec225c19ebfc1da9394eaa9b33b956bf7a7d19a9ca66a0f62755f6547de58e425926a8f7cb5271c9555295ae04b5bd83718d7ac5558118b909523c40b7044a5079a048209531a8ad7ea24184b98418fd4606b4ddf9b830899704c166c09479f9bdc997feb74c3e26f21e922ab70144826207ba6976fc7534d2cd3767e08524b5201dc1c23add924c5e7f923115cc7282e65ea0c035603e49ffc1c4ad4eab2939f7fe8ba9c5f17ec6fe6eee9e17d00d03f6450d62a1be81517f5f4327747d5f2a9f9e74dcb9f25a2fab87ba444d2ea9fa4d8da3b2532ed6e7518cdd33d983d4d96bb5a417d8ed8ea32fc0e93b1c4697ea9e929e23c14e3b3e62d89bc7a031bb8d948efad0bc5dfba3fc3c87afc637d7b4ac78934c260528aa1958f998a9434b31ba4cf8b0930633690793944df97a6ccbd3d826fce2ee738834e8d457ea461fe90bcee6c89d7f3bc967010fa5f1246617148a6e4c5676cd9c9cdbcf6a9349ac98d29183e3affd2c07e61282e6a4ecffea02d8b5cad2da115af7465be4febffd9f180cd465bb9019af6efd5c9700fbd68b56d9a6393c8fb94f2fef9ba6bd3bfeaa5465d5642f0ab7d00d134e380200f97dd439a4d67f8dbbf56af8b17e399bd622f48d7a7091afe7808d2e36b4eeb0f16c5a62ec4126a6b64caa86c3ce233dc04f06bbf27690782495db9f0bf83074ab9792e5a1e28755e7aade51c0725fe0668354bb0c1d8e9ce064c8e15803af88db14af9fcd2faf744d6a40fc231a8acd436d96e4ac6ea5073b7321df5541389e012fd9763ca71c2ac37992796936a999a1dedc636a64e9ef80ae552e196477d92dfd1f2dcae9b38557e2985fa27497482e294ae6060cd5dcf673da74270a88e11673d1f1b10add6a731208c0453fa33ceed987b39d1a97432c8e5fa89de4b04c8b057366166ab2267023e7490480487515727404423d3a2b84bed8805f84a00e8ad0dc059ee5ef415fae3333e458f7af4c6fed400ccfeb3442ca91283073775ffcdabebcd124a11617509c2a0340b0b3ac60c32fb778a3e495ce75ab61a1967767891c9319fa1560bb8ab8231618f46514fb110516aaa0e853a6e783014223eaac3c36a1e30daaa2a624baebec276c6d8a4f787055a54bb97c0b4575ca93867d7752da30366300dad0e6ea04808d5f16c9137bfbb8b2f741ad347aeb733a9ce5fb9ffdf67ade8c8d994b2d421f610d19ac899215627bbc16532d82bc54ed5176c96e83dca6987bffce6eb3b441cf1599513fadd3d34edfe9085e936b512bfbf104429a631a11767a2e1d87ed5167c08233a1b6d7f0abba49ddf360b78746a8e46653f8ca705eceae78da125389e97626c7ee34fe719b0e992fad9a5e29d5b52e94dd93f4cb81054d957ec93a9d9429e1850981146de1a50fd53ed4b38854b62edeb7c75d8901c54b07fab45d3bfaecb09c1946fbcbef52f596e282d0540b5a9ee4470d37c24193eeab213b1b499f8b25bf3749ccb6ca56e453c8df3dc307f7a02d8902359b41f18695372a2188f7146dbac1e3a5e684de913b0aca57c6f638d9d21f65fe9ab713082e2aeaffe61607a0ba7c3b59436ba4302a3188096f7f87bbd578db6958e9556df504222dbef9348258690d1713830d81e8d2de4385d3e1f8b7f30d7fc5ffe5169290ac7deca703970acd72cb236d0e40f28cfffe1e47294d6f0f1fb310d0cf100723a80c795a00913ce60542a134058bb8bd7904e590dd5960b435f48b1654d0374b52102fcb0d87876cb76ead8d46b551a976be4955c515de04c765b29e11b6a89f9baa33b8682b70df4ecc19db8a701fecfdcff60c8b92b20bb995d2b3e76a5fafe547e9241aed2c290ed63c39380bfa7f604c3c2a10be6ece56c42a6fb24db4b014da41fbdb255530c611768428ecf47cf9b250d7c4e8f7324246c42e34e1e05822e9e6b2d557a74eae768a83016766b3986201d09dd06bff991e49131bd4819c2a05fe2a1eb91dd4266dcfcec469a1ac4b82d3aabf98e767bdf356026f98768deded335eb2df7c10460287aafe78f6a1f50b2556e51f95d5650c91e476f016ace7b008152945ad68c5364f5d4d48c3c4cad705a6ddc0fd2a69f49e46c97137dd41e64cdbe032bd73962dbe51b58a9079ef73def80df471e0d69e03fc2e95e9f5d26cc94066b8d24bbd0d881877e0f8f0d4a31af67a7424edadcb2dbaa3d1873bb0aeff3d191c929777e9fba86911f302a6f360a93952f5abf99748fb13ffed7350253aededfbb0cc9c04f1a50b4db486828337d68139edefaf2809cdeeb0e190105b5042e5c4ec3a4d3e3743fa38d5986791481d8e85f0c0f5ebd553ec45eac516805c5c118eec9acebd47e712e04d7b0bfb53b8c89210f5a3d306e27c5a13b97b64641cbf36b51fe1ecde74451c745b5544c4690cdd7d5e60f24fe66d5f601003fd275a18838de28eacacd45e82a7712a1ef8fad7530b60b054651b2d39407aff8a7ddb36e214a89defa30181c7c21b6e3e00d0b4caf269429fd540ec7df103ad8e0fe8fa8f3eb91d72d59f93abb25476c64989ea68c65e6c92c2b1e75380916061e409d82d3ee51a4fa37364e4520134402a7deb2403f7198734b1442886a1870b7d60cff7821e5c3174646ab73123386bc85f65fb12a7e9074eda6b00257e517ce09940d5504e2cec9bb8d13135abaa461ec0379eacf6fe9df9b4b87ad3851d3bc2c4dc14d73a350f0de755d460c9520270a5aca4de9eea28e05e23a3cc7907a46173794223e90dc7dc06399740d76bb869d8a7dc6aa2772e164e9d39e300fb488eedfce63f47f4810eea04a561025cc5a2b20392260b21ac8deecb2d482ca89884c9486c40380b8d75d863d4c20f51d2ac1d6a68bd5b94b23535e90670b5d38e8412af910a286db0b5cd3c24e25d7129afdb917f625a3358ba11b61ac16d36c042f30abe8e79e1398a7ed1c9c11e43203d23926490208091b8e4ca18a674aa0476a1a740499f476dd0de06c329b0dc6bd3f3139c54cb6a504d33c727e3206abeb1772dc91de18c9fe91e8fee72c24094c61a11089eaa497f0f62083e3ff1afb161620d53ac921fb51289e8b96e0a0bd2d27a18fccdb04e7ae85f2fbe54555079f3c26d9dbd2068405ba97e9f8dff82f3b8aefbe886e019cc8417e0198164c67e3341738687593ed1ec60a5d2ab400fd9365438305b833224aa72acb69e308ba9f58d4f43638dd8a2b04b5a785f3538d744b78394d0afb7e0df7689fa48dea1e0269928ba10fecaf5eacb6c0cc698c296de5c07869ce7ae6b2f41e2e75bd64b026f6d77654c96a2fcd5395eda3ee61b0f45a5e49183bb6140d1f9c6c47e6763d68c4c88a0bc4dd45a6172b14102c5fef4208000c6006884197fcfa33757883711a13a146272c55be1e4015832d783786a4ff278e827bfe9edf0059138690428ee70f3607087939e215835b0ff881cae65104715e8d9da1eaa391b671526bd518a4e25010ee0a12e4a841fe435d3b22e471d8face72da6264d9845fa646c52971af63adcd8b9a98bea4a6a55af572ead325b4de9c12f513720cac2c8b569840e960fabe76ddb2fe4ba18f3288f53127433ce14176617c2289aedc20376ae3a594dbb760e106d848214ea9fbffccbf039fc07adc68255e7c6597093e414582085eb9685a1aa58c772a4bf428269012f0708848a8962d15e5c613b3ab840eabdfd5527a30f22f9172b40f2be7e98d1350578994659a8445e36347620e9107871bd82647b5e2ec0dec7bcf6013a81154bbbf6456946716317d7b11745cea71f1c8596b7b91f8e34af5e53074a5a124d34bf4bc4ca501f3be8d2f2b620b42543d9e1f0586893c7f0f33b10610e3d3d8bf953a4d357247db37f9cc85f0cafae6088eecdc64ca5d0b83900da62300cf6616d2442b67ea7dac3cb1c3caaf10b7d80d79357a6e57d808d012bf40e18094f1a24c4d370bb19743dfc8438c370f344552e1ea8b15f75452ea90903331fb2189827f717baa642dc6cf69e8ec03ddedbdfe21365cb9b7f9aa82ab4498d2181cd8f6df3780fc1b0ac602af2bf85c3ae4fb3f5190aa79e12819f75e9730cee46888da0f81e5137ab612ebc7394140451f282772b1e5e4d677665f7f4a768af9b49f39b77843f5797bce719530c0939cb4cf099777570b6e71c02cebbd2d98a17b8de5c45c1ee588f80649dbe801fa99c4e7fab3b6b2a4354099ec11a2a62f4e7face13c9c6f3b9bd88b8e983d18c18a24429dfe04e2bcb6fa1f2937d54846ab7c9b44e7c9f591569738da7109a93c50c184ecd4df0a1c60d1a3c1411dc25b31b6bac1fe52ce2892558f9c24cbdaa9689c692e645dc464c79e9ca52d2962b515c9f426119a94f2b8fe778ad472562196d661b9534867f90cb2957101137210d1947b52bae3d9d0044d8da87975d9ff1252b88351847ad1362dc649d22deb05de4fe702ac1a0fa04a0e8e48f00c3d92dd5befce098665a11f556a5c52cc3a802d3cf15e92e5671ae56894aaca8b40fadbf00ccf509994d80e54e5683de9ad75155759a8af8db6a1ea03b379320bbc450ff38cd260572f5f98686afa4c5aaa210118499e74825301180c7c865fe9205c3f2c032e59c35ea45691f69e2b720ca81a731baf2a65d85482e7f536e634fd943961701496f2d3adf836d1ae1d641ca3e2a2dfa6340599a72d9ed3531dee1975bf843d41ebf6823e19b5cc94484121d51f6f5eb9dbd0b0c8eb4bb5f851a0cb780995c6acb28d2756a4fc89ce99b20a6778e3a5eecdc2f665e7a733125ef501da34abdda19d366d43e24a2732ca82713588a51ece8fdd5ff0df068e590fb743778bc69593765fa630f4cd89496e185e5f92cf3694fb4ed077170ac299cbeeb0a82beb7329d54cb2419a6463e8d20018aba103a10c8d1d1c27affed972f0afd66c294c4b1e4b4bb04283a682acc8e9cf2fe98e8a20732c2cf85b9d9d4ea533c90f28b3312092e7e6fceaa00374777d335e6cfd28586f52d9620b7f88800ce141d3d9b57bb88c36f374191074894ef04ffcc7839efc65b235134d14a6bcd236d75df9d034efdc406f8aa3aeeabb2cd42469968338c4737ff7c0ecccc9fdf3a29222364265d81ba9bb7bdceae598d61ed7bc57a7e2e46ef9e69b679a8427aa1c56d08bcb5c6ad753d0715c2cdc95c5c88126e94c8665c65aadc1720144256f78802c59f3dfc099222651ef07d42b956aa3ee839c3b583b66b439296c7a0325d4396bb234fed62094a1427a7ad1ebe0266454d57d3de7cf31accd9c13edd3e5db8feb263e8c56537e8ffa08b8da08cad253bb4ee08bbb04977;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h630737354ecc22645a82a522e906fe0f1a9e206d9d91f1e910e9855b32805df5fed502f38ea07917dbd86f23b7f4d1c45eadde4346f809ccc9b2aaefd1837686805f2725313cf46e1f6ea979c720fc64141dee5bfa65f088bdf1a352f86a7977dbf132072ca218050f39ca94dec4144f0e08f88e498026bff028da0e94404319b87d04c20c326ff88cea1dac00226d29bf97ccdf7627ee918b1e206f830868d97eabaa512080e1d120a535b2e9c6386f1acdddeffa88cb8be7fe7988c8dc756f6ea25be9d43de25413f8d98cd2a21be6648ec2fbe1b53d393d2ce3e4b9deadfea12cffe69364ba4a441531e0b7e6567e29ea577689c5d9444db50d03c7537fa625fe51cdc59bfeb4df71809cd8de56733b252859f52b1ad275de13ccfe9c94304c39735b9c306b2f4d931088a61d8389de28f081d96cbb892408a79a69a30a603dc3b23a089edcddf4061ce448419c45257703a93b8ea9ff16cd888da5803a571ea222fda5577dbc6d23386f0f31b5d45d5b79b60c35f1f9bbb89d2b0d257a22541fa2965d331b2fcaa5b354ce900aece4b1965812a723df108e38a189b89787f2b1f82f5586e73064828617896b03a158291ed28866fc20f886055885a6451b80476d420d3cd244e88e788ac7c506dc61f1776c31c28b4ee7b62939ccb9481803d684511b4f4944f008fa107c51196b06302d51813ad9c38d7a1c15ea1b2d06e8ad4c1cc0fe731fb7820cefddbc4b9944c67fa37a25f456008862799c2c1a5e2a18e706fb79d1d0ff0a8f8817bda80a433c91b38c01e0d6c8d3cf678da1019e8df5ea807e5386fd5a77ea01d2963ebb72696cb236f9f051875b024a3a2d16750a85c49ceb712ce4c68bb141e2cdae0beea27c6abe4b70909b7818f6fbe72a361299ea19d41e374cd87e2d0138e28b07bd8884e91c1353795a341e83867afe60d2a8306411c4f156033da3162ea9ee8bf4505dbdcb5d033280aba709b3dc8d973a5e2702076b7b47f41b9b2577f7e32ba63d42c1341ce983a2c352a918258bde1dcf83be956c0efb12399b18df98f8dec05c7dfde126b0e70624374ee0c06d58fda883d8b3de6240503fdc067c478d8789c2d6038e43c9807dc3a25db953f027bc7aacdd149763eb64e599831603539f6ec2c558da3a5c14af1170e4667c2c80b2ebe74b452d05a46aec7319ff164a28ea5b690f12371a8d38f60313f9b0820682873a326ae57a3da7822302a94b721c1a06c213e0740638e967bc2e7b3dea34c79dabf3404f5455e2954ff43aff598f538e1288302168c7a4cc1fc259e53c94b35ded8b969e60c8290094223b4dc8ba31d969039e8359571e27478ef11b54d37d3339fafcdbf010cd21a90b618cd6a93545072149dbdd079f6d60350350ba30bc53bbb646f9c4d9da521aa52821f78b97b0c19b90ff41f87c4138177a411184b85fc84297cdf7796f025c7f86788db920c361ef22d6c4cc9e7c6b2c9771d7bc1eeee34528d6ea927945076cf86bc8da786a57995223be33009ab523acd34fab501884b1b562a04b12fd3d77ebdf81f44aa110d895750e8688a0197fd3ad3bd2ff672bbcf3c5c69ac8dcbbcf7c5ff93727994425e5e55a119c95ebc0a123268a53942d364cf5c5117d1d09bb8785aee05fc2bacda7b8171f9c8b71171f64de2d5ee645b0dc697d841dd8de42d42649e10f0c1da63dd3bc4c5bf50f36789f09b39a01664b8bacb5201366c9572f766122645fed334a7826d2d3c5658da771e58dd09df1676f150759d55714d047e5d16a7a29c391ff66494d2329115a5966f7676ceffe63e6a9af5c4417139d74e1779d8614de48a12a0f5cde67b3f912203fced018d2e6652a72ee38c5896861faf39c44f4d41ff51d1887b54951b4e0f7b9e060e769a71956ab637b61a6ff9313feb5331952ec0dd29b43d147e27c4339304b46936c2ee616f572a2a5a2858618778057337e617a32500f8dc8b554b8ffb58098e57a1f2cf2835a9873aa72af3d019fa97491c0b7f1e77e0b7a3615587c53f30d89493a091d2d70d55d1b739c6fd269d53f4fed2c6c6428f58bf3691a7247e632d2ed1f74ae81aab2b09d41ac9c532a7d98d03a4cf63b9718ac863d88f70b1a7b8f936b1931b542d0a604642b4fe5fd54487664aa3901372cff3f3a5b0717da1309d8c196cb616201dcd3b426d421b751b2afb47d14ae869328dabaeee41877624a1984b1d10477af4db28dbe7ae3fac1961e6c257eac5b1897f0d0fad40fcb076b311f8ac4d11548b7b0a57faa7afec012cb1fe47d1a584a6efc5de20d0d6660e28213d1c309112e9d26c9d51cb3aa76ca48e834a56edff7fbfdaeedcb94ba0d58ce55ec472c11d39cb9a7df39f914005811f217daa9b39d1cfd6109eb2ab667109e0e30397eb85659468bfa99e7782ba484fae5dd71ac5e95d268ff01534521b45265cdeea6db85cfb216978fad4683a941ee3420830112daa021da4ddaeeb5ca190d92ed2e0a416bc39312670507139dd37d04c40ffb6ca7db3b437c6fc6d2ecba95eafa4c70998ae23f8e1b63c661969dcc1dc7e2727366e198c3df2c4734983e8799667ebf5cea30b068712f969a972154e355b2683e1023faae76bcd46ff041cec2253502d5b22d76c989ae4460ae4704bda19b7503308a3f3bf6be1e97ddfad9a205ce711810a907a7d9aef2b9650a01cfe801b4c1601003ab092c78dc1359b2908cca98d03bc533282c0517f331641be0e2cd8b7797d433f677ac91425b8590e189a2dd8040ff7c397b0c7afedd3972083054f1a2c08b542c6608b16dd166749ab94b49e1510d4c421b8e6f72ed46ca0413e7df45c05065645251b9675b2e53038b4a85bbb26971b648a79b94d52b5a6fe853adabeb28303aa68d8ed3cfd4c42664215c3e19c5fa6c70b63a4adc3e5dd42cacde27d36ffef99975ad27dee67919d6ab071bf6b5dee432ddeaea2bc369b0519ccefa2ebce00cadc2c0eb1d3120ea71889b84c23de1cd1fafc0f985eb72b524c43731586a073a298838b95c5605b9505bd4a4d3cc108ab4bd7c2219f82b0d497f51cde8322992a42c0e43fbd9608fa4e1a73ee35122e8e71734bd7d70e44eb8317bc60dbca951809f97ae78b4c59183c486a982acdd7d4a2993b913f1dcda2f19a4bc6663716fd15717cfb3d92e7b736ee98eecc6889b4a3c4cbde27d5bca3a9564bcfa8375907f7b1013560854f0e0152e3ce384e5b24b447798b5a85b72e4ee9eba034853786f18adcfcfc461744d23f2e06f165f726a09d7a0892abb0452664dc5fd4eb89fc0c944cb6ee23a32c7c805386d22d63b7ac305333277b662ce08e02fde5a757867faeb250b3edf1dfb83b19ef2bab616953b13830ae82ccd515406ef3adc7018d90dbb743a3ae6c256242e97c691520424c3b5e4c4cc8a94e6ab462e8478a3c504778d6b5b6831e28f632f7e750250ac6b9f2d69f25c9c7008bfcf587eb1a0fdb93822b7f1d6ee304ab0f01e4d854f31d4006062d6c21eadae087d7e093b17cdd0027d6abccd5684df462c027bdee04a70a95363ab05da80b5a231f260726474cf40ecaac89f26a0d044f1653a38211391bf9f8005fe9af956b09e2595992f24ab625bf9530b772b7ff96a18c950b6f3d627041fbe8189028c7bb0420c9ebadb8dbc13454fa566972565f360c268c27b1c8d65bf5663533b178eca3fb6fe003051fb611b9fc4a24930ff007b8ecf46c4252aae81338e93a47f6680c82fd1d5cc4e0ee490507562f349321385b4b7c9fd2c605fb61a7cba2d9a92bdebd134c79ac99236e2045ac41204a341442bc3aa5d83df234583e190e696d4ac26638fe8a1ed2172de5ca224c97cbcc46c9117e0eb9c57fad6f152700564b04f276551575661897f9e1c895976b45cdc7d1e82a57510e09f48c98b033c4d454ad18d91b7a1a62813116ae2d61046d62bc961145359e1acc7e7033a7306faa018a7dd107a3848f3eabd1bc3e94224125a65266d0820d9a47cff0aa37a8014c2d33d2bbbbcfeb936a3df58b521984cbe759ebe932d68c6bc9e3b0bea0872d4e5d38771c62959f99c97ea7177c051e532afba977c74fd7525b8e93d2be2fee9d064978af0824b95ce3473b5e29933cd0a1d0c8c2098139af47e7fe56336107be301041b682d3bff023abddf90b419f729c02d82aaf2e344b6fb91836108f460454dc957ca61548f1267958257953ab50e0e380894a3e3a934af9fb224a911b9c3b59b8ffbbef0b667624d5eb83e2d5bd5cdefe7711116ad4a4468bb58a19ac5b7fb69c5ae80144ba5e520958bfcf4557a66a902079c9538c4d01eadd94294d83413845aff339bf3b51cdcf549c51f559db9b0de5334a645731d65f979226787aac5f1133d318426e0aeec489b8ef60b313694d9594cc6c2e50230158b866c1a16f6ff88dae945a4c68112ab640dec8e548a008d5e2fc459e09c0edf21723066c582bd6a021a944c7dd515eb9926654e4de91adb920d886db127b62c0f4a22cf812f172d898981dbdbe6c4a1b0242c8961ea6a322aac9f0dd28692a191e56e58ede7e5cd410112b620ed3c66086cfd1da787d579201c550df386d693f4ed74641d16dc42cc537c1e93d71c9a6a010a45e11a8da60209942ec4661ccc06879698c2837b4f6e0ff84a1328738b94d946e160fb466fe4be5a3b9b54a299b810245c7704e7ea6c9c6e7fae24ba45cdd5ba84a965c697e95192aed87087a3ed84560b62af7740e196fdebe3f2e33c2f61ca2371cb9b322d67affc34fa3cdfe4219ad7fec7310ccf0f834dc4fa438a9b2f4de765ddf474fb6d968b2886b1cf8bbcb6f26292ca88cb6c43984859d8eb4a94a8d73b9860195f288273fc6549b579f4f2bb5ca573fcf66095a2a35b6d77b2ce6e6a1d2629a03b9b092207fc6b258264f1ff64430d164b0a461694480a603874d6fef241a56c29f8f838d1067bff9a0e90606cf200ba36ee4dbc6beeab25e7f205ed6d63ec2a8169367ccc2a3384459ee0a39c3023bd396581e654de0631af48210934d12ee5e26363714418ee98ccc3e8f20a6a2021cb94805c66ab13aeab3cde5b1ab0cebab610783ad235ffe13ed62526db29938976b981f01736dc55df1dcb50f918c24313c5798c00b80f2cbde7d4d7ddf4572f2636e10d60a9f0d6682b97bb92bca34371478e367ff357b42f0052fe4222a661cca4e0e45df41e9efb4e953c1c124b408fc5711929db3684448d8935bdd53b7ad9d5bcc2bc3a250e54f3aea092487d06ac1de3392c7067b5f8c23a52bfed4953d2ad2192ac46f04a36e263cd426df15b7fd68cb453464ba605ee230565fc147fda57eec17a1a5d354c565a05fc894094b7283202de75e0aee2a258ee5d37c25853f2829242f5a1bc1b85e25079ea74a4bbaf5fdb45f5765b811393b26e4a16fb4571d63ae38e996a2a635f7e61456d0fae24821c83cdc0e8c84519a5439ef33e51ed326acdc5f431da1dd47c4e8863614b613da52d4c10ac841af9f92cf0a8cb3ac4b527370d9e9e2a4af6b1584364e1c20591b027bf295bbe0207227925af253b98c5d65e6023610ad09380ab0eacb0f15eec123436ead021e89447130b1fb2ac1f9117037fb2750cd1ed19ad38367c62eac307e863da29099c8f8a402aebd0e26e78f5d3c7fec9e04ab7400026168f15fb67b2e819b78ac5df3808d8103515857b52b4f4c55f32232d74d6f729d32a71228d73ca74b6fd8a0ea5963ec0e9316ae94cea8a3cd3c41a33b01c73848df0e08d8ad81c37af38b734eb9ff33b5a6bc81b1c791b8b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb8c741f2ecafe831bb43190855fd9286b0d45843f26f1b5d8620feedd8deb80d9f7d8f418b414b7e3204cca361696a1313a8c9b2ed109dd5470a937a95a03f902b8db07b92530caaf53d33b3a4cf6626baf88693a016f2d5db764eed4be108da341db3e307637470a7541628d8464f0238807fa8d0d0c52f5d38cce2f12ac3512fca71dd2f228a10301800308d803feda662c2e5f02cc47979a0ad92967d530d551f25a3da007f2b3d8e7266bd4d264707701b1434680c450c87098b91666335151055c8b293418526ee5b71f49f47271430f456a9dfa31686c4bb64c23db8fa54a2fa228162c58fecf49162a13c284e3c51b92ee082d245a2b5f0eed98fafb9e41bcf3f735ce922cfe805b5feae6a11c2f61e89c51c238ca5f66bdb0ac4baab85715c6775da69523e80876732435440893c0f4a493c027e819be2493e3113d6e4f7f5c9955354c0dde2c840f76b3e278732a0e6791b5c317421e8df44ce12576c274a1ca0dc301397e9013e68bc47d53828b0303b8288862976b03a3fdf87db7b77458e2859e389b3b4892ae5827a12bef6320e446d84f5d0fb1cb02c4874b4c56d5f3abb713f517dad8bc140bb31d6a832ca0609276717ebc7b211dece5de505fa00d817fbd0aede1915bb2f555ae6ec63fedbcc870c0f9f7ce1d3ef36ad82543a87ebd3fd2e0ea176181b9b9280135da85e8f48072222606919df133ec5745e3f500ebb673b822152df1c93ba77780251a97b6ed03d603d4b0333f874e2ccbeaa669ab775bbe195c22f7074427e5817afff16df577687c0fbe58d130cdb69b7c1fbd04b5a4c5ca33136a414e2dfa5e329eb6969b1e98d8861cdbf781a37cabd7eb3c6045ee9a83803aad5d91c19307e28cef8864bf4c255ebbd55ed35e79b8f3c414091ea8fb1c21a8f6bd684fde70273f8365ad5a6cfda3d34895f26ab2a5931dd1ea4906d4149b0bf9ed5d1b0a9321427e2aa8ee16e45bca14c9bddf081d13425c243671536fa6282dd83e2571065d6714ce133023ec887ec50625482f8cceb6f919acff71d7e5cf690617b0765781a4c0ce222756f0da3ed7fdf7936dcdd1c04d95012535914f8adf50951567bd0275b76fd4d2ef298732fe6eeca44c27b188160d369bef2d75d5f8b5bc0368cb5132b97052b56df826b4c4b13197db4746b47f419260985e3a821fd4323b9ed6537d7ea3291347d1198670835cbf75cc850642b0ad37b3c98e0f76480433baea163dadbe577b490378a22d417e7ce478e7cbf55ae251fb3856c18b16ac4db58a2bb8659abf8f47c5d1d3f4b6382b0f68477e46b024c7e781e72f0337663db12817e15c768dd4fdb3bfd779760344986080ffe419fd699e5bc126b5192a0ba8d81bbe052037a4df5bb2e483871575430cbd621ce28c3023c04212c849b864693a0dd1e556096de60442e7e11f960a47e6fb5bdb43426a4cc4beee61914acc82f7544a18ce33b0ee0a8b5e624a22f4a06b0eb511bc3bbefb6879e2e89f7fd1714cfeed04de6b85cae33bfb495b31f101f7a8c2819a37eaa823f3682e621186b133a6f8ef04d052b0b038ea224520c67c98b8589e814a88e8c396e1b8462fb4c62157b7d993d8603a26bac1d6559328f1eb14a3f39a8db79bfe193f598cca45ac2fb2d26cddc36d4e3107a090f7975a58af086ee0b100fd5e3b71f509fa36ff4f869b0e292333f691c5e7992f1a418bd2715f032ef01f9567248b6fb6f2851b83e4114ffc476cc6a3af9c8ba92d771fe2d5c8bbd278555de0cb5056a7b9b7820962c22979c73abfa3abed2859c1b10ed25d42950f9282154fcb74489f9d1156b24378db6bc3c14b1e5d5a237d0a26392e2afab7f86f6d7efadff50b920dcf62aa3022f27261ce2b23c782ec535315b6d85fc4303b6580224e91471b8a164c2b1fe85d2ade36692bcc1eba6f981800a6bc377cc775d87c733726e2e8234da32e1b4ecd55c98db50915ce083521cd16369feb2c3b412b6aed9aacd98bab433708cb3bd9f598bd12e5411411dd6c94c06dd1e0e19a06f07b83f2ccf614a1b703358b846cd1aca8bbe782469aae5fb3fe2090b0a8c24d787ee149d223e8b3316c618a704f473a3de3ce48082d3c7d33b1f829a3cfb1253963e59dd6b5b5425108f8c1ef06d3b86499121094f7388cdafbedf05ac34d52f5521c73d1972661ba455f3411f5f79de7c9fe5454cefc5c58b34516271d37aab55ff90a30bf4fbd514789811e53399dff74dd1d724063c48ba2eeaa893b12659a293af7362db3bd1493c6807b9e16d4ba2adb2f2c2c12701dac60867684cabd74d991ef166066460f00c5d8f6f71128d2e5f3d952ca720e18165e23f5db706b4c01fe6781d22c5e100a9f2b4be9baa9345b1532e3ef852bbed8388738c6491d21f20b13b583c33bb1c5bdcfac6f5f29c4b6f852ff265da75c6297cbf6d59e926c431fbee45e68981dd1c37c5a74f79ce34fa9e55c58b3d75e19bee250042a02db2fe22b81bf8e2ac3e15c6e9a5a07b0c8ac500f036e7e0968812179696b44fe4706d92afc2ab47766e40c061b0e4d83e426aa95551ebbbbdcfd2835380a4bca67c0733d00d0cfcc04825b0df98a5212d7d1dcb23e51fdc83f683817694872e9803925b1ecfd0e17a36b256418fe944b14c0947ceca629a303011aeff3d3056188bc769e41fcddc17a37dd4bf4b811862750ed2b49cc9b2ce6af06aa6eea5e540dbb57f9fc9e523c1aceac9e95ecc29bb16699b58cc06ca9bec767324895c3aedbcb54815ddb53cfbc8c60dc5990d313d81449add891aed319a867e0699062871a5f88f1c8eb8db8bb21832529878444d3b05dbed2710bf6b01789afa251d0e27815069108b773d4e2e1d57707d0464d941b19a85e66ddf47462b78a82708763af2cd398b7778dbf344ea40c5662fe2a47f934f8a540e6004a17a211f154e65e5be0239c3bec16feb8ed8b86fd01a5540057f4bce1667afdac63188e199cdc02d19318b3ebe3749cb352de93778464204b9bbb58d8b340e5a65342f8ba936087487c9a654d962d3a0620267391c60eb50988557e115910286a692e9721a661cc46e9f370df282d3f4bd2c3b8806cd867d5e423e931f2996757d8eb2988da36704f802c889955290f781ef799eddb8c5697c4f91cb3c096aa6d1615e2928a98ab5ab4ce8772d4bf1b17a99590efeb202190ead17182346dae3db33e641cac77c7692f96aea5f886e256fdd1014acd7598544bf0b0ec33989abdf0d59997fc8a7b500ec78ae84405645bf38b3cbc7a5a5adc318e51baf092527ef21c4b7426c77554de2d7e7ddfd29c0366209578ed768ed71d56d634a1b26bb6c0c4e809522ff332765e1e33c3ae9573efc502d35d6683752ad80e060180d2ef2d0d09c5ba3013a15d9290c892119469bec3841118c34e7efe2ed4e19728b0b273b03742b4debc23f2bc2df8438c8f63991d9aac92135e580a8fcc5055625b9e0fb9ed49a6815bcc2618ffecc28cdddd7e4befeed893364ea29bed652dd26fc0a2d74df2c67fa512f1983f33f352127b60e96500eb615de67e7d064b7a8cfc050efbb000edfea49e7e9d8e7d71fe1175c081e36d24bb1a6eb27880b4fbc87b57da26f9380149112eafb8d827b57cc0a10338c1d58a88defd056ecec461db74983610f7580226d9c7b5e36356808bf10c4ff4c63ca9cdea286374fcdd5045b32838086a54478ea9533cd03d0b78c6f794b7c92ad4719c86098f73eeb5eaa1c52905a9b894b61df63e6bc88a5a63c4240efea67da233c0605d1615637b1d418e8f20b61a21274f71a10b651ac70e1ee372a8e7d1146883df353eda60e00ad91fe9066e227b56707f8c82a8421940d420e6dfe2d2e3cfff7237f83c2f545d9f829298e84559c158f6211798e1ce6d1c0f145815927e9e5da3af3563bcb79b1d6e868e6239bdd6897fd325bc63fcdafb315403942c7765993c153439f177a27ec38e8661d24d3fcfac67e2a5c7a548f821924bfa48a6ce4da4fa1e6b7e4e16b897413667363d7e98c1b68958e8cd91c68f0755d8ef2f6b7eb870eeeba8e3c4257997fd22590cbf8577e4882876ea10e61d7b4d32ba69228469d9f3b4063935384f1812fdfa644d85df78ef0cae029ee5ee431a835cb32844751b677d08f2be5ce2fecba62ed18779580d24f6223fb29c1fdfcd52131a5c202f1a30ae9cfcc83bfd396d8f78de0689aa28be0a477f2e9eead41b798f8df9e04f6f8bb1527f78044323c6209d72602fdee7dcf635710a0558a513d483d221bbb7d6db33eb84a5d4a3270c1e42b9702bdd80926e85ea5ee2a5b42a1e235abc0c6bca36cdbe3f5c5f4cf620dbc6e9dcf0c481a2a1cd6f048bde6e1767d2046ad44b3096f54b14428647488e6abf04e51ef51139af00490a92ee667b3a94efc6b786cbeaa811e59cc1dc3e23d1239493d7bcb5927f5c56b9e9f977b1f894c62c994f854cfc00620d9ab32e14a4de8e3210324b95f3c29b428bfb01c01990953949d87133a9ba70e5e1b271d45f04d915471ed1cb65315631d6266e5faff2152bdb1c375c83bad623a3c850bcfb82f52b3ded375d322ff04b9785ae514128ec520b3b5a3043011ae7987c8349cec34d6b8ba6d2dc8b4734b4c2a874151c08c408a5fe5dbb8a26e35ec7872ce6b929c695362d4661d4a56be4f32b323667d94f80114cac743ceb6ebd173e063a2c4b14bb19fdc080e0d6906c01ac77348cd1ab2409ecaa6d379f4416e5422beaaa11f9b9a99bff950227dd1fdc8dc31d0704584440d8b631abad1bbbf34aaa5b21c9bf65f046c628db968dc93a26bc5213efb12d36a3ce04b0bbbe36fe5e2f06730cb219bf32ae820369e09860efd6702224f0c306e271c1bb3319119a34cf1363b81faa1571e715d47f78b8b25ebe051dd89255eda2827a4b0a4cfa515eb354a6b762fda84ea04b13eda72b57db133f59b1ec17aa98736f94a7d09e2ec57c0b43339c7ea34f2b02ed8cac299a08942011948bdeae2d36e069f7190da6d81556da2e2bc2f9d477c34f5dab2001c2a5621f2aad7abb099bf860bd15ec7e74b12163ed8f9d4977a7e134f187d4b4ea644170c0967bd2ea88ca894bebd5eafe5105b11eae467e3e4e9f93693bdba287d146047d2c2e26d4ff227e8f62be92c17891037edf68bceeec3f0facbc7fb833562db9aaa181a3ba5c1e2545ddd55484d75c99e06d4ae95f5d478130dd083dbf3fd37ccf9fd793144e05cb12d40fd1770dd8298ad38f2838ff7baf92df7b45a05156417454f476ba2d4f712a25929a0caae0b38fa67aaaec8a26abfef5dccbea62a8193b6ca94a12d4e6aff8dd3e00c134f2ac12b44d799c03330de085dc4335f6d52961cb253518c09523825e14d1d73dc0025123a70d5238dd578bf7977b7bb4ed4500d5a3c66b97b7dd4792e966ed690dad82ac9df175d14703e92df93598eab2febec322e1adcf3b71e950c91063b7b9e15fcb5253d3c3dcaf15d7d5979ff486272f6f45d2a9a7f42138284f4075a337026922be60b73c83d62027e1eeb808c1840b24477ed265c89e11358a717e8f0c1507c44b46098f7e87dd144ecf9a8a9c86d865939a7af01a3672d6c7813d89d65550776309dc451b0480364e233c5b5e8c1848450923c686e76b3313cd27b6afc4e11c2227b24fc44ad889ff047a9c76a8894d3a5e8115af4bab5c44a19b76836a154c2fe201c6f2aa908b7980b85c6dbe370ecefe9b37770566dacd62ad6a5e0495a9be7e74df89eb4cfac8856b9411c9ddaaa5c588e8f57212da72cd64a7b5d0e9a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9afe8568189f2ca3a390a8e1019f8cb5c74e596f556728889ed45c79c89934a62544f2719fd3e600253390fa0236fc0386618d5fe3a43ec1ec0c6d8dc22f4c87339419086b2310bcee04173bdf5297684ba24ff98680bb909de7ef5dbd18d3dd141477e7711eb41253913893fcbadd4e85e155dad9b7f06635a7ef698718fee9271db76eba28537a0cba744dd30e92c0d52734139ba08e527b253fb1dd34732fcfd2052fe7f9523595debd25410505f053a69a4b8489a3ff5f265ae1b3bbabde2bc6f164ea9f5c59f6831a63df3c08cc9b730943246641aae3cc101d14f69c342dbd4b33c11f001e71c01bfd32e3d9c5ee359eca13cd505375f05efdcd97ea0a3468b521f9ab3c488e6036b3122c926648859f6e065f1d7be0e768166e04b630235d22e5dcaf566cdd21b47dbbd308965ded0f61e9469405e20ea815a5928bbdd176c1608fb9ac05970e2e2f9c1b3cd26c592e7847d158aa8a4f64b5371f9bdc3c1c3b6a8e4a25a555f27ec6b401e6399111c06165705410cfee27f8e4b365ac80e97a947f1cf569d8678955a9cc7502cb4fc030eb45068d8b366eb8e9d45ea17788aa8073bfa448443da13b66884af0d148f94383901b680c3d4477650fcac5d052a6273bbdc87e30764be14b2b3dc351c09d5d7b9a8e34808b18d31bc9c0a5bdbeed4a0c4099c02207bf9fec031a64e7356a1956a555ea4da57a35590cb529ca1b7304097200101adc3c7caf2d0bb8fc023fa10f9f214396fb7579a515e696e328d093fc7029811473beca766e112683e964ca6194463b47d19996619997dfc48ed27c2db276a22cf56e09b55060eab69a27e42ea536fae457a3ace5ed88f2e19eb2b87f289f6a75cd39e0835d2f392e9bf5b653d4f9ef89afeab2693ec76086b186ccd1b0ee0bff8d4128f3dfe3bfb21b5a7bde875b37d7fc5627fe75f3b12740d06c665f520549fafd9269fad217dad216526ab54763bdcfb11e0abf21345296bab387d88258584373ac1a64428b91f7e760a785fe3d0daa36d391aaee16fb331f932679c24ee0be7af7a76e63c7ab76a657ed619f01c1752aa5ffe6d7d2ea68bb91e7234719bf5350600c906b6ff296b8b1beb6134db3fdf3596983348fb203e66b7b5a761bce68c7528098c36dee9cf8d9d63194ed0abe23674945dd7fdf98d18c04d67405a8563081815c4b4d0817a362eee676c5d9146584e701ea152c5a52bca4bce65d07be3892871b97a6af074fbff3f63f84ab0fbac6b4ef590b5460cea40ecd349d26f2fe1cec51ab74ea5a482025c0d04a53bc8dfff1982146dc733acbd57357f099725d3b33dfe526eab8e075d887b5a7a4dc9941eea27a129c8f6272e99bc5e6cc0dd8fd4e6948dc924ccc5a5a4e6c2a52e3f21f61ccc036d9575c8fb7c62fc0ae8932d738ffb050bff0f971af770ad15fb82729eb313dcdce53e547b20db79a7f8b2ccdee24fbf8195bc68ce67c5a5352e471e4f30b9bdc7052dc456b985b7ff445ec0a97bd763c0107df362a42446aa3c4519e334b14f70df3ab19448e546ea8c9ceef08c42f19ec25d29b9957983e890f240f9ab9dac3df8031af6be2c881f555a402c9f11d7bc0c68df194c44f011b85d79c16ab71556eb6f51ee60a8e0ae8e6eb4c98c222951082d3844c517d918814632674cb37593dd644434d18761c938314d0280ecd595925e00242ad1b6477389d1dd28734cc438e3b095f68b67b6af76ca92ee769071e60e3c838c0aac762dfa73e04a7462628e1579bd756c841f23f388e124b78c2567edd1d70eb6719a4d38039acd5f96b00bda0fa1b417eb2a225bc4142a02dcd96942c93e920fd67aa9f8050d98c5ec72c0cbfc7d28f457659d75b54f76bf9402454e52b692353a8a19fb39541806b2ea1664d48d1f17b296a41f1ea594f046ce9009f641f9e8f7cfbc5ed1af748ac51efafaf721f7bf58f834f3523dfbaad3f04cf5d72ba554abfa0b430e8b6a95baf0574b15bf3efd20fc6593fe4f0dbce1cff19b7cf0bc850a79e2b154974ec1f5f08fbf52083d38bbc3c0c5f0ceb542e2377a7e2c59337073236517bcd7163a4e3cc10a7b5e796c17cd221bbbdc21aab918ff094bdefe770f0ad7bb7d71089bcdeedee0b2f2dbc90d844d718e40343881d5bc49a59dbac71a6ad65c5557af04589d0f76828f24a0f8165e3010e300a1f7f13694de04b5b00c141f6629b0a611db5c3255eec912e4551dc88e6decb0f8888535783757895d249e8778c050c784f6e1aad2854b0733a3b6170e945e1b47a04415bc4f08e8ce995b3dd3fffd64dd21bda758bc2f94e46b37dff2cdb0d43a97bb1e0208932284ae69adbc29ad8644a6163b7ea0974767f5e0d1a144f898edd47f5bfefa989f3b96fc93b294ccc5165e5d633689723a8e11c66870e87172c69b36343256011de5e2612e44ed9b07c9069c61759d65b6084e08b8e9fdcbeeed621cb392df8cce7b168519ace154626419b9df49f053638af0e98c6c3f53b5e3217f2961e0d855cf36f18c4cdfeb56d38793b088f6cc60443d32dc758f9db1289d26254c11b83938fd331924c5ba0906f3fd16ec5c66e79a4188776dd58a67c7d2cc27b107960bf7bd5c79f7f48e543e84eb8cf7ae55d95e9ce37ec413d3091c9464b3340c7d0b09bb5fe66c0af185c294087967dd78cdc6efbea92f2cbc45ea035731f2904113ed638d98eb011f1a3fae46dc549c14c95c3b21cebf2867129b8c6c8e9b5298c4bb987cd6bb43800e2b1c65f066175dec07eaf75967c02311cc912a235178ee8e361e19981aa4beb5910ddf42a237c1bba2ea14818a65d428e32fa37a89b73b6f02f58ee53cb36a714715385c483990ebb23ea8781a622e38fdd767135d9e61aad0055e22058de7379e45f4e1fe95738f0d777aac351a23c384780c9cdb932075e20d9c3852b92563e6e122256e3eb29d6fa0449fb2b4e7d5cdfecf747524d49505f7b1cfed4d5eebc3a811d907f545cd7458be896ccfb99aa6e81fe3a70d40dafa7dce69ecb5b44579e6369b4f29b3ea344ebfd3f1bc1cfae5e76d46bc58eafada05f7ed21bc58e22b7c20fd8356e118b7a21ae9cf95d14c32608837d581dcbc979e916964553af773070a9d818aefb559f5c051358db5956f144074db138b4bcbaf455ecff45b785ff82e222192ce3f66fe99e284705974bf3da45502498336dd4f899799b2e9430c1a4aa4cce72b6611e309bf7474b2d9cefc3644f7a69e16d27db2d6c0a8fae3a3041fde2801fcd90acad8bb51600165ce22ab0035853d1c08ccbffbf6d4c3f871a8bac8dad89ebf1c6de2bfca1c4fd4590a6d321cfc2a24f2a223474031070da6613d6d3802140fe624d9f069577c547287f18aab9748ebec15dd88a94ce1ba25e2d91e55d0ab75cc359aa6e7f079d75ae9ea5335e72252424835cbcfdd0b1f40c92620ef7cb1c874f9e12856cda2f71d7595fb2ad768b9d0d632ca44a4887543760b496ad7d236ae3a7ffc15a67500d010a54a7b010ecfa6bf4d33a083579ac4a845d8895875b7e1f20de00de8599845559afad2af486e910e8b730b583945112e53cfff1f3c99f55950bdc638616c8455bbd9a50942b41524de703e4a5f197e9205773e927b1f560e9f3a82b5d50894e8a6b26728f392468f1efee793456a8e6a3ed537d769256c563fd30da9046b5b679d133ae6edb5f3ef6fcf4842e675a3ce7d08d64f6cab153e1a02c97256a3d1607daadefefa66dea4a237bdb2c17b6c7fd3332bea7a9964c26815f40f875ea50677cc8f2c3d1c0c5bab61883ddf69da95c83da35bcad42d3137a3fc483f2600a6fb5632b3229afec45c1bf09c0017205ea0e3b01bcca07b369fcd83736af71302d8405c627f7aa3f6aeefc318ba688a98da8550319da5c6bcb6ddc1d79565e184d0def15dc8caddb53e8db00b5b378fd9c91ba6165f607d6759a735afe6356db3bb69b9c5b0f3ed2a1a953caceeff5177a2f4ce7a59c27e2be9b71b7e7af4c2e90c4e8614164b6bfdb39e8535d9fc56d19304ac3ea53ee2c4823239f328662b6efc233f23f480d48d20d86b8e226dfeeb3b9da12d4badb5e637ec1763df155cb5ae178d27d4e46c85065e63b937aaa015a36a9de8b08fa4285452f200bd8cce21fdf93f0cd5be3ccb16417f3ee9d672fc08a8ad4c892b03a7192bb3f6a324e97cf4ce0d0aed9166097048f85ec34ff2fc4346cf22a88a5b4c08a8e7060252b707a76f45f249c2ae3c81d34266eaf5a87958bf09465494659ec96bbd35c955c615cf1244eaf17589a5a67dc9ddda9a49b241c1fe5e47e4586c3f15e291efabfcc385087eaff7c87e6c42fcbe178bd1497d5e95ba448402b96e2422262749efe9bd0e8e7c024396f6554f6be760cc30f45f4618008f1b6ac301735532c114bc49a29f45eb79b85127fc376d42d14948fd419563fea352b736877808eb26c16c406901a21537cc6f6f6b83e0987b076cbcacedde0de0f0daec46bdabe3bcc62d5308a922710f810803da7899d056383ef03849e3ec11e67a5cc7c4b28a6fe05773a645e02c1862bf72add89870950e8463f6be6f7167ec3cfea8878e8114935571eb1a124bcb274e8d74cd4dfe9f29e3670526468b127444098cc721d5006e84ffe587703c6253f3950fc04035800465e2ca243ea4300358549d2c7e0ab3c030f95c021a8cb1ddf7ac3acf63648afb21f80f53fbcd9e3d6e345b3d721be1a67c30a9bfce6b6222ae929b9a86ad73889d5e133c9c85054e9752d562db3b8a0aca891131c7f5130184272ad509f8044d729350c3c4772d05410b72ac9ae2a472d2c4911e219295a3dfcd053c92dd00167f9a8a4c78e7ef4e05610ae615c4fb890c11128d232a93ffffd98d71ac4644937afbe0cca0c010777bc76216d8c4011559c634890ad012ef69180f38b454b17e59855047b23e03ff79acaf1bd5ec6ecef369a4edd48682a2b7b9a7e75fea2168dbd7fc2cc8201b522efe1cf88583fb18aa583f2624b29f0b3995571e2442e708c6f4a814b20757dda4fe1174ec637d36a72ebf646dc38af6eac99ebfadd1c4bb5e701013a5d79befd9b4a959d9275638fa42273aff0117b01b727ef0769be16b4965303691f84f0618e6da3b091001420ba43acec409942e60f787d74ff0877e312ae2c46c14231269f12516c3f95b0ed91da1672d56c435a5045230baeffdc0f6e7e53be4b9b8c410c717d39f4979c3e3063d42094945a08a42ce06cc5c55770a85ba96d5fbd2077239b0f80e1423d9c0cd34f48db682745d33261f13799dd784727ff2f6e11dbb7f103172e3539dc4a570016fa0bfde7f9ebda67ef929a2dae862668768fdff0ea0fd6a4117d8feb41482e6410a0ff54069a6ddb6d67a13c7264eab20acbbace0e2e2f6c0ecd9de852edd29331629c51c2854b6da9673f4991e7dbca9659aa36e6b4869ec9d7a7eb907c2f07c679f0f8f45c5d038e28117255da4c0c2140e294424474f01d2db0c033a0097554040988f6b658271e246ad8bf9abb90beac5a77bc6c689a90d20f355aabcf6cd851e46b6f868430518f9ddd5b17ad859841a787666f6575a12905afcb33b1de96d363e1a3948bb39f46ba4a9a2526b759beda60132fff56a09e205044d14ebde72a27bfe8ac5da4741cc455df2234f590109784a3bb98cb118cf2071b979dea1fb5d6e7e873447aec23748713aaf658f76d27c9892ddc3da7e7f653baa09ab6a3b2a461dce71f8e34c92155186cd8c2c172788841a720847d7fa2be153948d06915edc5f21243d8e61582eeb084d42e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8b940c7751bca13d9ebdc3d9f58502d75c20d4c3a1826f2fcf23684c2104675ef6d9b4c41c8a78f148a385f7496153b62f7d6f62fdd343b033bbe89cc28f65962b8bfd465ec1859f3835f3263c50f999847ba877882fe1a66a49af99d35cdf1ceadd59752645dc1b0780a67db84e20d0552557504a0b3b74cdaedcbcdfaa26869321b639b61333ed5e784fbae4c62e757997ad6e684d20bc55fa9e12abd4d1778dd5b02700e7bc70bd4bfc700d08e4afa5809e9af88e5b388b7557753d9c3c72939fdf62aecd7738f0fb964459c8993ae2661d6626e0a332e982465b094c71944bd38c51decc6ea49c382ec2630ca7d134315fd668f6e1f358c6582b62b73011ecb966a543c3e987844ec2314acd14fc90e1cde13b42bd1d57025e18760ddba2f10cea63d36cc6f37eb26c81e47c50fcee88e61c0552f576f303d0bcde3330893fc98e9431c83b9762414b4ba4d0be6245ff3bdef9c7403445d7d891493164acc78e0333dcfd2f379dcd23bac4989e4bcdc8fcd092884a461ce9e6ee7eb55804d58bd0a736950020dcf1f9cf2f2ab3902f97103226d95813b43caf436e77ffe05a0f8887760453154209685bbf74ae40053d410b04b2915561a6149117d92366b09ca6ae8685c40b7186cc48f72fe9528b3f56dfec81f07b14a0d0a1bdc8722630e0d717104826fd7472bdf5e134d6674fdf59ba0f8195e3ad30e8de1738353c806fdf65227062b7f650c8be93b5e6985bc32ef602da91ca6cde50120c9cd2e2c4f2b5eb0c6ff4cb9469ef552ccdb059357ce52b48db7b002dcfcc1ab6d7c76db322a8bdab82decaf1a8648c817f83b005897ac0c9fb754fd1a3dbbcec8c77f492cc3bfef40a83b9b0b295b4056b6085cb8cc2918c6a424048a7bb20816f9c54a3f7556e2f905281ac92b1d10007410dd0c703ec0614dd75d28f9966b33498e9bccf40749692cb75f645cd933e96c51be8cf43574d0d1ef62f330d60f8eec1f99c1d8e1594b2a62f93bb75681dfb35717d0630c1009431eb611d8468d16b1f59f15db470cd8fee702fecb6bee1ee77636f2362731453d1293e472335281dbf4d4394874a4de57130bb9d5f25b3134702b1353e93c2b40ce313b3b0f4b912a0b9aa527ec7f9199bd51001792c777e463899d8ac44c6f9e798687079d8ac0bf319f25bab3184a88c72d4e01484342ed7309d55c5c0eb3c8417567de2225369d540124357b5927f5b62082d31aac3963734d756ec83ad5227b40b0eaa959c96b7d5cd077ee951ca0c56c02e486a006a0a3f810c39f16260006e21f83e3369f79f59a403afc3760c3429a23fb4c8f78ad76afec245cea194c40aad9105cf1eac7014b977729d97036b3a1fdeb97c6d6b64dfa41ba937be94d52deab991deb5a593c2ae64f590d9bcd10565f4bced09d0aeb7302993fa2cd66c24b833fdadff8f5e9b16d92a8ca8ceeb7b369fdc1e17ebada8c4e5cb40ecdf9afc70740891a356dc6e6c07384f7251a53a6d01bd85e9ec0753d2b67a33ca3e7220be09d6a61fec240a16d52a9171aeac151197fef3116d2e7059a2b12bba659eee4e5535a5920da21b5b1e3ca60bb61b024fdc2d269be1bf55814f6cdb352fceb3adbca0afe858740c876c6f3fd47fc2cd6f1dc76ed64cc9973b93dc605ffea81efee50d10be533a8dfa70495287b84de49e3bf2f6e7162078d663b2da05d028f8bb2b5163384da1b8008f4b28deb240fbc45995e06cf19c150f2ecbbbf2a0045c0a2c3954598e5cd39742a485716f1af6c721626c5de9ac94b17404a0f80baca5aca097183b50476cf3f9cbe2f2ade5a87feefe9d0ae1f41d79c380f0d16ef0780ee1af12c133c8c327845e214078adfcc5e25efbd2bb18eabc1a86c1a991b64e5619be6c9a537250d78ae8353c291b7eeace993f1a073a3f15ecf2504c727a99063018e5e5af998c6fb47c45edc131081b0064186ba56efae89bc7830a9529c63ba8d2e52af33b386a35c10650ab709702f376e71f08d33c97e7229f66921d5adb46124e3569432679e345d11ae722931f291ceada989801de49feb604edaaa97f119f8e14598df891a273617c2419aa9f69224d2082404c1702f8a4853f67823dd3ac3f0ed95884fb240b5ffb94ae3cf9199610d048751cea5003c2ca743308ba3eca5882ff3a057fff478ebcb80cd8e997a5ea3a60c5bb04c5e7068a3d02653e8b267a343d3b5aed2f5e819ef551392a2ee4b2c00c13363ebb2b9aeffaafedc37d53f05be82e7e6e708c3d58d0a380cdd1475f19a5fe7c6594e8c182eaa4675d5410d4fc7fe6a89440c03aedcb28a20698ebd90d50d0d8f04c1f00d47e06bdce73d4184306453fe372b1ef0740d20445273006316a8520dc43ed5c361843e0ab6c5b25a905893894e4247ca83561e14d3039a0527fdf69c7e89172ddbf30c22f2b6273fbcec599329ba567c05c71839a0852aed3fe422eed26f25a2103f939189359a31a3c8d831394ea091bbc10fb4b4b974e2b4afab95a9634b92c65f9c3f890d41261e95e8dd56dd5a35d82704ff1878efa6ffdd1718e2758e4efdf6d4545f13aa53a0dc3ff593e01daf0c366d37909d777e99a33859b32ebcfbdfd33687b03ecd18f23b78b53f8708199a5fa1ba828a5900b42313872f06a97873a7fc01ca2e422cb5917b3ddf7aacd5fa5b0172be75bdb3bee5ccd07273ccd64614e43a00bfa362b06c4b60488e809219474ae298620ec2c79b56450a1afd82b4bcdb2942a230c00e8fdffd2dc0871885f88bf969b37478031a5fb359d4f66f6f2aec66452b7e844ce96ca46ed611fab23d346ba3d87c6d08d01d90e397bb0d375ce00f4976fc39ca3facb8d4d7f279a16992c60ead9b18f525e8315230f3301be4e531878b2b33b2ec00194e6c88a5534bdd3b85e76d32d367f2de8156c2089c3c473c61c082b69e5f06ba64a1ee8eb8a14ee6cc344feb13016c10cd9603a364b31b3c2aa941eeb79a29776bf268c0b311ada664349d68d993b5d670ce4483a0d6ad54ba1ece4d01110b6a87126eb1e0804c751aacc71649cf90e178d8b3c1618012a6ed5ba711719c552253d98164ed4fe5cbcb12e784059c3a6e306c90894a6548025a8abcbb7c786be8305bac62ffc504a390d39960c295941bd85075b67619b8af6c31d4242a6b673e87eb2830b1c95ea018a91de2e3f9d6d4361f0b21d50f072b076804381cb99053aa110b078803b11babf376da6c0eb4eadb058a69d57e0198e21ff631ac31b39ed4c766bb8474ad188d510b378c2d9b42fd8e34fa843e8e29fa169044026ecb45263f1f396b2f66ef1de696ae11f670ec09f8ce177eae2ab08dc465940b4eef08ac1774cf6c27df73cc86c083440deaeba1957834a00a1f53b8b507f3e18ceff46b0f8f6820aa3c3fd6d286381b08fdd4eb66f5f5ff0d37cb39ef2aef5637d5d38a170f887ad616a45abd9df8c71a89c8c689ac51ce50a28a88328627d8dbf54168fec7b83e1a552051c402b86646b23d88eadcb76376ed9f6a47713125a7ef8efa2e1ba08cf7bb2a83442fbedd3be384ae87a30ce60fd459facfac940882d57ce1811dc83b9041c25b375f571175b520d8f20f9ad5df6c6567a1b704911a306e4fa07832f73448990fd85d6162dcb1c3365f482b26a69d9a0da6f0107df1e748f31aeaa10466e9b3a0ab5d41543c1817b4bb8d84f9d364b75fbcdd434813875c17e8bedfdb1a733498fbe61fe71636ebcf31eed9d6480ddfd9b257a6c593d639e5191bb5977384753da606423a4c8ec1adf4a5b15a15c4576858d26fe5c55d81f045b426747c7d8260723f0a8758fd37c2375dea21c332f28d1e10b889b47a4a79c19d97b3fba26cea1eb9ecd86ca60eeb818e9c41f8a164956086c734554cff7e57a0c02b6faaab326a784a9b670fee34450c4e8b5c41ba407b5210a0ae72abed3ccf2e2a3cff988f444a9523a61a4d0a480e9855adf929f6713be4f4db75ecfcebe4bef6c4685dfb6046d73a52e59c47fdf3f2f5e3fd716140f8c14c12d4cca454168f6d77b69a2bcd794ec2b2d3e3fafc49a4f6a317488ea47b72cd44d74e22d9f00d07ef13e1225be7ad125aa78452efc813905b88f9782ab0fa5590d57593c687b7e87a5479acfe24e6a6fd009438d422d4a42ab8875806c4b8f769fa09f12034781d5fbac813b4b2fcc108af92c3a42fbc717ffa6911fb0cd1db36114e7fdcdea3576f3db613fbe975aa4a8ba219778e7339de938880e86d05719a1d5a07158957b524e6f717a5818ce6ea56f51e3d0d2283f3c8384fbd5f49af402dc7438906787b4bb571f8851a286747aa9cebf97c2e33e1248bac73baecb893351d61e6d9a1903f2843718ac8ed43787bff11cfa88859656fe26dfc1b5fe29239e16da007fad61d242f9045f427d9b02f6b563971dc2063dedb33788de66fca7cc442a5e3cb5e1c2c7b5df4fcc03e88b6bc04978664e65649ae45f77bfff80d50477c3e93afe7d05aef4377faea15e4b16f5bb19c77ceb610a61b366be7a055c1dd509901fda7947287f939debd2e208c5dfad7ea2307768e3841cb86d4a73edd9ecf3c73c5014095996f08f9793bebde4f0088c1ec92bbcaa8846e8897f8f105ad3bdc5e54ac9aee981454f32a1240b95791aefd1a59e451d0af1db1f43df0ebdbf9fddc2a19cdc6524235426f0a7e58a7d228307f468293b225680e8c7cee20c14f606ab58f095a59e3394f4a1d981d6e300a8a8126feec9314286dd782d1216a416f346a10f51345d0ccc9e5efb09fc5307d4f14f76173cb83be2cb64e33574da36391ff1a351dd6a1aa17e0459628ab78db336e4ab29e4c9df584614d058e676329ecd1dd557d50cde2b842c3b6ef5462e72397632c2ac9fa976a0c7b5a4aefc461f329729e5c077ae4ce6dc164e3fe5aecf1b0b95f26bb88a9ba2c68f925c2b9eb728b532e0c96700972ea28c88add3b712999bc271b623c2ee9b65517b55abf2678c0f60776a8a004dba6702ae390328d042e7d406aec556c473d43222ec16c0bafda5bb1a8265ca8dc9eb634b97c9ffba7a694ab1872eefa6cb59199ae97ec8aca0ee1af0915f08afd9ff226a88a140104535fc44df03581df09d69d825409dc49d0438895520f131ae7666388f2f689ccdf899410877e189d68894d7ac597726329465995ee0b91b7edd9ed44bd2f73e8b1b5a1e9c2845af2df9b10478b2635387beaa470bb136bc4c8f09f546d0f75970619eec988642d4d8a42cbfea9996884fba1e6cd4b8007d4adc192c8267f391e9d966ddec2760649dcb8088184070116abb3a88dedf66298da537109fdd85a90ff283a580408e69fb0f8f81a86f8fe3e56fb812e2e771f2c783e20066b1d2b0bdbc815a1e59d0b1d377900d730c5493b66804f3b00541c9aeb517c96c5fd88c1b220b519eb45cbc75120d407b6dbbe9d33a916ee325e3c8b803e1a7537c0ee9b841583067e091ebefb73856715e27357fc1cbeb5aab258339e6cdd1eb8f4834643d9656e8e1a95ffc7f83cfeddbe32ef0c72e120b37b6485b1b2daa7dca13e0aee7f66dd572fecb7dd70bbf90c2bde9f61a333fef8425bd9b8ae557d90dd4f6ba58dc7cbf94f44186e25302fa5e5c4adb72a593ec85211e38843ba3a6aff96751556b3cdcee32a9988ebbb4612f181b02a11340fb963bd8004a6350ac3e0e3088f30126ed51673bc6f9dde81497cadbb3b15cf0f960f0086cd2d4b8b53637ade9df147e32b90d1aa3d1b21a0d0b68d3116ffbc8a5c0498b9ee5d8dfc2ee8305b040cdecfd7afaccdb1e9a4b7c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb8b8663531abcbd5d3e3a9f7ce494d479351a2660b10d08f8ecbc8a5a98f6f3b2f062393b053cdd618a29d5511490ba69c456843585a67bd803d3d355e94a9cc1fcaae5cf5cfc328c174134af381d0a30e363bcdcb450077a9089dc4c8ebc9a048e1d61fc50590fca8b681c483ae44a689835c146f89daf630ea5dfbb4a74705b393ecec290a62c77bff849f261f48deb2a9a24e80fce1a7dfb44a00c56d562397df2bb238c4b3e1687b00b68096b037b4fca98826c2d812c4d792a6dcc9902dfe722c984caaac1f240e4a622127f7330d951356d6a4bdcd7fe5b69dc4ad14e2fe2f33ed31c940d159a0849efce1aecc77005040a2f287ed945c45e2ee109ad7286d7b3ea8daf40b5f9714ac4d90555a1e3785d4feac45a2bbc731a92a7d6726c6b34275e090c04f855178175658229bbb9378f145671ce7ba860f2e1e483a0f7e54df8c38f145dfe6456819a80ff93b5e7ed1c3d10769a79a2b73a7359d5fa2e3117c782093f223f252f5ccd1e6d102371d978f492e4e7acbbd9f731331d60eaf68df43bc8bebda3b621b831a5e7faca3213f91ea8099d2fb43984f7bb4bff56f19712d58ada3a35ced3069eef8cd16d43fd5cbe6ec935842532014aed4a996b3ecb478f23acb0d51e364f512e9c28207c94dea460e3f890bd02dc18e8bfeff269fb4a0d202ed72b28ade78661cc8f0ebd2c87f1790a81e136820a495d9ec43051e9c8a08ad168e2446b6c23a982f05c8ff4d59df1a749db9a25b66a46f2b0a4d839a54418a73a6c2a48023f856a2dfbb398dc11e99850aa5aa3b5f05e095b059d8bba66932470259d3d1ee86f8236edc333433d6f18de8c137dadb7c8efb5ccaa719d2597bbfddab75d4dfe15e1d619b0f576c5d8f616cc99f3cab38f1be95f282736086c31d0cd7d0f73156c60d4279576837b356088e90d98ccc67f6671959cacd74bb20e5049d04c3663a2799d1238c79df27f57b5b54450aef8f5119a2017bc38fff5ccb97f555d8c0b6e34b8f5e888aaadf634c6daf11eff712d60916204bf9b99d7755a8dd48ddfe7c33a328ce238cc99aae14553d3becce4724e787d88041c8a72d72083ea5c59e72eafdca12a5de86ca58d4d06c7fb148b67a7e2498078460b91a9005d8d5765f922a00ec2e9eb61cbf8507d696c51dc520f232b40d57022db910d8c3872d66e7b5635b9589d03dedaf7d260616cd9a5925069e75db86231b2165b32762a38db6b26a28782c10855a2a3f42ccc625278b9ffeacceee7610e6194932be42f44131e5685c9c2a8ec8275f73de19e8ed97e0cc496a4020614fc5a1f8271441bb60e8d3b60d07b3880e2589889152992729cfcbfb2ba36f92068dd09bcfefcb43895c403c39093d73863737205453824787accb81a5a4d1d6c06bd3507587f9be5875818b3279c8cb233de6e883afccccd593fee73581db9a88d2ff641be1047b61584819af908026f6d04eab5e011825e070dcd093f2901c60a072e91ae674bcd9e351e4e64741f483fb89a2c81127bf4daea734645a53b0432eae41cfab7d334d2aac892d2fa5896c0b258974265f83edfe22c56b3de3f033e00da0887afaf0d51aa0f87b13b27f244f7fadf1cc2c30f5d0ebc1bb3c5d1ee5bc3b37ffc88444d43ab9c0a44221ae19a5543775daf50194915376b723996901aafa4a8cdd73fed812bec373edfad5ff5f1b91509f62aa82ca00ca37d900db6686531f293f571332c1f5f7bf88378a497090ea4816e9e0d367133fb48f97ac128492bd34a163b8e1676d99ae8947b01fd60812e06bb5251dac36c8489c43d22a9253a271e9dd0e59212bd5b2260aae51707a4a55b5f1bf2430b1555b9187a9aef259d387c2678a91862714501ecbbe52005399380b8eb7272d0b4bab20e2ac7143043d3a7cc20fd3c1e4fcbd767f7c7a98ec20f1d401e990f47c9df1bf4c0450ed1db161a9cfdcb94f0fa19f7e8b68a640270bbf273679a2392f52afdefbba9930143a1444a14b3a4fe572c9e7ded365658f5abb124c908e487f4c7b2e95991537201439c0356a51116f6142507e0dd0a75ec74bd89c1530d2358c04edcf33cb38e79a4d69e2da296ed500d54927fe6a35e8d9db5515e67137ea08f8bdc9c0e4dce44ff6c6aa9323865d3e868c88cabac45a75f5d299596d04c7f6ad2222df7fc553740f93391af60f2ab3213a680166c5b17a38ef8faf498997ac6e15211be90492f7354b30b73b4cd5a728a5aabfa346badfda7832f8b30b39bd8bdc53c2107686697bb3686b18a8c4e08eadb3f83ba7c83da44da9e882444c51e65f528cfffe87d40baceab11cf257a1a2d0e06d0fe5be9d283163776c00b9479886c97282ed12c5404183cedbc221fe53a86d427a6ef301406a00a8b26f368fc9ef7cbc05f2ada6d00c2555395469d4ee65faf3490e3ea43c313972ba4e6cbb9c15a417a8a260f89be59c9e34fcb9a70de7dc5d7261a8d4c8611448ba2eeb67b6fbdb60fbbcbf29e8119a3d49bf5abc5de2b0ecfb7124b68fa2075e4dba47af9b34fe7b522701e9d7887f8c23d7d2c28ef8ab50f5ec18d30965545044d3838015ae5e73b64b85da8dc9c1b5259f3b5642a647316296d4f77409b72a5b4122e665c8d93a169e3eae7486e3e3a989c2f666278f9c10367ca2bcde4bf69421a1fa464b31b364fd7e48be05e202907ef4f33451624df0d4f36ebf890ddeb8f24d4500d45213de4a51529c5f894f24fd41c2fa00348f77f2cf2da952d7c02e1c93c52df57f4a8ba56821539f5f0f67d8d6880374d321a131fc1dff251bde7b045c95bb9ff69a03e46b1ac30751cc7002c1f6084e520cb95af3f28b44a2626a978286bb39e722aa911446e4eb947d5a33676b38522c60e67b4742470d974f52c10893dfefdbe4c90496faabbb9ebeb7908610c3410678c62075cf21aff383b1961980baadd49cb3a1cdff7c1cf6e3d55ce0ab7b844888273291df72c243358ccc8a7b4d9b51048b64a4a8579d33890f581bb528449d1ed963b8ecfddb42ac547cab0c650e3257a29ed277a10e518682651765f302a10f88cda6f05181387553d59e0bcab61d601eace78f6ba4ae1a6ba1255d1b6bc9f0eaff262bc71e93c161a9974b56c27d7e54c7388213386b857bd89225b00f1864c7ebbac767a4c70cea005a4c53d5296f5da7cac00b0c7d649f48a97e8e356537b838d49b92f9245cb83317b90cde6fdaab03814edc9349a5d96ce80c3deafe70c9cf49c6668f7d212d471fb90c2f1d4808d892a137d12d0ef856c7bb880fb94ecfed2e9ab27701b8975b381639ca127762664b609e5d61647d303ad80612c25c294272ec10de6a594b79b32f9fec588da37f62f213bce48cc8c2acbd35af1cbc24779e39010f0c171cd5fec8d6a7754f365f03944c332f20497ffb054a7da2e9de9a1c8806e0e15943bef65de8af395f31d0430460764a734425114540af9a18b6a4679fb052f28a2bc30dc191905fe11f3e17b553c6c27183ae48d91f03d7857517313c5c4f4a82cf313d580dec7280add662cd1834d247980cc2256fc88e52f92a37df3c8c0f52b2682bdbf214cc805739eea8a2b11fce7596d2b61332a81152122ebbb5c9848d287b79f1b7ad254cd7b214631b92ea92d658025b5e9efc9869454615ad2f1befbdfb883ad5654cafc0ce40b0cbd41609695870e0bca07752c394a353d9b448b66c78023e61b368613e21ff73dbcbfe4151d0d88040e5e0acea464b0ad4212a349e77f07a5c7adfa15a5778e4cd0914221dbd8936f39fea1635561b242199b3ea5c9af62e9e99472bbdf3585da84ef9bb37b5c7e98e974ea56dd8604f4dec94d631f845c307f5ca1d2a72ff19f477a63dbc4d347cbe158e923271a5d7fa95c8e0e249f31e3a7b318883165ec9299ddfc983adb2872ffcd642f7e3cb5a98ebbe672d319ed4f83c879d30f631982a16a54d9a89349c345aaaf195320db4c883edea964a5e0a7a5af122d32b9edd9f6df98b8a3f81bad4d7a04d9793545d5fc385905cef464443241fbf561439958899933a76e199bdfaa3720e032d91e3ac42edfc81ada970f8c8ba6ac04e36efaa50d4f297f408e3b99076782fcb9d98e0b590000ef8a52a7f2a5c163d59b7d162995d44b812371dceb863d83672074e65b49a46055371cd8c75c46ab7000ec0c5807fe16306b289e923d1220d056b651aab158da8ba548c47808cccf1e36988291c51ae39cb39d4a277fc040bc8b46714e3d779ab8e4baeba8680a8dc4311ced95d715c4ddadb4f79f685dfae70964184153a50e8a135d9140e168cdf70b486f475ad5ba46c9e2c101b3d28a37b47ad050d66d660869fcf86d3c7fcccf7e0fc0ccdd1b1204367279bc951fd521d01a1ea7ced645bf07a4fd3e3f8c2addabe6fbf93d13a8886b620e4fabc2cd4f16567d3cf4e7101ceb8a3d716371874b577b6a2970332f4eea08ecb1be913297694615f0083b5d175d666119fe4097f5b160daf401ab55de58e89c1bc55fdbaad0b9edac89a449719b4b5f6b6d74209f16bd5cd48f18f2971e3f748686483d071f1f18a29d3857908eee5c60d39be0f794781f11534b286cd258a884e6290b429732e41386ef999539b06c5bf278566088da157d33ea37bd1b782f2a7d694b4803107ffb78a47bd751a8538d12253ea7636677befe6460a6af53ac84e7905dde0f6c561ef3bcdec462865dee6ddcc4282fedb0dc7edc7d993f9464134c7e78983ab082b2149a081731d55eaa9ac66c37199aa10486b41e35c725d7786cf45e1b76bd969163051e39facbbba48ab532d7c8dd6c7cf9ad4cf360d7726c90d85a2d7d76e5792f94b64017cc7c1ffd8e6fe597faace0fab0b3692c96d7c24d365f319550fb48754ca4ef8f1fdbb8a1ff4ecde793b37a97a58f8b0137990e3b74845471614a250853ce4ba3abd0749c91b706e35c98f635872bc336442960479bfc74bb886d8f6a846a1bcaeb4c32522f9bf7fadb4e6c03fd9390290e8a193b62825218b63978598c0b518db7f402e5111120ef1ffbcb09a4a139aa5aa6f930d0c73a742e8c82822d2b9788c9feed690d855f2dd5e45f817c08f75dd8bfb804a18342e4cdac47fbbd3d4264ea1b5128b341fae2668eb7f0b84f19f0aa4500d189cff93cf288b7876db2ec2ab523029cc24657f65729a20bd92616d194cbcc7eab3270ebecb50d6eb74b6e95849e73c2c4fde2cdfb8284d57a1cdd1ca5067d89f25ef752f14f2789785ff505c501e26770f42fac0acdb734e46dec6f892f39a2bb92d210e06729924b166b7c03460769515c4456226c873682b69c59359e84b97fcaa5b66267e4cdb3cb55ccf2039fde3d3c1f03069bff683b432ea9d834ee521f63203fcacf62485df169e52e1da97be6ecf1355ec058ac87d2eaeabab2b2a270c6e609b3107264eec23fc78d347b1d70703cd0917f1ed5bf895241b3c2da059484b008164b2c5e0986a9d0ad40b3e3d91bcc9b11392c84b0e35e267cebfd70a9ef86ab6cb8e8f533221f28c3fc7e3266e7be1f238c005a8be6f334917a1ebea061e6d1d8b2ea37ca7ef12416210b2ea1719b6b0f5c572e5f2cab2cf552bc0e0255b63651873e8f708458e6b29a622493d8d7328c9de930b70c7fc311421e8d8142a49507f9ebdca5dbb0640bb440eb5ec2f1029c19822b26153ce17d3377b185d7706af4a3d1813ee91a5bf58c0ce10857af94a1649fc042368f52fd2152c89a0e986cedc82a4f230668694846d5d90a48629c8b21d6ff99767dfcffa954bb591fc84b05d60735ada6eea9b4cd25d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h74961ebbb67914bf7ac5daa9bf562bd539ac83c8cb445e37badd65da179e08e17ec8a662eab98d6d94fb0ee084c0e80485e742ed51bc3a21cf69909970c71eec01f6ed4e87a5f689f7ec8428791948be361eff66487c7c7823eb74b6c823c88b2d72372a602aa6d068aa8ae446bfbc8559ecd0d336cc7c9d0f75f2e56f7a8a8746dcd6300c0b7f94654865d2e7e7440bc54aae810abe8cbbe0b5d30028759cfd4fd28e792ca372bfb6aa4563831429c2ab019dd2c101a3c2a53f8eb30aa7dfa50f20a9c4a008c8b08f569f195158bd079a49b72a22a51f9a9bc98abce905dabde7c9783e1d92f48d5c2161f215b0c82acc2cf09f6eb3a15796056dde8a18facb119e8da49de5538d88316dabcd0d1a7008baf7d171529c5d439f559fa9f31585c78fef240af679aec69ab8b44054534b74672660dfc21b946532cb9a7e3b790d012d827c679bab212864e78a0d26c843919bc66d5658c46c418a7063f620510c05ee0b236bf6eb32c841f21dffa0a2ad4e1ac5c088fac6b5fb708fe8e5a09a6877ae3a747416e2a1245de37e767e701c31e40c768c8bbacbc5028359adbb25970cbd338a62c8cc0c76853019a66f766ae554cbd24eecd610c7e1463f5cac7bed1d3891787264963a60df01da4da166b36c67ce52fa2a638c0dbb2865790dcac2eda3f53cec07678217d40d01c671f3a87cd121822f8ce6a520f3c4f4c57b84334023ec5057480fb3fb4a315791b7bd1a674352fd7789992263368206870980e44f1b5a86711f8958a6c8a37620300a9e36be1879295b9234fe0f48437a65ebef4d72257c96d243e2ea6edc79b7ab63f1f2473d748a138a7b2ebf7c9197010f49d0fa32218eb7ee18a015e44437db9f039f7e162ed79e80f61258f7591b678a4bb5dc22bd5b24c11265fbc7a1a70887c939026b371290b6645a8fe7b72e8aae0132cb11011ac7a59a65d2cf41b636d2e1e24006453355a142c9efbd9c22534c8bbd2c7db4d8c16ee2a9f1f08f8ffc4f2863a348d2d794acf51d2c69ce813f502a972d6e0094c58f5a11049e3303632fd3f2dc819c95ebe5c65495f4a73357d55487fda3cc9913887b11a7f5c8ac311c38b3dce1732863b3a497cba84b6bdd98a884c8ec4367c513b9b3c74afeb07861d1573870b65be738ebaeeccbad338adc747739b0ba7151f8375e4827c37d87f0d9786de200bc8e466de2e4eca37dbd2fb2a7d814b0129fd017872f0a6a160c5a42074f06b393c3bfd38cfaf274c3778e86cc2eb6aa777d388328fa9c14673df02dad9e66a684fda0196631ff487979a793ff809d2f81cc0c7f24727ad89ee69c69bb44369f0df1e7c256f624a696725f70b236d5740ad2c03f410ccbf0e07d622db7512e522384550c96af83c1cdb831f50f3cb31a7a8c514f2c54e41a267b11f33597e2ada05972d8d2aef6a267ba719970f641fae4e6e8ed086a2a712543278f8fe1eebe2e678cb70b294242af796849a442b24002cf26fe16fced660812206e8b3545f3b995e1ea23eacef1ff954ae787a1ecc13e730dc0ad5eff7bb4bb61dca8d13b820bbe5f0770f7e06fa260bf2600761c188b71c242920cd22c6ea2863bb31fd17777f549161c3e899e40aca06813365d50f14b7c44f68aa6d70f7e892db9363dc4b92147c88e1d503907820682bd5497cbb50ad12000964afcc79576e28c17919a30fe9868fd63ee9bd554db3ed39684565afc69cd79943e0b63e0c2c5ca6b27deea1100bd7140ab65b54913555b29e256d4ddefa8e18565c2306d727622258a8bc0ed6c8fde71fed3a4e83dbc870d457b841d683bf629c0a2a12d9649005d09df0ccb63ca663eb4d82938c5df77eedd0f9bc2de4239a10e4fda5c27bb1ca086b589cdee1b9167f0018f522e4a9f4fa4cca91e3351327fc128200ad1b3c5d9856f29b8830bc77e2ff2ce13f431ad4b8cde012b7f864944c18f8d43a00efa2bb4d929954111ebe01bbe26c18fd2e000201bdfa9713a4bea6b03c9b87f83e730873472ae50c62eb22daaf19ac153ab977cf291f2f5e54c895d8686c388958194c167bf9aa5a3947f0c221014fa4728efc4687d8cc6885fb14f87b21f2bdc4bc40fceceac2840c4ced32f366b6621db419bce8a37fdcb890884c526db15c48d9c4f421c39b01675de8951aade3b1e2ca8611de21be258987c6fd611cdc4c557fa51eda158929a8ec3546e48d3b9b57f25a3d6d826c878d6e5bf4f95509554022a1a04afa6cc2aa2b5e34921444b19963c8ebf29779077ba963d8cd31d28b37dcdfb94bfbce37f5eb694f3407cca9420296bfa75b751e3e0986dba1be7122168f53bd3f1ce8e8310b786c29f3bba05bd6473d0f560c77c75c76aeaaf7a53b0cfdf964f9ad8ba86bbf115496672aaea228435a8612d18e93bedab21820bc22342e6a4ec16c514e594917c70dce1a5746044fe02fb8f0191c3c34a70521bed64e2810559763563bae1f520e2d920d5bd36ca766630088737188a9fd280a5e063f5efb07bb676fe2f87fba68e188f293a0f20bafff91bb4c50f8d96f0494e326f8dd80048c58de3ab1344b0d6ec0a1a22ed911ff1e6b10c031395cafa06d4eff728b0d65622d7a1e7cb677a87f913187e9c73dd1106440b9ae8a0f413aa47e88b878ea1967bec553775b2dc9322e2a1cc7e741f79a9915b3ac7ad90609b9fcc6bf283de22cf3550ac74cb1b62b12e3c65eb38e383e7801af5a68dc84bec83e26c0934675a84a92649fe2148837e1c39964050f473a74c62b0be317efde7659893dcb05ec41c46ac0d4fdb500c08183e30a0a713fb26cb102ea027182fe05446e6c9d197a72a1c9995356f3cb1464d0c60133f56814bfb1e7ef91c4d1a5d9d1d5f790d567429eb436b6b28805b27edcc2b9a2d4e4b64da880bb6630c02150fabf5fb3ca82b83d14123406e77d6391365532a68d206edfcff31730d95fbaa53ec3e9d34fe6c533346ddcdc1187311f894681924e43574f4a1a515f665348ec0f4bef375d7a6fcdf4e13e29bababb7dd98f97a2390fd794eaf94893b933f34a56c8012dbb7b74a2cb691cee8d9530c20caf64b634747f17340e1832cf226f341023209b6e2789ddd22dac8d9f4c6274eb7e48605758ad9afb27e8ee9cf624bc3c846f07a5bd958d665a979d62e0777468e8f9678173357ab3ca31ac9867c677d873dfecaf35432d665540bb68fb5b1025aa206da31d4a54ebfba0ca559a5b6103d82df67cb6962f35b24c009652f0da09948b7387bc68e5dc4ce44e06208defcbace6056121818d7c5a21f056205422aa2ecf4aadcc99a1f3ec0f0a4f6bec1005a6ed537f1257c84ed950db4c777da957cdd581dd37cf352a7dd1142149ac716f05bfd2d047331ae3f5da616524cbaf361295a6d52d1781a93cc6c2cce4297972eeac5e86eb88e93829dd37cb5484fe9f137e369f4b4f4bdb1f1b684d593aea500ea683cf852de77c20c30125cf48e77b908ea92719bc66a4c1a33c7802573e6898da8c441e0170b3f387585cac87c35fbe4a46860df565aeff0314d41c862cad07abfa093a37b370137231535496418dd0bfe0591bb81795e9107049185617d6b8cb0898a691db78cf095fdb7b30616af8e210f018957fa25840b904ae041147986526719fdaf599da29619b7ad312bad4d1074763d0b9e6fcfab48149706298c2a63e9581f1af09e582a7071d6d60a4e02ca5bc1330887ac40a3fbe215856e59d90efb693104dd7bfe08067f52d75ddb2027f72d92e508c6f5de81589a3120986593dbc09de63e12c2ee9a01f374e891e3ac803005fdb0953c221fa2897c24623a88818c567df496d8b76f204a9cd18f915a28e300e3d155ff12e0e2263088f39ce15e67bbc7a350529f3c2097e99afd3f248ebfd261427c027c9d130ce4bcc417f8faa6355b5e05c54f9f20845bcf1c51423f72bc86b2220d07a0fcd6382b342f491f4adaa9735116d9ba13b2c5d1017bec60b417497c64356c9c2a6bb19e6559f7b7261e766b78bddc2dbd50191bef10cf11ed606ff91a8f78924f0e00638d8e98b4af601d94f7695d497a26a5c20a50ddb77bafcceb761f0908dbf92c3e4c38b2bb3fb5c35f74a555b658c8cf05f0ca8df7a12d545f8ea8548f9b4cdc0c592c3499096a2f0af758b08b5ecd63dcf6c6aeaed7f21b3b9ee0542bcbcd23376403657e15766da4b2eb49de4cdd26c85ba08ea027277f4558d71c3f00d70ce322957355a67688c79f3f86a3e094dcdfe4531c7c962487298600a81addce1fc8cae001b035c10ccbcd81b9b9884ddda5ae88ae195bbf8856d2253a3639c30aa6bca14377f59f562ca9c4bb9ed5f40b80692f9c4439cd49cda87d4080882cc61ef52b6f77c122b57345a1be1a7787fb6fea1469dd49559d69b0c1c2b3dc322349d06fba7741eec6b74aae7c3985a30c74dcca070e17734e3bb287be52442421319c8da9d8d6ea547eabd753e92b6568a280762a07e8f83572ef8d46f209890c8b28093930eb1addc7adc2afa0b58828ad9f36790967161dbe8bafa419be170b19e7a3c0a49cce2f0676e4dee44c51d2d3d28d239f66cd001b191c0247fb5323189023220971d1e602e6d4b815d31e563f4015ee54ec99470d2bd1a94bfb49b0b8a1c7ad66da2a6ebaa0bed0a5733b4e71a5192443253c650a6ff9665968a49f9d7983d50e6d5f3eefd96340e1a5274fbdd3ec53520ed8d291807936b232d275308286f173b051bd8448068333e3b550c19f05e701faa27cf57703277b798140a638d4d489e10ca94c15cf4ebc0528e30de3e94b5ac7365a0e3f48c16c9aa2e1c149a76b3729bbf6647348db10c96f8a1542a776e23471e68dd49406b0df86ad8ee78b16d6f9ec5e25f9bfea1a3a019a3e08689f21ab046fac8311c8174585a783841b08a8782dbe2548c325132e510830579ee3714a077bde5f1d66306ccec99f6da1b504ea4a4353c2ff38eec50c635ba0ec8217f02931bea35bfb43d5697cbc9981e75f867d0c20fcdc17708802a94ece70b166a22ec0f1bfa1045e9a224d661460061e400149f2c47fdf45d58d7f51994c67b46fca94aa9b4e339f57f4c00599b14a9adcd3f0e4b4b89869f6fcec8b1e688150590da25e9ed748515405c0bb19c637edec9f2d14e53fc217cb372b100484b07480c82e58ded9d2449efe45fa4163eed901889929f1b92e697e191c583a41c33bba4c2487b8a6c5a5e17a7328e0e450d2d063af2da978b56e1902b606d2e03e6516aeab91886844e78a77ea6bb20e985777b48085a4e272823a526f47b896e8f9c82fc7c003ac57fb0dc2cf9d2d24ac04a87e099960ae919b318cedaaaef4454dd2208d56e36832387448668d464b864181544b2a404fd0d78b94fe1783189910a8a3ef0024baa81cf8a9bd7cf3fbace29ea182d8828c3f46344c3b818d1e29312096e26a510954d85cf02968069fd5ff3e59d3ec657b4738ea920a045cbca9c125b6c6291912e7bead1cd47dade80b4bb110777601f7a2792b1495ae1e9ba03a69bb88248fe48c13d34c3b86bee7cac129bb816725f4629fd7e0723aedc473608f292d1d2b7e97bffeb7a156b79eb819394a5e4272c97810ba2f8d78fcd8a6fccd27a139aee5cce42b28eab806c392184af3016f0fff655da58ac2e0648a260931a3efeef5a6bba73d3702027d4812834a569c262efa8840d0073b34f433f3c585e50e61121799cdffdc58a09205ad7fb0a31c104bb54e2405356bae2034be1215fb89adbb4f404d3f5cb322c13e3ee6ea93212b926324e6f5a50c708dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc73ca6c966d536b5686cd9721375070d49f7032c716312451fc2aecb506674c5cb0a40951d2dff8ef2e197ad492956813e3a1661124c68125cbe04cc7250803a3a179b96547c923a92470cf0c1f0b423167fd29dfa383b23be75bb0ce91d5d3c245974e889880b9fd1be27e0dacfaa4dcdaa19bf8fc978c2873f498765def0be7b933cc82dedb9cf7dbad336b111f78adc2760124d9734a95a428be5d6147079a58e8364cf5aec55eaa23ce4e98bc895073a197340804c851c62845364b3309889eb0398f7c4a18848341889cdad510000b3a233e79ce41edda55a9845ca0fe25cf1df4dd076800222212baba028210fe4db2e40875e5bad454de7bf17b4ebfb109ab239793a8cb1743dfb4657353b7ef21802042df03daa66e004acb806b6085f3e172a63269dbdc706117feab8e6dfe2c639da2e356b8c3646b0040ee4d3f6b7314dcdc761ce7cc0c4a3956df8a7cb11632a221fdb33570b2ba7b413b2e414ba6cef5812ed165b2a7833ab6ae7ccb552cd3f9af5f63791f5c907ac57f1aa377ae13f211df2a0bd8f1ac2f75fd9c7b534f986ed199cc626b8c09e54bcbc2d2f5a498c9fc929bedcfaf987af4f801eef36fabae15bbc89c7851790d86f519394eab8b2115f1db1f608409fce8843ff57ef4d061441528d6eed52f6caf806c2a50d4c437c8d3caf5c91db4c33ca9857017c12631a6b6947aaa5af18065856d4399e701efdcd7c14b16d609be1b1b7e8d1d64f78a86f20a127e87f1048334cb5f33f733df488a59068b2f9a66167d80605d8209edb8663151db6fd2086e65d4d9ebef2658b30bc65d1743fc53731686fe24b2428fca24e3099d2210a713681ad263f479b9abd5801295f5eb187cd20440d42c5eb27d0897a2fda6873ebe217915c9bbdb446187a6df80571f8e236b503fba2728b65555d5412af20c411ff56711662506587c337fa19a7aedd84c58ced1e920b733aeae9d76f4d8de87669712fa5dc74bb04dfd2106c538b2099861023c524fcb0c63a51cba87719b8f6a36639ae5444bb42b8cedbf804b3fe17ed7de5d8281e867f8d3f4513315512b55e51cf74aa48a10cc6357ca81cc6decb2b84fd4ecd546c60583c5fd7cbb50a15deeef92411fd7a3008049c67e8bc21b821de9d54018826dd452c1168cd8b79fd4bfd6d65b00647f861bd338262743c960690789ed7f343301ef1a1319c9bcfd8448cbf17e32b53abdd1a52c4ddd49d95db1a7503cc2f05a97a0608d68bb855d33aac4e984c8e5237dae090858134cf2bb66a957e22310b37ae5c0585b375e460424ec427668113650c22af56c64b405b6997490c6c0487c561d0ac0afbb4640dfa7ebc951e78142335a383843c909e2e12328a4c5ab9868231fc672bc7187f9e1317da49c1e88c79de29948ead09ad4665c7f26416670dcc977c6bbcd4b2cf61aec188a53c0e88c8a7498fd079b67f9e95175b7bd351b3d836b46c7cdbce797ef56027b4449715329b5f15c7675dd7067e26fb907029be74d163ae1bab83dad27d13de8bb1c9c59eb1532e66136375d90f3dbda9aefcd286b2e8ac5515607d81a0553bf3fbae36a9db75aeb73a9e340f6d90b2bc64fd85ef86a65e2c276381d0156c269454bf873f276e14a2f6f8c3f5953b9fa185db7ceadb0c4fdd1360562ad06201969b02e130a8e290d360ce0dd5b8c0d0535d965aaa7019d6dc92198775460b053e97d3b147d61d697dad4648792c61cfa6eaa062d21a3b42192eaa65f87c8fe273a635c6895c5552ed8852e19ef5d97a9e77bc869cea6813858a5dc5b036b432ad5cd17b1b922eadeb875a6397b1aa1c3c28505cd3b392b77d48e30151983527f6ec7ae79e25ba763ae7a45be1c8d02cfe5b1ef9abc098b9c38c437ece95face1cd82493f730665cebc408a6cd97f697b7aeb17c55fdc817cf16aa9788f42dba211f542ca982853c9f6ac6322e9f3e10ef202617ff7c60fb3df76c3260c98a973137af162a1aac56e7f376efcce181efaf7a04956592f1d81531bcb77af5ad4bf0ece2315c90239a6fdea28c47ac77e2e301026959bc5b7966fb4c703faf7c4e7ba619c0c3ceda51e288ff9b1ef0e014d387bf43b77974acf2c748414a69250cb31b15710c17ab608ac1ef2da6ec332beff08e748421dd24445bd6319225b6ef4211a5515e0e3720ad9fbfaf2428260e32142e64f4523610a1c6b38811c82f5fb105a874ed9330512729d988ff5503e6cc66d79c61f418a3ddbf8bfe439038edab69ee03f7a28d13729a9d7a87bf3e90297b55ece3720fb319ab36edc3bb3dd1ca10f0bca5a48c7c47522dff82c7165120c300eb7804419952cc6c9055dcb0b864908c42db3a3c4209c0605d62769a8c701770eedce68764e3158b51b3c90dd96316e9a5c188067db0ef40bf31ff86cffb1a1e351d983352d2f0af84787d424596a0fc55d7278b3d3379925c3c9d491238e7b53e82627cacd49869a324329424d1252011eb7d0095fbc17bec9f8e58ae65644b7c627bbd8d3c4b921321276ede6c0c44dc80af9696a5554c2d9a0e7767f5e19ef4ca4dbc602873db3b938eb0a044aaaf713a23c30f0e450dc9614e835b29b00ade9587bbf97c70b31b36a1ac9f088aa4b7f52f1d6fef78d41c5c5e19544089ca3c3620de3bf6a06f976a10cb7a2cf960b48d71c996de8760f799ad1491c5451444a31f44061068d88b0ae32624a4baf742912299d717a55b4a3ca6428da7074764e8990b7ccbff97d8eeda47c846ff0935fc52278df116a600d55ecf00c7e010d6626df8ead624faa9f56d5c40c5dbff1a7824f34fb30856c03311a3288fe15a1effe007e252e7e98d9d3e8619c52946e1c7e6eeae55f67365a0fbc036db0949956631f6c91af2d6ff1ca1b3012ff14d384d2d7efa3a026ff412514fef4d691fe977ab5b8688139f36b5802e3686a7866d3b98c8321aa956fe08dc25a275347b7cec88c7ac28c0413f2a5115134d1ad3899f625ea7f79c42273476cd05ef454534701bbff19faf2c711d6b2c628f59b8426ee68282d5cffd1dfa761fbacf61b2d0782b84a58e0879c57e89bc5e13c4ee973337bef853cb315a1805951e85897eb9713352fd41830377ed6e700885fb80242a0dc3f94f6a9bfa53b8ac61088fc08b60761a6a07fedb198018e890d124ad3bae4d670ea01744a5a6fdd4f616510dee8064c760915a045f635eb44479243396346f91cfeaf634ae284a0c1f35a92befab6b0185bbbf776826974b5668a844a0c9c10a4b2a283a92dc5bb4615ed9ff60d45805ae862af09bf97ce5cf18d94813acb1a8cfc7542d9ffae0989b154670105ce0801dcd3ad567366a172c57c7a339a6be353a59796bf5bb27c3e627cc17abd9160c58b914394cd91dfc6c5ed24e0c17611a17a161de0bdb4f4466965e047f88d897c1e379629a4be194d308dc7ed51c71462680dadff528a6a76188b923f6036077881883ce1f19bf303becd77eea347fade9dde73f4ddcb947a85d98fd0dfb34a7720adc24844f8b2dfc1c003262fb637c5abba43a3546be10a6dc4ddcc2c74514fa0e793dce76e1f323922be643fb5af8c3681f07f305b0fe19e6a200eef8aa16f809f973e60740c874156812bd972ea63c4262030f0f45ce88eea8dff36b7e4c613845304b20be400a5558e2fde971dc4fafb85cd0f0ab609a4b7555df2263e7ce6d15cf2f07eee9f28d0ba7b28abca57d3b0329eb4cda18de689bae3adc6b38c41787e8fdb3381a883ae1e9d99383bef063a6d06d3e4af6b14a99dce677b118b426512094a37df9a076b8a3c73abc37d0db4b3ff6397f21053a2918f923141bf5b15827056a4b6ef808edb8217199483d9fedfcd3767c864fd2211ad10069a7dc439ea3bd01e4b1b35e37a2133da212a6b853a94efae25f459c5e20b4d79def1385964b554c947c390078efb4cc4f4fa79aa574545975ab0656ae4c13e488190b591440e3cd97ac348631e9994743690dbc9767e396ced7bf6061baed37e9381ad094457267d106f004462111ae93c94d34b2dae561138de6a2560ff8973956b0bb7d9a0de024af0227d080b73f8fdb1d34afcce435d9c50aa0f3af277ab4e183d93ceba4390d022a5c42002d742fe29a109446d5321a2f64e2f842993d000d29ddc28f67ae6a6c1e711f352c5d9ab7af6b7a06614b028a7f6bab9c67f9021860d5feac4fce7d0e7adce8521fcdd4334dcc5b73b9761f0a1fca1758b9b415a6662b067bf976399979bbe38b6a77e8e1b10b1faed138bb139a97b6dc243364ed01da5cb53aa0fd7b1af2a2a4a58b888fb07deee60206052f682494063d9211f63326d9bae72dd6af4b810204b54c9c83829cd41033c5caf820205ea7e83c3dd8a14437c0cf55e2b199fc5763637b39729a08baaeacef73897d02b1e1431fe71a24e578852d9717d6d9c272c3f291de4e3d25fd505891b43d7208773bd5d8ef945e922df2ba7a608a7d0f4d63eecae70c5c2ab7f18dd659bfb35559f727cfbee60d22672493fa5f3a0bb11d05061d73c94a3015702750d67d237462e6c272185bb63fdeb9b952695456ab969de952e34c0fa0f7da8fe5c5ab64987226bdc124d0cff84c09e236850f3e41e7d8b7af9d9b9697783122715347edfb9fbeb43b6cde1c244212fef93b84a0d9405db36e28417e91852168bbadcb4993fe5a8f8169cdcf7d3eb8b6ab6048b634c3c188e7b8514e9400709b863b31682ec189663e02d6053f1e5e937d90c17b14b047bc67b030ed6a8110a4c53d235c6209c753fd02260e60a81942e1aeca19cb3e3b293ce762c389bef711bf19d1d553b340c457600c2696ead0b198dabf99244cc8e7a044b8fb0ae53901bb14b271e3539a7423f6ddeb34e6c7da7752bb2c4b29df83a63f3301db510a4620bbd3c0111f2ea65b84103b7ea13270d67ed972a3421d1f43c31f7ecce1c265a3f12d4f28b91fc2caad7e98a7741c056bd803eaeb8d647dbd73a3730fa926cab1a99282d29323fb8422a0b7d0bdd88056e7d59fa16e99d34a4ce294cad0ae6f0e43306807e30d954b040955f9c5a13c28a31f2950020f31a64d4c7465b938bbcdcc5d342cd5b01a9e045c0febef12767064a793692dd52c5b0bdcd57afc6c1af9bfdc34435978fae94f8608babcb6a0b2a4def1aaf94b2b41403146b4a7d5018f608d7c930530bac4dcfd0319f57cceeaf9f57076fe485332e68d75dc220850a29dc4f17edda7ae9870ef558fcd8a82d36bf768239b0e8e757cfb6f0f37d35924aec1325e978417cfebc733bfbcd23b0c0eafb8a11ad7f56d6f08a3083b4d8742951c034a366ce3a6c3ff6dda86b93d948f81ec6d07190cc890c6f00b85f8140945ed23555940a464056381f44ac4b93fbe2f2bcd0cb16ca4170344409b8dcc08b4b9be337bec6ba9e73d7913e5ac3ec0e508f978ad27ce2b83c2743d45d94e268535e3852a53649ef189fb299eb805b043ca97e7e434b221fc1cd3dc7a8bc7076df28be4a057effc719dc5535fc46df3f6009764a63047c3129441087eb8183b38f59ba4435612e9d2d35e567e7b8dcbd557b4fb1ae63965c3430ed46f0ec1abcc47a415e20dddec9d49cab0ef0c855ae8f2a5187cf762ac7dba2fca48798b75f9bdb68e99fb99a9195e03a993071f7ec84bde1d7a718e5d7f5f50e1f91084b74bacfc6c76f4d24fa0d1c24b15419da27b42367dbd20510ca239b00169c75f41ebc68ace1553f15b59a682fe405b69d6c771dd4b4d00041e618749b4dc107c9024363c8ade9a84ed26c80caa70ddde6cdbfdc757;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8031d7f12fb0956d201273f9d3c5804f049d101a463ae4e19c80414c7cf29621d2db9393cd30a4b7056fe0c98c66fe621cf594d8e00eefcc17ef14aa1bc392900e5a2b34cde2c3901c62e6ba21495310ebfc9c75c495d61c8c800f27e2bd9f37bb8e0c00c2dd8f58ce654ad7e153e6a77d54b646958668800000a234404a557e9b75989c515f352eb1100b1bafc491396616433dc187fe87a0f0102edbfdea035d2233c051226728df1b66bb25d7d910ccda14b8151b6584ff30d6d5b577f41334034dfc24c8bc94ed16a31cadb83299928c117ff5743c901be95c74c5b3ba2718372900d1c90d1e7d3605130abe15a0c9b87da359d93165fc96e574a4cdf3ed11180dec7e58bbb9ecf16648e52533c2dd8837fd1bcd07ce63df8b3dd9c8aeab04edcf58404a57688dd268098129c5596d3ec77c7926bcef83181071e6b1f20e68f8bb53befbc20f475641d77260a2f689b4300be5445b9b00a17e5dbdb9a2ce244f67f0bcc18ffaf401b2d7d97575b2aa3fbf62b25a99fbabd395f0664c061c3a3dfc99ce0bd2408104412e3d802c40c484090f9ace6a5e573efb20573da401aa58830b29139a9e9c0947a280ebc3990801cbbdc06861aeb77c5b84d546f75df37adfe4758aa5d845e8bfa618c0b4dd1f4069600e278da7eaaacf294bc1f691eff1e6018a8dd62a247b0460b79d00f0dea0a060ef1d52e19ae77e8f7c39344cf0de8af0a5124e87f8bdb61f18df938e85e5d6427f0b720edbb0c3dedea3b742bb068cdf31ff0c6bf1110fe7fabbe584a6bdee59012f566c3275af11dfae9be775a3b0b8b8c857618f37ef319a53c45b166c8c2d8cdd4c8e5b6d2a786841fb3d3b70c90811b398df79533b98c2e75ce78b26c6d8cc3fd0d613d64d14308b8558a228f30ca5d6ce57d3776fa62dbdf8b08af7edf392a371460206d936c3938234d21280bc6253db1418be60547cc5c997c1bdf4d7cf5586b902ee96ef811e4c156b8a78ba04d9de27d3331142695257ffa3e5880be83e385cd32cdcab7372f780f44b99da36f4e167790abe8c26a86c682e6c5433fd2459fbcdf126b0802453c8bea8a0f1d069cb0f34222bf6d812fb427550113b58fa83d1a5c7cbcd52b2f14546441082a69a2fef424949510890e53af131698f53eb0a48446086edbea0aded97fb1464d7f545525b58e9523df926962912203fb881baf4a45a73061014238a3af6a1edd6c8c29294298238ee8dd97b3c6fc8f936040e9246f4837c886d0b4385d24538ee265f5cd4e6a69b74d0d8157e60d8b5cf811fc35599716d6fa02c700aefb0296570135affb1a11ea62f5cdb65791abb0447b3336131f96ff061f5302338ef5ae25bfefd44b94ac0c65248790ef5ffc45289daa07f0bef52747b4d3251d66cf79b4aee71e2338a948daa052b0c94f7bdb69939898dbd89e6263aba21d3363e31f5412583299a7b2adab0f54628def2aff1b83dbad117d881a23751228ad2224c7b643b1c461367fe1b9da3504342f35eefa41993e146bf6b943ce8dfb53828cf717754acccf09981652bae22cf3e65ddf8359e752cd417cfa0158b3c8142cd60cb2a4073ec6b0d36ab8402a4ffae5678a3647ef2441bd5dc92bd1318f6ce582bccaabd89b5eecb93fde430a8c8e354abb46a2d8a12aaabde0530ba34972c39ece1a8b62efcbca970e131925a927cf798855e220d4de10ca987299c831e078dcc967e61afe13cd00532795fbda760c615c17b7041d10bb9fb495401452bc3bcc79def9676f6c6e46ce03d15885ea641061a6da858d51be29f5b10cdad0e96ecff92a816084b378c818ff72bd2ecbfcb150d36427b3e98075c28cc981f32e951b2783f8a1aa818079355fdbda47dda5831b6e703066ae7199c322b7add6baf4b45374d1fbf908bb70a9d772b64c361b6beb9461c8d25cbc50cbe1a015572651e090818062ce85c9fe9c8a99ff62438331166e377844fa792731c78a1daf18262e2b4539276c8cd0a345fb4649cbeea3c0684a5cddb77788f2a776b1ce8da8f7a966c5dede82df0f65069f51df3e613d3ab2beb93d12413f0339baad559e6584827bdbf2f7c7454a12b3d99429ca50bb4bc0e669c0829cfa1b924735a82a1e3d96b26ee438a1da3dcb359bba5e08d06ad67302d36d78705124688523bff72b2567a87892114ea83efba2871f0af5b4f4400ae181d04e69492d89e020a4a4e45066f5a4c2c34f6a1680bced382082ac08b2b932d98553777aab3ed6e72bdb3b06613f4009aa02a367027546bc70c33c468a3fd77e8db880b7a9b2a32c64fb84984b8da58db362ae45c162db46cdc9dcdc98025749d6dd59ed38fcbd1b5e2f67cfc1164ee87a9f1d6cbbd33eca4fd0c1509e9a9769b8822ad322a5c0b40b281c9227d1f1159182d4795583d556971e8f522981e611e981ecae803e86286738a625e57cac8ee41dded96f39e11c4ddad5f0792858b2b30e04c2c40ef47386b05fdf092b25bad50b7ee2231dde8805e649a031e3fa27823e856d369219131aba127680ec6b0b19e1ba2a6ef68caa9ae29964116369ce9756fcffe7c11fe5f70dd8ce0200751c9753f1129a1ea6067da5f2e59477e3b385ee0cc3092b9b690c83e70aad8436caa9f313650522a58ed49998665da29da2fc1e2722461b18ba353efb3302fd80c6d3a41b63f3f589ef0c846aef73affb8dcee47c5cf77fdaafff44fcc5c3e08b7a00644b441e78b7d0ff9fd11801a5a3eb8b8a7bfb0f57d19aae571151311ca43778a626f224d64683ed5f88b886b063f26d2b5799672efce43cbf47fd7dd1707f27de2a492b92c4cfd43109ada0515225c769edb0c22524b0296fc78e21ab99944b3da10e83349bc1ad0acc0ec432e3403a9b0ce3fc55fc654d3123408311472b92f10fc90f1021e35f75f0be241750b27a36c7397dcdbc900f405e897bc74a3750c7490c24cad0e65a43ed744430941a10b6c5cd85f8ea9354db31fe291adc214e035a0cecb5575c193c730fda344a467b14a656ecc6624984278487c54f73c10d19d20ddef24809ccc9feb1ff0df49bdc614e595af9df7caed4069d5c468fc973e541676226118d42725b7196b888297017feca40c819d540d6700cee7f1c00fa22a9c73434da7255258896faf9ef9615abb5e524d3ccb2d0874bf1905eaf3fa8d4ea7b61dcf4c8f468c7dadb7ec6ef427a15c4a06fa8564e3086f7608ea17606b7f714696e6529adcae25db1f9bbb83784068eb0e71142cf1b9a842807f0f9fbe10da486b29c9f9ae57a1a9ff94982b08a6e61e45991d275c3c4ba8ff69079eabd359cbe5c392c17383be6574dd9a359b491e845c6f3602156008e9cbb335b07bbc3b2bb3a56b7382432d25269a668591f825e538691f41860aa8976322f2fe281a9e2f76fe5c92a5c44f20b67124a99159e8074036d402cd96d6959a4973cb5099fdd470a20431577d4de73abc71e7695bfcf2137d508aaafb7a6d29328312865d777315ffe627bd9e43a538feec6f0c2e047840baae9392f5ec26a2a77c5c6332399c65d1ce58391cc5925976daaf623e5c4b49376958b1482e432472000b6149c632c1c103afc95325ccedf484ca465bbf0372eb9e53f88dea2bd9705580c7dbf7b3d843795f133eba68cb45561b8f75efd568295ea192fa505b7a910c1f81cc41c2f7eed0b64de7a82e51fec64a6c6163338a9320f41f6ed3c9f7021d25034cbeb7b662a0cd8634b18b918e1928ba5008a01dc346ea3d5528bd04bd9c4ae87be86b443a04e3af28176090f914f686cdeca71c7ac2028b112a10b0d71187954ea7f3a0d4101a5c68c5bacbe524daa6241790cb66c93cb0eab783c1d2973edda07cbda606348b797a47f3943d3e54ab3e6045f4bc72d8ea0edc5ddc4e852bfbe1426bbd0c647445259829d3d4b484318359dc4807ab5b92da428479583d46524ce324bc78b7c5caeabc00791ddd8eebe091f4e78d8aeeed109d1b4dd971ecf4fe640bb602c270dd88d7f24e38d5e844cb7663a628f4ecf5b38c423adaa8640325db131a835a3ddea0bd4c523ef1b67152c237a4957968adb134f73c52888d91eb1eb773fdb36968c5ce7338889b4e400c6683bc71585c5b90acf18336a16904b33b6fc22b6f9f0f51d00ec1c0632865be3dce55b4ed70bc3a59c83d4b492ad264e0f71eabd12a21959f869af7c9f72169f48243b4a70f783f7d00f32ee5ecaff63a0e063fdc656ee04af75adb1da8ee1ddf83ee3fd33698444a026d310607443071a8951102024147b42b9ee2a1152130375613cc648babecd03751d96e88d9555babfe878a8868aad8f71bbccc109fee114a7239fc87b9322fec50f38910aaaf0f5bda55d4ea368380d4a701707ff936e68a557fecadce0eaa37012a4f47a03feb8a5b75747f3bb542975d682c1b25a2b3937fdda5a791e497234673c1dd1168a76aff643c3f95378c9dc3b2a5fa0883347e38d2d6bfbd594f6af782e7f4f2e51812d6ff5a1c79496dfefcb35bdc2d2cffbddccf1a7a49147ed30bc242bf93d0434fe6704a75f18b130a367c1bb714a88b22457694014417eea8286dc6888dc9631e0c31750721be2e3ae0fa3172b1a93dab5df460aa23aee6da58cd84d5a5e32ef7d7449f9e8acb949eb76f9903a7047d754d1cd47adaedd6eead99d2e4f2a17a1281d77c2d1df21962ee18b5f132c9263c522af08f29c8e983fd6d81224da1270bad0d4a11d03e107c77d0f632820344915b7e6c5f73ea8df812cc9bebd4e0b68fe463054d1a0f56d57d3d4a59b46db6b1c0208214126046e5dcd427c87bfa50d5c84c7b09db1d6b911be8bbc9fb32be5655022b0fabb9014e4736903ef39222aeeba80c7311e02874c63ccf39eef4dec74af9b9966ababff50f2d6e2e686874c0bce8809431da169f9567440411d9e0b20546fea7f7b849236502edd998846d93957f5a75da02e8557e6fa1cb3e0b5a460f585be030b2096a9836d348c3094e47b36ba3588dc2f9ce2c55979cd9682c6578b4c2d0df52c3bb29fd2d5d976c023db720bceed1725c56751407051e27a365fa24eedc8a3d2a937ca017cc82835e823c34a89f06b3f2ae85d68711ec8e205294b6b08ea19cef86af3f967bf58b9105914c2077eb5d32b1e3b799d6a66788c503931b0e849a32f0cc70132d974e08e7323c23dc31d8b42b13cd07ede149c3a9c2ae444e9050e92d5e74de773f18a48e145e181fd4cb8ba07b0951e0c5b3df583083d5fd61e9b492c09480a9977b0e32ae81eefe773b2df0eb4a3a13528b0bc2ac9428393de52ccbd7cc92ddb63ff287cdd2fa9ad3d6f47a06a235262e0d945a6b1a5598f0a31ecd0ec631edc4931b9b76d0016ca08af99f1d287b37dc4a3a6e8c9f99219381b200ce8862057b84242b984b7d423620a72f10249efc9dee7c9ccb059a03828a82b8ba62deb01e7dc9c8b169dd82be427fb512e95ae4653b899bc36db4e34f99a41483ea25314ae27d3e1c03d63ea3f6d4ea9860651b453ff9c34db4ed2d87add3bf8ded02fe93d22cb410f98b5bbe18520b2a00a436941c76190ce25de1d366f71ff4f496f0157aa04f10065ef66afb436e868a4f8b03d509d1df419aaf350ef9f1d0616214341c4402155d04432ca39064d526d78a1a05935de94e5d69c6ba12092db15f10c34997e78c5eab4f97c36556bebde492fd40c844683d8bca71e667d3a7507ec5c13dc0e84f89a70533c8876ad85472c738640f6b95a50c8837d8e1cd269fde3d5ea68437c953facf3b2592e7f9d25543316dd443fdcaef2dc2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h43260e3b55a49ef9835d2c19d912666892b476bb42eb4f58a6d14648184323ef779e7816248e1df010f37472b9a4b7a620e34e5a2a3754fb2f28ee47893a23781b1c5b1a9549cd6b2108faf338cf1e1689aaf1777dbeb8e013bc53f71a82bb9f291c4674f6605ba985e368fd8bb2d084820317af87570c2beb06238e3366b451cdb872cc8f8a2f09e0ba1f0ceab7c07cee46f3497679f2b8c8d29279cbd4ce9ca66c93b86f254a3700f26497905e996b417ce2088d7807d710f16d5f9130f2729d06e0049bfa6488798188e9898271d4588556a8258560227d53f49a1329ce725ea33dae1059f79b99938690458675e85b6d3d076ad0d8fb6e17c5c5ef2e763091aed708527f7a6402e9407082bde2d5fb0e4afb68cb8dfb9209aa70c3a84ce863e73855ca96c1b5718292f3381253825478e50041597f3ce76c9c45f85b311f491043eee320ea23b58bafa9a6fdb30da0130b5e8318b80e6ba68ac7d85ecebeaa94ff42be92dfc0f741375a95ea5983f4f36598f7437c667dea4407feea2e0bfb01f250e03e7150eea7f6db53dd087d139312d5c566337014098ce9bc0892f2a25cfa70e7f9062a0a8397a04d6e883a5a27bad680a220967c78fa24b92a3eeac3a998c2f64d6d08a1b755acbdc5eec914cf96c59dcc25c0d02bd13a6b3652a94e14eeea1cf4485f39c6cd94b71cab3a0e7d9666ca5a07e4a145bb9075d26211fa80f4459e9505fe18c60aafadd1efbc7ac9b8f66bfa5a84689bdc608d14cc1de0530efc8162ebb86213e27346434efe3f09aacfeaa715f49e38ae9e19cdaeb55cd44c6759c1e5b7394c2e07ba0418a49c65e4ee1122e07071cd5dd5fa063036459007f53c0c3d9a4b05efc3f8d4edacf2cdd3a681fa1d71b90bf0077802240d59bf1a543b646e0383b05f1fc272391bcd993682ecf1bf0adb299e9559806e9b689b82c3d35e89171bd94db997289d1d0ff119d68bb7f3b2fed89b440837cd6f783736fd6ea2d6a32cf74f2ff9383adabe4a50e100150189dcaa6b75d2b1dfd99834028ea743b49e2f012233355d5dc1abfdf606350faeee9228b350bd07fe616db22a33b9ff77fb47e182a283cf0318fb3829138e51b0db0718eafa61d2b3279523a15dbc077c729d846472424f72fea2c3438321a19d02baa5de7354f758d217581f6d340f132b450764d4a2f5945632fe8d3ed8b5059f4223c4423a726f6f90e4e87b906b06156b1c994e9813acb41e826efebd12212635db9380de7eae62708c5390fa8d6dff9d4124cd4c9730ec3948dd555ccff9e09837fb1d4ca73c10fe17e0e9581af29a658c6b3746877383e1fd6b2b6dedb502af6a06470ac46deddd86266ca6a0e2c3c5b25a8f3c3812858714bd76c3645c606a6786ebd0c48ee0df8f3c4aa1f43cdff6ad51ebd4c45fc215d62ab922285d025a4a80bd37a98ff6fb8cab8ab346f647607cab21931b2c82405d9f319a8721e446b0cf5ba9917f2afa9990d2813253df80416ec42b7bf5a21beed229810b8995e5e98e41edec850d293de02ab81f4a95e933c44672e6a5a1b2c8cdd385b41a4716c71b52027ea365a93dd9c5b92df6479ccf8932c2612f5f5761aa6d98adc218f0660f78feb650570821eb5145c6b4da4b4c579292b68d5afcb21513b2757da8544fdd6a497484be827e74ddb2a8942ec3743cd8fac3026db9c713a609d3e331bcea2c80dd5d7e86e1f223921d1a26de2597f1887a45bf6cdd16a5d5d2359ee5fc6c5f957f4793d72c19737027c35bf62be9ccc73acf547d40e89fcdca99a5ee427e2a521d581f7baed5b7b8500e23805ceb9127b10b506e18936efce140430d49a61376363cdf192c52005f25be833914aeb8604ed63f131693055f3e1107228203b49d7daf0711a2784460e02c639851507d095ce881b0719a2d4f8174085fdd83793afc6ec8897a3908f8fa28017078bab6d9e87dd9bf210776780370993156eb1535232c499c6ae5fffd5d35b630b128311d865d9077f9913cc6f4e0ebbd494fde626a37891904edda4f5ae57bff460662d57ca2305e7b4d1689ae02007809375bebb0a3993c0e449e9b578adbe5fdbb8b1f81d0d14483c45941cc0933cb12cf93d8fde34c5da0b360598cf02f60fe8bfa18711ae429da7c7c25ef1140620e33775fbda63d9d03a6c298da889c88ccefc9389db0777ffa785aac70ece5707acd44ba23b626efadc99502a8cd0c8ba42d7e93071c592e02b479ffd480efcb87ac99fef7b3fe8a45affebf82efd6a735d2dd0afb41204e043a8bcd65cf6223332733b11e678891c38611b89db9b69e69e21f66663c8a991629436f497dd56ced654a331cfe952460749c7ea73437eb919ef00af7e82470e9caccb0d64622cbc70f908e66483b9ad157b962f47f5ea7ba959ab5411b339c778ae29b1d4cbaf1809b66e82a86cb957bd4ebc3c9562f1da7370d4bf2fc8cb8fd19becd0c5ffa719056c7b12b5360ba926d66c2adad58845eae9a440398622d09ef27f7e4cd3d6f39510455e6f6253a944c63ab34f5cc883c4a81b2cfae93d9d40d676cd1ab737b24f91a85d97b96f3865fb1460704931a842b2809d935580e5f549c08ef38aedaeac6c121fc313c504749b59ea0fcca1d0d6d12f19ee85c7017eb3f23394a8010c3825b51eae4300c719a9d9d3e903e806bdf795058d3b309ae07f68b33725739e6e709a7b13d2ebe6920096b2877fcb1d482b00772a14b9919c34c6b64aed0286983904463b6a56047851b08ab7904f9f227b04560237f34bfb1b1f6dd4b39b04e04247aa1594299299b3e2b85371f0f4a36b36f05886e3cc942f07e2551e68909f55bef8ba918b6092e70ff406f97a6f93a7b92f16dfc975e4f85ce63a605d54d908735d3828cfe0963c6ef88b3ffe94078e44cc21ff1ee0a2cc3b3dc51784f0b69705a7969187397837faebef577a1c1943d31a167472ae84ff535bb9286cf4ba3b0605ef25795b68b540b6707562729bcc304385c5d2e69a4cd968c3d4dae2cd4d6e42fde098190c3c88955d4ec746b23307acc300a32fd3cbb894be185cb0bf2117538785199c14433b2923837dab1988ce841ddf1df24c496a071d2194e373c3f86beadd022e05857d722757625f0512920c0e2ce66ecb12b08e0c47acfeca66eca4954f9f62992a00b73c9049852e70527b4307e134eb19f8072efc8a3053334a27e6ddaa0f3655100aa5064a34e8d0a638d238431197db9a59cfcc16f3b43294186b98b9a98f0b6a92ab78ef48efcb64c692f100feebd00193b18fc043a949ccfb548768b498cb74cb775ebfcdd903ef820415caf6720cedf0319e87192d8be2babe247a5476ab385a5c96731920ae5f49f3bf6d8380792bbd2e3e7d5cf09151ed7c2fa5a584f1dc2314fbede7f1851b80d66de27753b0c967ad6347de370cb8923480b5d0f1f7c6b49e03f85f94f4e47043ac67a4a8eeea8f4306b25e6d72d703860774a7354e47c81c13942f4e82007879453957c995ebcf55f9c95d27bae766388d99440add116556e2bf3a3a46903c09c6179bef7a42052d7627545049596c8130d308270ac132beb0515b00c7535ded73cda2be86f8d7c36a0c1bfe0abd3e95ae8fada37368af48109b1c020983450176c8ec8e22b6725de3482049158da1933e8dfefb0d197b8a9fca242b178319a449c6547a210d5b2ba910fc336952073e30ea6323342973ad8ad78f46857d7f7f994d2ba759d2a42280e2528c756ca7c532db9623859c5a4fbcbc6815b94cb9f537d04a3c35d28d3185e24df91349f21782d65bb87fbcff0cd4475d40c7c2c55f2430805bd7dfdd579f3c9b393bf852b3020cf808fe340251da05bb17f081d6157d10ac92715f761abe7af07daaa03d297729e302926105eb64fd26881ee35e5acc44fd342db547193619b7cbd1f324a8cdbc0e025e6873c236136951fc22c28a532b718726f145b5c7fc8edbd34263afe5e02311514a0c49e43e028e8a55134c10b88bc6d54e615c7a9a0964ac83bc72f8618c9f5bdc9a410b393017cbc3750da9ca500b780dab0f20f413f1b881f4469c862f51f1edb6192bc298bc56bc847d9bb39537a649b4c554e7cfed205c285167f551599b32b1c639e549f7522b79df5ee37e137c3de80117456c6afd8c3e2f4e7f9619c69035310fc42039bfd225091df7e583e7e85a8ae362d200cb9b7d2584289abaff0cfe770854dc70e2c340a0e62ccdd3da523087bbcf4a831bf7b00bd143648034960a1746478ebb0529f7d2fc779c4c66ebf6e8d4d220a2d3293ed4bf1fc1a413be4c04a7a9e72f0d92cc76feb7b9bc2f24df845402c7bdd778ab9dc7ba0fed9d8d94d764be651b91c73b46f9e3e0cdb922db8d72c53c0604c902ed84f5913b53439a4cae76943f514e88384d9b1bd74c83317ec06256562f0d631a1ffaac660d0c98806f4e38fd76dfa1ecbd16d3ff55ae366b8047333bcb1a8f253b48cc26448ae6db398a5e44afa17ee2ea200219a7e70ac2064d4c8821499b9714b12b7df097427063545efa5c7223cb514db847152a5aead9b7432fa587b44420ca87d4b8385ae3a551df21c87fe0ab71efb687bfc91a025c3f192eae7a1b2e34f0188ba5db10c5b0b16e2839f6d0aa35b1186e3065ba528db5166bf873a097c6553bd861e661565c93baae9236e5229c305bb86b6d8ab6600ee2b2c3198a965c7a001eb1cbd3590041031dc7968b9b59232a41ea1d1994eaa0ac92691e324b63ead3469628e36803098c2a263d9e6e7e818b1a2675d5b3d085a38579abcd8e1e8bbbc829ec7f18c3dfa65496824124849c62056f6119a4b9117b4325b78355ca79bce9f4fb7991da846a481a8c58d63e85b9f98828cbea78b56792411a50f6e955598b57749dbe2bf28cc0ee5776a50578bee8ba3a7832e4b74e8d2994a44dddc1ff24c64d0be5a615dd99aea3d242eea713f9aa9314a2fb39e863bf7eb3f17d3f448605990f7ef131355617198d5787b08d60c865a004452a2c43f008a9b29fcdb7aafcc3819b1d792422d82858e30a5a5a68ceb058986aa80b957e26e1716d7a02593fc9d03f113c096ee0d3d055f0e2d56dd7f1938b80581f1ffd233abc20e7c8044653207d8bd1e5306f2fea30c0c14e7bcf866986838c00d76ff1e9e0c47623472d7bbae64252cc36d7535a57700e3aa85a4c5af4289092ca46cd5993582bde14f1604fca75df49405c82a34400c6da20a92491cd2c78ca9cd918692cee61d1e3c6b52c1ea37703a0ade5bbec3ecfda338f4edee58609b46fdec56611ed256eabb572e71e9d775a25f1a8b6961ca390b21009e0a60482b669428f0c24389c94410303310b1a1624f1d0d1eb00eb033f0388db7c1e78f246a6a54cd83d55bdf22ea2d4d5471dbf7b2501f9f94a3ab9824bb053da613c26a98c0d579328371f0eba1ae17168bbea9b06069c3a37eb169e65f8ab32e3ae254eba1b4cdb7dbc4e8491c7154614aa61cca4e68e233b52d76930c4eb23d08b7fd8b42480a8b469fc258380b0a3072a1a43b5ba0d1e79b1382ad510513d093539656e44abac264079d08ccc403b0ed78fd6f5f1b806de8527477a44e354d385d845f83feb6a101cb6be8c6a64bd63f8025644c3dd8973753f9287767bf2436a0c1d1fbf6db2d96c9e10c75db062a3ac579896d6d3c1a1f467fc71633d1bbe8b6a668e23f79e1ecb371fc7f51cf5b9564b1ba88750eba8317f264c59be6396150bcf9e58014ff48c4c12ddee733bb78fb7947b8777ed01964cfd248d13e2d1d3f3dcd63be407eba8ba9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6e357d5cce6950211f428ae1b5381e36867b6a09fe01d4880ca2107df3e666fd16139c1abc09403990d24d5572bb4443d0105361fed81fe8da8fd24a06df21720ac2c0656ac947ec7716675ff2a0a462a192417565b8b624d0263814afc8280d63b757f78a34f65739b9f4e7f2ec86de0ac90a2ee5dba7aaa4e3322461ad9eb6e59b50ce7fdbca120f8ff488fe1fba844532ac409b04e58cf982d77bac2b8b02227b43eef2eda7bc0259576a93835c822dbca1da8d2bd505b11effb342d3c259689a5adb46ad33d655a8f940316353103b660dbbf7ad5b4c2bf33cb319e9217633e33addcb7d729a6daef07253b354d131293e44fac8e5258f27e6bf4b35cebc450103a8a927c84424d652ea86f08660e0c007a3309d2db47c1a278be0d2cc8b62a607753e842bfe07b21e1667872a6a9228bb663385a56bd5284277318ba4bf5d68b7d720f5316b4d9e69a7cb2940cc0148f682a95462f2c6bafa60cf10ad0709f69c013f67e9000f1a00442581cf87b3e04a51a3919ac1d7b8026537486044a4d37e230dda401a0bfc631a390b8d0fdaf21db50a405d4396c49c5bae2b0995056dc938d0a690dcdb750becadfc67fcf757ec527295bf73e1cd9ba80c53c636033046f7a126f1a57377966a6d44908f83d22c72754a06fa992bbde34d0338e1df4b85110ab3454d6a7e2a6e8e579433d4968bda43b5014887ce97a08bec2aed3ff2b59529fc87995427acf9d7793c1347c3ea9e72cb744653fad7df210bd808aaba5f562a3f503df6ca8a8b2c068e6bd26fc6967b5f1f5b9a6ac4db0c38b607edc49a0404c9e601a75bce2f7744ddbd3bd887f8a46c1ead32d202a68e91989f53ce8eba191bcf4afda9cba532a62564867cb0f675b9c8d6509ab513491bb68962d5025e6103807f9a0571ca7175bb21e44f4947ba138e847903931539d5550c84fab9b0323ad1ac9c08950dc601893c203f2ad0d8c6fc6c91ae8c17be030d7d442449abb34a01e378ca8ec84861aa3099b3bea3b793749c6245dec073bc5141987d50b552a75ef1e18627755ac8de6017e07488b1ba4038361162c1a4e094e6e5d01d9d335dc81fcba4ec47bb9ace320716b4a2e1fdde97f2cda14c7a01d5cd7d1bf7517442a648df1519a399cf37c00a3a94e5c05e43f2180af72aca259dcded7e63bf2d2e232716b92f7472832e359b2d50c5705b208ef00c61af5f145e76ca2bea17d5ae31fef05e881037fc28216998d410008e016c69c9f45666bf8140e85dec12278ca9fe2e33551c2e2dc68c825e85f45fa302ad18f49d3def8e7c7f889321897cdf20a9643ca348a141410da664cb3a7ec5c37e6650cccbe9e1c831b098de15b1e473b43975898af43d496bae9e477659d54aabdee08b6297dc0bdc71a42d078d9f6734c4f342e5f028b5cf9e67e06a50e3a20e8b344c2dc173c452d500d84dfaa6ec26894302968c0fdf0c0a692653b25d8261fe46fd101f7b2ce2cbad17dfc067c916d517755678cc473387e30990e62a5da11dff12337f3ec2dd72b1e981d5d96eba5dd1d2b22ccc1db950be249cb25516c2dda1671b7ab387d25a329339edc4e4783902a6fe2f045a253b741cf47f9ee98e2a98a9b7c9a39622858bb99732998838db40a91acc4708ea3d08819b36404090c34a6d9d0f71ef911733c00c7d6824355b08b546cae6e0c308bb4bdc0f5f21400328795f769e6391335d2716f4d983dc1c70e1da8ac83dc2d5c5a08de138064af002a75bf0821b902615ad084c5ce9c47c0493cc05dcb0f4e64795483169a4fd83b752bb451dbb77b5c9e237be865a38fa71574436151847c38b519d295a8ce868280338386f821e028d38710e9e57f54d5561d620c3db1374659962f14d3ba112c111f45e9d52851ffd4840b073a86b42b6295a10d8106d89381aa9be41c91c365de92cd86c196002931a9dc9845adbe635eb2eebe25ff8ce493d6e1699e23a90af0e72e5be00453d040b282a9ae6fdc9c2f3eb992591aa518a9b77d30ab6bd57996f11932a3053b399f8141ab30456f193ae7ffdb0e5426f8856ef2c6abe28174dd81f82d0098609faf20c587a5fcc62603268abcbe229aae33f98b8f5790bc53d1504f1ec85b0cae6051c14ac6fc22bffd734979ea7315b41cb3d6a267439b6d89f2eb23c21fe02226bf8b84d642b340fbf14c0e8aa532d5d717a0b4b428d5ed88776ff7aa32e73b53369fbfd7452c7021e5d965746a8576bcb0adfd1ada67003c6024a484d31af70ac14cb893bf9799a5c9b7e245ed4e3aa9b500a34c3b8d81adb50cbd9992b97c45b8c754e4a7e117b5f3c3f772e431f7c2753ad468ba0f08c5ed2c5bf0e3c7f0b98b1903575df8bad35025801d959f3659ffed23b799d306614724d63a955f93e59f4b747cbbe187eef72c7b49a90b3a5c1a4651750389537a8695c3f24bc33876d67a455b56bfe0ef12110d0f7ed305460761cf1b683e4c9eb2ba1d5663a879defdc0231f775fd10b72da059cee4569bc60609a8ee483d1f75c483b22145054a34d30c5fd23e8de8745d30d92b32934d02c7e7fd64b4584efcf7ff5c767cb1f4115a3f5e22ce638251e96961a873f152a6d36b41217ca05f081dc631e45e5ca423ef4a55a647e6f16b5392ff9a7485d3885c500b78f6a3698d1c2a32cadc7c49fd5f0481466d5c940dce61db2249407180a774f9a12908698047975dc1586c918d39ec3e9844d4a8389e8db67c45be5cb95e9910e5c76ad228d38f5f07d15919d7e32b21e41c238acee6178026cf6011bca3cce4a5b1ffa27ac4176264ef0ef6c012d530eb1e681bbb3ef33854996ad160d61fe3b768dabf11aa3cc3d6ea8390615357d4654dfffc7d5da473be943439434e93e6eec475cdfe789ebde072b05ff9b9d280d39bea6b2573f07dd6cc917bf3b00121e4bd07edf2db97c9de4e748b9e039be52d1aba32f6f8a0f1cd9678f60140b6ed05e20fe65f0157985a632210e802922ecdbd96d9547bf669189cfe2844a03aebab32611c80bb6e3ae1367345e30cd40eda1a5c12f056ab6ac7826686369d86eac3394a3e3d8dba3ec43cb275d957cc0bf31c43d5b839048641ab285af0ca5603d9cbfa619814a148b1e4bd16c626472c7b08cc1000842e42e3ada156c019ed6615391ba11cd1668364d6f6d6f98ca774e901624ba62de7543471858853740c95d05002cbc4a015e86055668219a4f9762211a703eb667f1f47fc14192f4428f0e35acb885f6853458c0bce8629fd8d2c8639b3a6dee8936dc7871bc7884ac64fa52b474199abd78ff6ab56f231944afced8e083b1db2f17344944ee269a800b64a2bacaca4ff44e62043d827a878d47e44a8d60089959bf239a5bf138bf565da38201bb06e679c91d67ec0e02dcd82e013df6a33a023598b540c56f86a4d3427e5f3c879e9453bfeb6404ed1bb92a9af139b64199d310cba6b55c0c73b766360a2148744e5d369f75d562991c1766ba00085d384b5db60a49c6dc88033b553331b14ff1bd7976f539ef95dd021561ec347d95bb53e9c132097dee185c8aac2f741b966e0792dd7e0f4ec7724fdea8015e1d8efd19211ca1c534d661d54dcc900079a76d42282ea4b66f0b440458f54b2192570e44498c3868414b26d3052978b9cece614fbc9abf5fcc2d9cdda32fd89fe8ec9759a57c2f4388ad0f1e10c9ebec41bb4809905c4ef39f4317e24164778bbe4c0f43db8add7379448eb2749462d42313560357d28c93d4097a3a83672f34b803792fdb8b64582ccdc6653ddcac31a414739f70af78d019ff428d2969ac410d9b4b9ebca90e7088057baa258845db19b0d66cdaf3c8de2337b0ed21b303446edd9dcbbbd41017c49f4c4d9743f87072226c3d6545399b652413a19e61241113dbe30aab90f8a1d4d28ab118ce351be032c3e1e791fc73e3ccf21a28142728346c940bced2e131230c2989c23e7d69a483d2c08fc91e922018f1bd09217bf2f7413ab0f50f3729d8e181e97c16bd7825d717632c03f5948bab4a7da3a9917d10f52c94cd0ec23bb3a9894bce5df99c2d198786403215cdc7cd6a7811d2ae71f8edc2e9b67e2137e9c747e529c569d76d7bae017805beb03e889e8e966eb756fc9cce8c3b44b411a1bbcce7d734f14f49d8e2f8ba097d0e134b57407d95b21162c7186232a9b80181ae6322baefd0a29f6e7b8aaf95985fa666fcf73da24574e4e20dc2b5b622225318e7ac0066853c51704d19bafa513dbc2776e6bbc9e43389d38eed2cea72585a6b7d357791a1dde31c1e065dacb23bf64b5035aac74ce92a4aa8439edd9f13b029b253f3529834e46eace1f526ec7017f8d1037f000144988acf22361a2d808bdbc21dfbc41e1c19d24a834ca1f6e2d643c872471f791f21af06ddbb174993d16905f91063af432352e60fea90039830a1f8fd146347f50a52032df7477f807a5d1eec8e149420632288a036b1db9c3088847b467e2a9d2038d6a5ca74f61f2336d5ff2ef725ade4b0cb5a0bfc92919268ebc562b5832fe1310ecd4c7b7b659480d5acc5c1f0b5dbb10d6e12cf4f7c046547173a707351f869d2bd08de668065d5283636bdd493a6f9c39c0e1169362c4897de592a44454f926e0a05414f071697b45cff67f931bd74939159cdb10da91fa4a03b89d091167a4c0600d43c4e0d3bf60e89f58889e8e02d342ea91e1cb8bd18954ee4a41c5dbc64e1b192950bbd6782fd8ccafdbae5caba010ce0bf9f633735860af032c1100c04e572879dfdac9fcf29c211384f37a374039534f0e13d28aacc42bbc127333c4877ef4347d1c8fdc7b66c93f1a99e7107b6ba6b297cda95414a5a59a254e5fe95918ebb51eb2a58bd818f757f6dfe7d503d68d87c64080f59bb12d13a8123ef11c5e108b5a19c7f2cf52148221c4a66eb4b22dc9d996c7c762139a0d4f56cf9779c9fd3218327e91edacbf698faab4577e3f39472ab793a0a2e225e1473fdb4e4484d30fa249761d896956699df05fde2cb6e87e27ebac3ab41d7c212dbe7db6843d78c53b1b621d6aab413366e3f61e20d5dc3dfe2c98bfc9a5bd95029d6d7c5877083ba05629b85d5ac4300406977b9371dd874ebca9c480b920f02afa0cad8a462eb887754817d762685b9dd721723348ca5e8ed1eff5d4eb95e27c75e13a3ca7ab8c914b7cc8f46cedcc0636d8b93effbc660d50c5a45a73b35ab03b0565f0e56bd437a971151f1065bf384e9b6a547e6389ae7ce5de101f17c528fdd6b1a1abf1769a83af0127da7af53e97cbbad42e62b1d98dcfcc6ff34474f68ba12bf655ec10f8e2eaf6570d5c2b052651c78ccc1b4a45460fe58a85fbd3436cf62d3044c3723ba41c08c7e719e2e8aed9f3fc21e6cfb69a206a1c1ba87407a45571db94c3757166460db9cff89c847783ebe6b7d0936b58ff98132bc6d88202b6dfab5ef94f5f035452af51bb0842e3ed77779f67d60ab307562668f88e7a1514057df9d9a54f279e61ac4079d58d80b46b4844161f7778b7256d4f884bdc1b30cca0d41865653bf048078d2e563abf90d315e01d801821e0fe2b47cc11c72d4b5dd525922d9d639a0adff4a340cdb3c550d0fe6949bb67384882c9744a26a7c54970616eed68eabdf0e8ea3d98b220749afe407738d7cdb091a2145c65f3a10d2642b30bcf18abe3a5e93656bdb351bc2cee3825f649d397109a7d592ea7220c5ed240e39c625f148b8e9e6ac6da6eff28419897c1e4c46bed41f6b2e175dac4fa3223c6cebcfdd4812708280aa8be6fd53b6bf923fafbc3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha26900c483ae59b05d01dc5684f00f9b3e88077ac81d95204cac808c4ac8e09685552568598a2c1004d08f3fd57f2f9fbb4de860de97b4077f57e68b4a044dded499ca40c71eab9fa52ebcae21673f94cd011aa3eeceac912b63d2f428509c855725f44222f19fcec801b091c2d8e97cba65cef2aa6d865ceb2f7af87292e8a95ba76a95ebbb3504a51f80a808c089db37b57c2005ec1a9d9f50f129c85d0a3d874a19be08a0d7bff7cb205b62a55a9945d88d42cd97ef007044ba3b454cf3e28050847a7f06aaac20651449901e8e216c28edeed6c68c4c7986e13921acd9ac46c09af1931bcf5a3ee738f5cd39bc414a0c8938834f7fe530cee093ea69284da8688a759249b24f8219b70743e7acd5d1e6e483783cb65a0b386214be91f185ddfa2e05140f17c3b15181a09dac2c37603306c5e13d8a2d4f2f4b3d751ece09c0b382a2a1ab0d672eb89affe086b9ad44582298c8e7ca46ea3432b41d6bd6595424f734b6a95a8f504d86d4cc1fcf867d82cab60f997047913fb31eb654243583960ec4d3ac3471b2f20990799d873c84fdc3f9082c61abd676ee4d40c15818d31d4506c6db5365d8953f4f352c0605d8db1e9948bea39c8aec97f9987f6e2d3e7d9a6772e2a583607f4a7e958d1a8619cfdf20d667a169c26b2793b9656397f7ca098079a0bb65ce032dd80488199af6619c6d5c9be9b67f02ae6b622915fb74a28c00dd551feab6c78ea21632fd843b8e24d523ffa3c1746f2e48611bb3537d9b2953dc7f0a36f30a5d32fc2d186f32852d5179870ac804b3b49b9ce3df4901cccd5728ea14667be249a5090ee77c97723abacf933a964bc59f5f8e22927b0f1d288a6b1e4007c275ac628c1d54911dd885aaf05bd44f2d645b4d1bca2352bb7515a5ab6c1ecbe01e37797fdafbc5a4ae1e5a06819cd33b80349ffc5bca15dc2ce5ace4cfd44a78742164db6acea4ed984297ec169b1b82ba66c5d37659ed11ded6ff3d4e4758a2c057c9e1da0ced798566aba6777fa1f3ccb01683363076c1bfb6d3be61adc2e2383641409161c9dc1ad912176b7ef622e75e4046f93470bae60b8f8e3fbb4fdfd9f7217b41f9099f86b641b0859954340372c20912b81b025ad5718842f4f48f6250c44e96727c66d91d4917ee9fb618c2f6897ef14035e68d08395e5f7488b87c38a70f96c55c706db5d2149c4efabad53eb029f26cf7578be3ee7101f12732f9b516bccdf258806c3022d02d92754515d02534461ffdc487b8c28c31935675c7813224652d033b451b6b34f86fd3a97558680f47e7d8f0e20b154d2e79dda9e5c4a7117c87428e6af4a02041234270eaaf89a0879b9c74bb02b92a4c4e0e4434a6c942ad301577ff80a6a8f8a93487f7897f7113f52c9a1f1cafd46b03de481e87165183a4cc7dbaa49aa88524aec15f85d78c4f50f6e374a6569a7651a92e901adb9a65f975331b8fbf534469104f024b7e22d9f744219b550d001d808cfee03787fd368865f4f5093993de7aa556082c7fea5a2349a4dc08f4e2a44364c79ece4a9a8a63a0b6ae362ef4b61db2f8af3c1f79a4bdb932bd6cf5466190ad3844c887e0861c38a81e5472f730e086d7cbd51607e11ed6676d2dc2a75d63263c7f78fb90008240006a34a845dec984ecc516044c21258c71a8df11a6de472881e0c97717fdbeb0ed6a2eff0c62455d1c0be5c8ad223437d2b9aea0a552187b948391d4fd755c916ceff0a0e80cb7fa172ee4a3ed74e47b820abb9bc3e1d9ba8f51d77e9485b85b3ece8c7e92ab02ccc7f64a656fe32eca1539067c8acacd4bd528af078c8cd25aa7f5f233349c71c0a55758b58568a33d2935e442e4d70fdd694adebd4545abd24f5ceec2d709510838cf9d0df2f9742afc7c6162b0e3feeacf86da36be7e8113194ae38834cf20caca0f0aa068d0d1703479e4e71bba3dc889e800fcf8ab8e302da8bd7a75b416cb3e4ec5f13be0f1a6b301883d97440d6ac8d68411231b3b9568aaca13d90e6ee122763b15daff78233aec5c519be13e36551545c747dcdea6c32ffe607eb671e46fa20c9eb7ec342654ae8746f911fdf88a10673277e9dc7982a58e7591bf2162216bef058bd29c5091bb7dda6cb0d6d950c2b1c11960c674dfcf714aafa1c9d50825e79388e4a062b67973d42af602dd8ca8905cf11b89a68776b0329d0f44d217ecbc42beff2bd5091f97c75f479d1e28c610c99c88a8833b024db3ebb044d467265d7939076d70bb775fcb01d3a2d31a94ddce195f7a4a0651f300e63e06de52ee2bbef38ed082f51fc660cdd1819b83c502f965e1a5734060bfc85b1f5911871706aa7d6ccb6ba61dcdf5980942fde05032b0b262af371e12cf85ae92b2278b9814622c536c025fdaa1d9bf4b8bca847ff04d36c7665454915dec895ca012cd294a0a017df45de48df659f70314581b903703d3c6e67bc1b64e043e5378988f42a629675f70106d0f262faf9e56653e2317dea4ec7b05ee7eecd3fbb6118beb804541a4e62d647d32ee7e0ad245a9b0d9f360add7fa08880e745c68bd78b760055a7134d6d292960b05fe6dad8fb1185808eaade4e7f05989436c8dfd8d81bf84dd8725448615de252a33332d1455ddbb8775b5628ad1058e5634decf5cf21a389bbcbf5bc3efb575ccb9894b8ba09cdc29f017517691c334ab5ec93a538c11dbbf01acce6868075223ade2cfde92a7ca3b258cc524e7c6d0c761f659b340ccffe0e15ce1aa33e45147730e381c47d1e5152eb202aef0f2ebd676139848def3781ef451ed9a5d306bdfd4a370df78f58695e52758acce11bf8d41197d1f49ec45f935126999110e31641219f39061a476026898e2c5456d4d6cbbf920dae9d92e0c64b39c631158e6a2e6667b218d1ec0f400ecf9adbb748daa660aff79eab198e24a73c7210c83cc4c95cbb84542b67b77852458b414f22a8a7ae02a6884ca33bb360c5f9c69596170422b4470df1dcb94a0e9548d453877bee0800f136f44f693a9483eaa01fe89852ae19cd55d736ebc6c30dc7813f4459a35f5bdf6f216c134986dc54ac7e5572129c07561f960f04d12b2be7aa43c765ebb4737eb8d39b01878e87c5600d2916e8aaeed3b1795024f742f9f500cbd81b5839971e9093df195485f00d63df08fa3c716733dae57e26b4e5415324437a07cd3e595b0a8251788443adde850bbfcc52b143ad69abb1504f4256a35f66b5da55e006b67becc81f0ac5631eb10970a2da9bd62cc252276644bc5b0c3d15912d78713d0672617204334b4745a288b0adee92e65c60cfe0f0bb5e08ba79ef939650ed4bd8d8b018382148d53162e625c1ff984a855486d8559dace73464d891bfaf09de1d351a92aeb9d0b26f92a9cf3fb8099d3bcbbd6ce92459ef72c4cee47b62735352506f0f243ed036725b13b556b5d5c5dac1e008543b958334541bc3915c69e782d5a10264536d6420a06a6c10b3418fae094addace9af89e5236f71742d0ee56bd3730acb3f02e1c538e7c95c475ff0d1735835c0b72ca9cd916c7e11bec7da55c0b34e7adde03f04daf23f99a6e226cf8bba96ee82f24098a8c86cda8583e26549db9dfe4c0f4715a2d22e1e428ae666d47185c901b5beb9ceccf2e00cc30de5af4ae8cac22f09e3de872e0c7b448a473062fd3faf2bfece175810e0c5a3044e11f1194df92c9a5e5c896704ca9dcbdb5f2f7554a7f63a4dc84c536b557aa2b9775928ad58876bd43277409cda5cca4cfdf7801c3087e781c5baee172759a17feca1b1b47ed9d998dbe55cec3b0b54c1fcd5fa6365f155c9f3f5c35874304d1777c4b04ede2c44254b3c3c372229b9df06a325eb841bee8548385ea5c244e34ed3c43da6911bb1a8998661ed5cb0f2f8c3c0e6edb3b97f5938012f19bf331bfb277ec887fff33881b9917b989b65f2092b9c19a12d87030ade16d242310d506bf72af005eb46cdffb3259df19da5f87e5a287d763af12217559195fc1881f153eb22e9c69747fa42267ed5059169b796e9c5cbce30e47f330b504a2f30ee6c660e1da821b6982caa5907544986bbf02d7d7366be7ec869ac165c60e62cec28cb1c0f79167eba9f3fe794319ed4a7deb07a8866002ea1d5d1f32a4ff3ca399dd1ac506f440e517d1600f6133a31c7faf1b49fe02f20c141bd1ba36847eb37518ee99c862a40997cb45a352ccab8909c3b09f02837f952f889d35a10f160bc28d12830ee8c703652ac52eb92a3ed4c09495d5aa2e5e98082f02cdef57187d7d4732f97b18997a4f58e28ccf9356e0310749a1992c546f7d7ec684b107e14828be6db893a67f74cedc09f98918a0d4435d87e5ddca5333f073bd9865f519638a34793b0e714a8bcd4b04113c7ace6d828e1fa6b0da633d0f1d625bf7f3c25b19d3a50e553489735685909159df2689566fc4d7a98178e6644ce425b4ee4fdd16afd44a0b76c5b990f9ffa097a173fc4348535083f393e17a6eeb9ab7cf8762edeb3a63c06f87adbc4000a8c4763cb18557ea97257684e0043a604b499cb0424c00651411b33198711e5a29b038fd9b15d21e46d04a1b97502b23d0f950397a68be7ca2e3df6fb1bf0618e09ddac7f4f7d6dfdc98883e0a9b6a1a24fa0701a761381668dbd10afd515d6ad22e087cc9f02664a834f2250e51a58c121ce77d4488a4527844e8a7e6e1b7eecca984628dc12e43a205e8c77b2dcce2fd68c2c6522660d196905a802de8f9405ac6e78d7dc6c5d6ac4002fc87f910760dcf66d5c0d8e0a050418252078dfe08c24ddb5e7caff8ee5b034dc514585c78bf463685afa0fced730568c622c23d67c7d881b2036820bac9aea9514f6f12d1b920f08decc4d4ad7c3f8dc9bcb5dd47ca862daf0c2873b2976a03e91987cfc020753432101168763bdf25d316fa0045db4e099a2c1fbfbdc8a78906c693e09d343d2fc7b477a09b2b5b38e62b2a0882aa356a0c0a2eac7eea20c541c7ea25577e8a9fe479c3b24d027ced83f0f3b919d8044e161c33c164ed017c4bc9f5a4083e0c238030a4de0f1740a0ca8daac37806d672d0c8173df3b9e9c916bfcf2256c7b2ca23313e218e5b3f353f87b28aea7ec256e73ced3acc20cef15ec304b6612b570cd768de44966cf69e1d09d945eb69db621e22e1d41096e50c819b87339bc0b6763625ddd1f8d4fbb99f42574810a1788026edf5254f4b25db7e8f42b55e1b4ab889103fcffefa4cbc40e77f173c6bd4ee878ccfa6c74b582b8cba7095c99d50ae8bc9ea327028a067a5288505463bceb9aef0066ecc74871848f054894a55fe925911809d6f4d174addea10861753b464e9b4c9c27beb04d1266f84007c30cb55555415bfec654dd073405d319c057917cdd2a678846bf42d2cf7d8c0a761d673e9c05f5549cd7af7336b6549b0b88f9c6ea7d658efa23b8d3b6ba045f478f7af18309e89c3cce87b09f453a36fc347b250203150a4103b91185a32d9763cc1b07ef6ef51917847d6ddf65c36fb0cbe8185504b0b4baf522bb7c79d95617d80a1603aed8f5e599e691bdd1c89cf0f0eee0e262e949afac7dd692f06eec40a7c266ec65c93a29e02d0d4785a8361d8774a2147bfea34d714c65599492b6027a0bec9df2fe303cb01cd03c46aef1c2249db32620b02c0a7457a74b739e098da8dca7e0b3fd1c240b041ec96b3e5d6e472e2d1e8f093fdc154d1a78aead19f46b1ab5c534f4d5d67e28e1a3dfc14beb58b7c707832dc0d10ef9142031b85298789d46337bc20b50539b60f45dda242b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3b55bdb8517da6ab3fc37c4b2e54f29ebf8d3af2dee506c962bbd350fae333f4073227899c3db849fa30ee1c1357728e2544f645dd227564ab6a13a8d978172a67ee3328b1027f12e7f60fd11f2ce10502599340cd3888347239655c9a5e5a1c55b838751450ea09da43e93077e377db52027ea80ee0361d57e9b1cb1db53bcce1cbb9bc29e79d661772c09fcf060cc624fa01e84e1cb64c7e4b567d46e016dc56bd5b4e9d0e5141414433406aef8ba719250bd346348f9039333436540741a517b832f3dbaa64c0187a324ce31c0b2726172f103cda8b26c50f50bd1b0bd31fd331a51d14bd5ac2576141335ba3d799f6277462d1446f35ee9f9edfcd70f95718422602c9282162efc84fc1db0de1f9e03779fbc9770af3910762f867917adabc970ae3bf4e6bd883233ab0bd1f490360a211b0d17750bc71274adf0a0f77c07a8663acb5dc0aefe3ad77d53d029f99074d8be7fbee00be8a95836e43b25148024764cd389c9ef9c769356ca0c7641351ef5c2b39798e390b537982091bc47dce76245b7d085409c635dd7acdb33612384f7c7a821ec0b58444f002119c93b8b351e6f5072bb943f6f4560c325f687c52dc96b9a14d47575c1a263d466083aec6510356991840f7ef8c69768f827c39f2f1373a3d4cefb4f5fb7627409f9973a807afb7a66b9fb72d683b228483642ffc0ebe24fb6dac2d26903de9ea452419045bdc53d6b1ad159887e6d78c99ad496d6356c64f29891146bd692e2e0dbce81c70562be15a3d5050cc9df76e5eceb03f0fb9388151b05e668b1f7c44cab485c73baa170ff57e8546bd8178b7f67e0a4a62cd8953b1570226fd8220dfec34af4083acd817b9ee7339a6535f574a4050f239e46d67b21a43a3be04a475e7bed43de278266adc8a040b74ff6e84d5e9cb1cf4604d1a37ba3e2baeaf154e764ee58887cd1a57eb7a5649ac2b99d294d015439fa2529dcebded650317d77b4634ab9addf0c99c3687f5eaabafe2d9bffd1070c054c4c7ac70b236be4df121dd5d48b720efe5e1347b7dc2af293af2d42153281762342fa522c393c04e03f762c7ece42096f5fe7cff6a10bf51c34b10ec19e6d447462d0b13f6308c8c36e36a096f9068435ddcb3c1fd79c7f901df2130400731f1d38bea994f74371b60413fc263ea2c06a872a544575aeceed4dfae178cc37e13315bfaedb67bb3ac61206ac860784d4d7a52e0ab87eee9b12667b8472d30b98aab59c918890d91dc0c6aa0e381439ed7b8f1b8368bfd58219d6e0f2fc7998dae42c12e2c10dfedcb10d837f7d972ee6c8b0dbdd7507e547cd29e16e996bc38f597a460fcc7507bc6237fe3f468375b0466816905a0437a5e552e8bef232bfb3eb3fc137864b335bc207f8082fea801087dfb6161a631ae94df8a0704a6f15c178a47da5faadba4747b9d9d343ce009107ec3a060a6f47690e08c5b10589c174a753421ad5c54b3171ed628814f8139f0678b9cba58d59f503e713b409a08691febb73e3f6c7f18a13a9a1e6e0a0c05c7d53041d5fa5d6c59529c7a57db827463e8ba784d1ff668191e604c550e2041402c06c9c6cf3b2f243a2426e8caa6bf65b2a0b88696b067b7e4edb73c09c9ac5500ba4e7f899d2d0190cd1d0ada7c4edfecb98ee0142cb9d2e286c94c6508d3ff8cf0dad9930b412c716c096fe2cc761c7263dfcd26783b59698bc047c67787e73ef0f6dcf69fe8097b2ed094dbb6c013da5a882096a17e7a15fb92d2b00affbb0956f170c7c2f69a6f766956a45ce19e3444e4680e3fa11c4c6f0a2699d64291fd616b94dfb5cbe9413a1c964c1e132f0073f30c2749eb5af61f5d97d17b3f1588c09352acc4f9ff6be9ebe73735369f6168fa5f396200badfd6947ddb568d7e44fe15e4c490e85aff3a6430c95918b0dbcbe7dd48c8c4d330f1ad7fa9e4d2367ddd397416028c6a95e51b3a62f7a426395bd985268ce32cbcdc1ba4f5199a7cf06dae6428b3f095b87eca727cbd01c8521bac0dd6df8fec10a438bbd053974b9c355b3b548d3e243ee019b7482305ff607431a95f03dbd87fc944c286cb2600571742085641ded9bcc03c512020036c0796e7b7ad01a6049440f67aa1316be00d70a6f1b8de9a02bd6f09d2705c47b39ef6bff58eeba435ddfdd1261363bca8877932e0b75cea7b5227a23819ad20359b3027e6cddb5f1c028cc746eed70c777ae83a165977305b3b2eb74eeb6e74db5cc02b7951352b3f66186d027c6c4ec50ac2558e8781d1029ec4d86fa24da307dab7dbb8d21854f55615d8020cdc90ee1dbd7160b1edf8c0bde82ecb8b921ebddcd1800b35ab639a851b276a4c7e8f2940a10bbeeb90c45ae7582060670013a4c2ad69ff184c0bd0059099cf120f1460d759bd506cfc3928e4d1b2ff9c6d3fe382bb4fc3dbcc720f6f67cf2228b1540824e992b9ee05a0f4cfedb8f84562db318ba844522b84cc597b39147b48bfdc22c50bdd87e27fae2930ad10d9c58fc0c3c409fda6e9ebc375a8a724916a8dacb8f2bc23c8ddf005c58a5ffa69fa24f37c354c700fd8c03561db9140328d140669a05a502eebb595268ddf5054a22e0e87b3997a8d576db83e8b099d6842ad84171f9649ff293daeb058241ceac296648d06ef4e522c716d1aefbd928c1a6ea1abf928de44b56cff57ddf7b84ed5d594b388488d63f4109bbd85e0c6858ab90f628922d57f939047dae113445f6a571476b268da7ed3ea0f01c167bd46aa619185b1191407b17adbe39b720d9b7c284ed7f5e80a0abcd9f81714dede28497a51df12afeec4b5b263f168dd52fa964360e3b4960898c097d943058855797996aaf4f0388118aac811cca2148af894b4ad1496bf308d3ba88ee45ca30c779148d3cc3600a8df762c43b70fcd86d1c82a537a218d2e278726c54fa81b5fad66e87cd276b2933e5989dd98cbfabb930ca216ee4967a24a34ed68e47b1c33430a8d7a4d34c573cbeb2188f5a838dc7454d3f5b14871536ee46ffd357dc55df877fb4367bc7a20f133b3351c30373d8e684f82b78ac7b1a8f5bad8f58628ff86392a2a76ca27238a962caba00bea5755cf8695a48e2b2b82cd88736ef8c56ac2cf7ebbcfdba8ea094403a4748df72fbd313b38ce41b22bf9c3aef48d20d3244cba926e7f2ad950a9a2d5280903fd109568ffb0b4a58cd05fb7e6586d71a2789b14c4b6a1d9b8db89031fb2cda3cdb0d5110abc6996cf40b8fac6f29520a61c7a2dd1cb1bb3b5f5b6fb4aeda4537e1bc7e7bd823b3fbac6310460cc415419886847e81b1e68f4f650354f7267b7443649cdafe63d7e7b71ea34b7143255566e2748c36e1d56de918fb06160bfb99602c118c1254e48dfa5b88b1c7e7219666e63dc41c8dcedef8e0bd7709bd2da5c156ed1876e50496d5d3447f1465ad8c677af8e784731dc33d8c5a7c28afd5f69ad93b845ec3127aaddf8867a4f013c664635396c655b9e23907d2b22b309a99de84e8387c2d764ebd58965a3bbeb8ac29af4662df74c451619595508918a767d06945951e1b56a6e3f069f439447723bccef4c46d0c18b7dcdbd7f293f208362fdd2253bfe01c7ab0e9b5299fe8200303aa1387f184a79aa01e38aa263044c3c5db9151e06d59c5088f1fb9ebc374396620be0260d4082e82fe1f371991f174dcc1295c04a5221f8ce4edee83c23250b11e745141f1ad92650503b4cced8d83a53e5b2688b70f57cefed1a6b4267aab38cb9082acbcd479f86f685e08a87636447632c29aef6785232203e25fd76367dcc48c3ec85a18cdd35a8f8361b205d697d26dd1698d66ca87b64997a31c8d4f01ccea2bce39b4a33412b768dc41ee8920dd10f4c9d832a9332cd1b632872f838c755bd5de880c7be5a780d8c2ecc66a5ffb3af8ee8d804ecd7658cf48dde8f1e89e47ceaf7ef664931a41ee7aad8ac93be5732781c7be972ecca937b7b08c88fdf85b255cdb70548c389b6bd2bb96c5e8abb62c2a54cce5e6a4de921ebac174b2a2e0eba5fac2014499c03456d4f44a3872a65540c57964f20ccfcf9ec32ea2c1d9c1d643ff682fba5ee30e70133b6878b0ebd1f5443ad3de610dd58734c1b2fcb2eb8452d0612756af236edeb06938cd1c7554e1679c26e21b57c0200c975387c85ba2a4da2cbdf540e8ef652fbb604f8d13758b000633db3fdfcace2ec6ef77fa2fbaa6708638c5fccc69ff9da7a95cdb349cc68e0c99f62bb457c53988ccf6a3a5e6a9acef02a2eb58ff0836c0b07049c525ccc5d64eefdc62b5c596d22a7fc0f9f1aaaa376534c7cfdbbb7fc234739d604719fc94fcc391e2ca8408a6954ca71cd2485a34d81d105e155aab1ff21360944631d7eb5248ccfbedf46904f6c6ebb0e9e5dc821ecf58213809e27caf5813ee91758424be1092d22598fc8e99f0a811d851a3e952497b7d8d65c39538a4f6fde26ba9ca987f51b2ee352044b003ace669870f2540cf2cb6e32273930e624e5bf4261f9857a1d7e8d9499c794feb2a76bbde66efe30ac64f3944d0e78878d57ecacce18611fef480fd373912482e06e63b33c100ae98dd47933220f2c2c74b2f4366b189adbed94cea00bc347a7b46bda38df16421ef3aee0f2ebfe9c5a0d7e8cb41c784bd865a8b4dcfbc312a4f420c1e9103e7ca11c4436301800710b4a36c8078e9df93d9d67a925232e4d1f11f155b5e9eeef0fd1d25ec1ed48364da5be3dd5c0c09796b4d29da37de49dc530f98f4d3d45cb65b52c6aa0cf731617eb38243c8d47e7ffc87788f1189f026927b37e7ffe0827a9cea5ec97527cf0c8749477d33e2f3be47f2037df499b2bc4d93628b3f817e0ef13e1d904d847481c77dee4b98ebf324391e0fb3aebe7efe5c87f8b67388117f4bb60d5733d6924f6f2c348f576012ce35d6f88fbb3651407d7826acf8ef0d6165257c045cacd6992336ac113a8934709c6d9981c0ff7d4dadff1abddd4e88633f2e55e44536a9e850397393563144975fbbbe11c1d1fc4b12e51e72fcb3b53e71b921b2dac4a176b47f65de70f3e0856be044aaf73f826a01b4b398020f704619056e125f77402c369fa7a4a0b2cb50fec6de766e2265c3badef7e14bd38af083d1003758f9908f10fb24f885f1a70c4edfa6a50b0fa48e9b4907b84632ad468a4cd8629d475fc680c869f2a8e5c1e583252fcebe37f2e7779c4784b93de252ed96bdea7633fdbeb8166a0c7421eb50eb5a80d0a9dcb5f7ffba686ee7c8be2205562643710640d59f6d17be649dcb0a6ae40db028790f32f838d50db8046501420291fa1ca617d6d917863900addec60bca0c81dee321db01e6a7a8ee29a653bc4a618980525dec333176fd1df1faa0e7026783332c59a1c4a4afa9fa5e0e7f35f717d554e32f3099b0d590cc9ef4d4a1840d4d8de6d595112bfc11e46af003b7248d1912da136a7e1f34441062f4a457aad36d5e32fe3fc12be7fc44de34397529cff2c0c9f608499a8404ad1fb96657b33dbca16e3b345f1279208d3af9eb62e727a080321412526cbb5273fe7fbe4ee4c5fdcc6a8488c2d76eb382d2d937363e2ea7ab28603ca36a9fbb406a7aeb278f4a4cde9cc8427e8c4641a9b81bbb73e899d421c91549d8e5be33633d889665f5a97cf187815e57b11581a47bd971fe7dbfc7e35fa7a48fb9c947d6e5b11f48a33fb260a59a5aa6b017ecadccfea3fc7aa4399e02045c922ad3f577782da4394b45033657cffb74f58c1e273ce1a4d8a79bf95f868a817488c5118899af7c3ce960de9caf08af0e374a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcf100176ab13e881470b9e7547dc70315f326e1bda2b21105645356ea7aa9dcd831d32e071337898f17b46d2667f5a5408ba819f5faebaef005070c12f51d885698e8c9352d4e4c800cdecd753b2e93c8344cc9a2cdc98eb73297d3c1143cf3b6ab4370f19998631aab164ccc7dff8da438d93882ad9b21c2ab966abbe4bbd92bcb3176b7e52b00043bac78150cffa47a01103698910f34f3f6bd75ca736f3f75042520f099f275ebb21fa5d59b7f6f9f8f3701c6a5dd32af1e253c2b0d6a9c930828f26c3909eb8c478732dd2b20e26f9bc2afaa418b555746ee7dd070006e6f57b0dd8929ff659831d8c6f87138b5f34e6574eff9c997c2821374cc72e6ec43a360971e03427817819f43d53bd0764199b5b42a9452153b2bf0d8c202e296f538d3a1ebdd420304806c7d8d63af048cbf2907f5852693d4049816d23ad5ddd16eebfad0334f29c1348c7847b0327bf3616c32b1041993e046acf7b81729566a5f7520a2e3ed74ab216e6df3ad1fae33fc7dc4e6867c714f51d6eb998b3958cc003b11c8c39a8109ca179b37def0398ee1e6c810d5c58dc6af5ed484c19f25c15e10532028e045d643de1bc6e6240e59bd196e781d0a1cb490ebae0bc02e3cb13bfe3b3da36bc87f72b36f93082627efa95c652b644af9b640d833e9d97e55e5a4eecf4492d1cb94dcc245c01e2e69174e12a1efd99d1ef1c5f14e7ac05fb32dcc1f4918436532c667b36771f871d015352bac6489956182f5eef39e63e7b33f58e751883ae17e87b0ca70e778e5f775d54a1baaa1c15140dd468413176d1116e4f1f432bea4383107c66898fbd613b3c0e64f57e852f33bb31362995f2a2c7c880e5a4d8ca4219f9c383cb16763ca67ea904ea7ad22cf63ebc7cab34e64c514c7996d2e7a548e76069e556b5a749195acc8c998096c267ff6b21605e1d30a86c3a11857a3a37f6a37ae82a837bba7fb94e9ad68730303fc2d95ecd44f2b96aa9851d518ea7f67de67df1c175526b39f9d281d8570464e742c8797cc5bac5a7addbb6bf0877d6c20a3e12917d441b5ec9809eb6f267d87d6158e12adc85013c8dc9bad3802e117cf97a0dad23c64601293d22a50921d01d4981bfd6e123ea61732ee41c332c1d781befad4da445ec0baec1097326758603eced7b95e15a9c11f790bfde6336cc8c04eb29a1a0dd84a9020d369c53987dcc780e983ce0f1415605a2b9dfa0e0c591da5701308c914485364df822ab1b4ffb6f3c03ea8424798396584214acd0a108d5d8a35085dfaf3a2d588db9428a5defea92535eea871bc18cb90c0c959ab6ac2e6288553051b295fe7c0638e504b353f77bea488011a01f909e2140fe2e617a57de54704632604fa4012e8bddbebb7bc534d2dbb3ed55e32dd211b07c5c0039f0c97297e4edc414cd2ff573f083cbf4382b4c5e99e18e91fc97df7234e02cc3bf2cc47ec1fd02871e380915c338ddce044a35c8a4ce707afc69385c09ffb6219f84c7034e93703717c0032f375a78f65213e395172ea3fed539e986827df75ca3b67c20abed8929b0b7bdcdb87513516b633e3833871f85657124f9e0e4fceaadf3c3c91de1d74262906bbf48a77ff63534da6628d31cf60be5239fc8977ecd2a55f12179dc22e6766d20489ec13e34b7c49444a29d53930104295492f2d1ef7d4dbc4762678f542fd400a79cd8379794d2c254786c6a807251253a618e7e37ba7dd1096bf301c6b16ab0364683112d4e16aaa059b1528f9eec2cba7e8d497bbbdca44c4f0037dc6c56a209f903fb5261a7a5654bc6aa86bce207bfc656cf8a89c0b0e0ec9827c6a09c46945bdfeefdc35088701cfcbe83aafdc5fe14cfa5f6f5f7ed2f6ebdcb36dd74b601bacf1319730fe4037fd4338ce3e2f8197c7819500d292fc987b0f9ec918772b8026b611ff2c2844977fa2b568058fc5b738f31875a654d9fa4eb971bff360a7de2cde1f9aafebda68ea77d41ac61c84ec3564626fd38fcf8a84f5decbd7479d995346024812fc220c5720172ae9d3cd46d606e7d75d75d9e7c3e9391792f946e49b32371d16ad153439424b5b3964b6ec2f3b5ad3f8b047140f388c68165dcd088ff67670b397548361be23694caf0e6432cf6f5f2ee5f54eeaf3d86f93a83a4820001f8fc9ed9ae71f38c291913b8bfc58ae0d2b3b8c9d202e580b0b82c1651de16e4e9729bd3c185cc5d245df06bd71c02e42a1ba9d1da4cd1abe9af4f0dd0f1825116b499e983398dda191dbeb7d7075611833b9c79fa05ee0347b9c2967b6ad79adef02b1fa4d08fb7fa04c2349a9e2143e8894fa93079bfa228dd5cd330b6f2bf3c235b033d6d0a4d597b59c4dbac77b95f526453126602a5b4bc2d235d5fbee71eeb6c45d8a1e7706d03d01d99ee7aaef2dc7224ad65be1c825d666b3f23c789f679ae69e8a034d218e95600c4d1041203be749f4a4f1610bb99dbf78ed19cef69fc0aa94b723553b1f3c580ec695d2dd40fdf836fcbf9798f26ef8ec820ccf49f57a39148edd507eff77a17c891c4c386afbe6d428d5cce659b88e7e819c69002d249d3f785839a528d0b939f4173d989067bb57dc7ef60f39777dd7a21eede74f296aab406741b53c98be07f826d67b8774267e33e5b3a63ce0d67bb9e241bba4084ea623965898b911a3febb2455e80e818497aa041bc07ea687725851ae61e27f6b5870ba927a63fcdea7949d98a0084937690953a2c80336a66db8b7dec41ac5cd68eaad198299c24b83d6ccee6bc1ead2c9cd7b58cb9a7112675680256cba828c600b1445eadc866ded43020d61b6abafe2c27895584380ea1c5fd482abb098a90a5678c1b0013175a58d3b9f2fc2e4027d2c0bbb1723485311218f593e68c32d1ae8f5d3808a30bcee91874e8c0f60a4043ddc183936d589e4223b4928cbd8c40313328a3d05be968511e0d035f8f0a73441926d2940550e29d91d839a02278c29732bb61d1b678b45b78a4682c0015412b442eb0e30c0380ea8bfde7d678a6c98f8ad31bf8a7a47e5fceb9eda2738e24f2993525aa94d9d748b042d7b0dc88169137de4b0d2e1a222dce9e7179e1f2b1bd80f95a2a6fd04c8cb3473c3239b6c9f854f115660c1404a12a6fab0a66756d9a53d5691b6190872ea1a0c313ff036278a5aba45326fc1aa006a01824d0eb876f5e62fd760a1106b023cae1b2193e653b929a9fff34a54de15606eeab4713dfc3c6292c11990624a1f40655bdc371a63e8334165ffc58822d4d4678e74ab3e315e998d686971b76ffc64a701c43b820f2186f78763a2b87bfd867e5150c5e72f500997f0055bb31174c7c6a67281e16dae8f1230716a3547f64a5cf43e5184d84a14b9b906862dc522f383e035b13328dade695022c05d82f4b9d1039b69f4a9d069d572e783245663c3d0b717b6de077053e377b7b87201922e49253c48fdc8a15e5f6f016f0d39d56a1e62777bd6a0b39c2645754bff4feb156b0765ab1eafccb6a4a825ffd871943343ddbdc06473b0fd26219c43b7149e1ba2408dad01e4df1a8be0471efb618520fc368e84ddc552748918d6c085265766605b6f666afb1db589b03dbd3853274d8617ea55dde7a9adf5bd13b9d138a59c62710140a7b0f1b229cfc885128a565755f7f825fe18a2dc8c07b6cf67c62c015f36d1d828b00ddaae26e3ea7a4405af87742bb2eeca17b52302ba96be3c5f4aaa2f4f1f240b29c9ee3eeb96b4b41a54028e0af1886f77e8adc3bd8cc937e191774ae237b45c7341b4c2c0abbbad69624cf68dca647d97959eced1d81a30ba8474cfc4ff8452a97b25b0ec0f181d0f5e0d052f351f0733bee141165ef3bb1dee746d635dd250433fea414636b6ea197e70db2581d64f05b288991ce0cac3d5ce8a857c6cd5fcf58684abb1a20d1275f38ac3d39c77a10f5a57f88c7d6aadba7e5db88eeb2dce0d92582f8fcd0b13abd356a1b7d26899b5fe01e320c04667ba119f4f0ce3569b83c24b101438197bec65339e667e867f80f74568a0c7891acbdd51af67d2256fe2d2e145a5521745ce38461b1ab313b3e06d8a1dc7eb3fdf608495e303189876d28180ee09ddee7f06670877d674710d261dc89437654d743d72d26783d77712770514ec0e53ae1734a5526ce613b905fb3c1695b2bb5e0ca0da26404b5e0c025da4571ae97be5ae0575ac1f65b799d2559abbf74725428111b10589c02481372370577cfac7a6b21d4431f8415aa23e1fc770da1d8c73de9871917d50258991298be41c5b023200011040fc447e7a544b312a79cc1c20bae066fc03bc99607cdb65f13680558a966dffb4ab4a1c6bddcec3329d9a08cd0d053cbf2fc9e897c94ba3d6482f8a9b6a64276d5b9e01da0af53c39e23edd68ae443b609f9a8d727517a259922c20b10f010aa92518a893a8b310b255a3ae5af83f7da41b6659bdc48f4f908c4a8457e4291502c6754d76e0b71f52a504270f56a48c7cbb4fbd0827da93890b0daa3bf3e7ab64bf72fe01dfcc9ae50f26ed7f8187f335d3430938730a3a9c21361237a43753fcf00c98067b54fe6da64d17aedaf1c60fb377d2ae082fda983f0a8c43e62ba70c261451703fbfcd5068d27f2d2bee09bbca3aaf63adaca3d4ae190ab825a1998ad533bff154e300bccf7703096a67e071871aadc35964fe970d76c1a990b98ea03636858a3b7dffa1665d80204f39f0fd1e9a94c0cfd35925ca314ca7fcefbcbe58a27d86b80c672770346301eb9b2fb332d74855aa2f2ef056cd40800d508972f81a2f2b7f2d6099063c305f73fd65b87aead50d104c45e13ad68c012823d6de484eec870a78721940e648145e9e0b932384c09b1b010acabf98b677a557c1a6c7f737ca39c81b8d3cbed3d04ce47c05a984f2d84cb5605ccb2a7265c29d686763dbcea5b733f1622f1b8a89a08c63b5bf56d512bed296dbc32a12535677600e8d74e4d34a872e7d60aeabd34c922af8a6f142019d9fd42264f2aafbd51b96e0ee2e61fc4e966df77126c3307d22f129904e2bf3e1c32592442e6020049ca506a90de0de27fae6f8046211679ce31bcae27312eff61f612fb91dc64a1bbb8607aef094f3d8dd7da561755f3043ddb66a684627da6bc90ea35b23559eabea5e2a815dbb700f892cd0eb9202400631ac5f7089162c05fbdb0206cc1ba55b1acccdb73990cc3a6c4da61347c0ea837a3aaf47d738d04f97d8119a851f605272ecaab6be34662bbf65a2c88b7863f8e5659387a6f0479ea764777d1b6335b68ceb6547e2e1800624357808b93dfcfbb68c26387ae3d68c26a8064fe293c89af2a152721231ad9aac813e7b0baef9ff4316a982e707a3866ebc5ed30d91a00090919e23fdb2ef52fc1df3e2958a30125f1f5803ceb5ee207ba9db47e377502a4ee33b19567270f1034fed2216c9c65d37f01d7c7257d0fb7e75f62568120abd2444ac5355f6dcd04cef162911a66d9912ef8d64bc0c622b77b163a81f23966fef22c8dc6608d97814df4be90c647d397d64e6af07b8f91b7c59a093555d0b65e41729113dea31f239ef82614e21da12ce7133a70d9d3d5f23c4450bf75b975681fdbe1a20aad729cd2c436303f0b31e69d5c016aa8c00345b1f3388b58a348c49d7095ec6af0e2bb6394a44c64be50159642fbb237829e7031a0a2c782fdfcaccb122902927744f7b80da57584603f3ad2f42a5a5afef3f755a72b808efe7fc5926da18170299f0486a25bcff025708221bebdb1296df814af704e0006c6ea521662940d5cfa8e2b2d4ebc7e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h36ea29c2ae9519920fe67b14399625e286ce8780758bc88563f8def03c25d2c3c0953dd11756029fa041993ae97e0e6c54df8f985e3028f9937dbff3b58cb71b5e0e3591a22f91f1642bf4f5e8c5e0974309258f57fbfc460a4c13cfe9c5895527f190e8da9dde6d112f3b56390652938b5d535d60128ba89eca46a4ef338c7ae03e7a0476197df207f29fdc08c37481958f5d239def3ed746362b3dbaa980d80b646adc24cff7b8d6fec3e8249abf58646685258f8a4277a3cc41e4319c84746fb67a1200579ca652e18dc968984ce3e24901d6fc9f8fc93644028506d46c33148f3adcb789fa2dbce2a04692d293484938dd5e32d0a81479541acc00c5560f1f2c2a669ccab584921255d1c31dcf2ea14d72651f5ee55becdea0f90bf3f764d85a67ef486917c192863d954eb5539b439ded2c5706fc8b29c6640a81a6851313f6b44b5428eede233aa3d4679f3c0175765527d9ea68c5e4fd4c11b039a83242ca2f30bea112859b8d22db22c3740e3ea019f4926b90427d92609936eec0edfe1fa0d36765d4572c8534136eff7d6a382ff611c545d9d1e5fba0cdd95beab823473afb229b76993bd2fec203bab37e20b0c965da9ad08eae2592864b618d85e277d060fe1d336c19d398173e6474d4cd3492634cffde5d4b3d4a2fe6f10e9fb9beb5fa89ebd6d632db949945b097688b8e09b6ff91cd64c05568d734784d72986c64b1fe358cd58ef4f754b8f5e98cdf76d0b355edca97481f97c724e15bc6f36927b24136d86c55397c2b057220f9cb37f345b74abd5eaf12eab56af7a704265950c7a4eb6ce682a8eab0fb96dba75a1880b63d7b4e932f45c287722c68ea27e976d78b992080201aea975342956b97da54e1b6f72601105647e9a51bdb022fc8b46906d1e5049a357cdbdee26e01345af94857f338113ef8904d1b21c2c920abde6785f45c0dcb6837786798dbf9e7ec7b061e6868cbb35eb31d14f75ca193e8533fb9745feb1ad12fe6ecdbecf0def6569f2c31114cb383f0666a0aa07e9af7bdf87f611c3429bfe7a17af693a90309113e62524e189cca549c32da0596e95e6f5d5b3fe543facf84db166765930e3abb65c390b895e6a970e53f50d7d0ebd3446472fcdef3fc16d3bfe583a17072f532fdcd5d4d75e6018a02fe2fe07177acc3179f491db707d9a4fd76fd267a9ded538bf30a1851c2bf1373d44cca33d08f1736de36de22fb21f9695f2f2f2ff125f6a9e75b47f88eeb1187fc6c999e9698661c20a1a65f86533b105364b7a5e0104283036ee6353d10db35f8a6645dc5ebe8b3ed88029688c42221bad04edfe85c16b27bbcdfc35da066df0274709a09bc0901d53e257eddeb62501ed1d51784943b53a903552df9453628fcf7993841a448ba3d07c251ac587d2e3ac175a2bac07a4280e068c36ae24f484ec7b97d5e40e80b07a7090c6e7fa2c27dd85b90386f1ff0417e771c75849e6f573aa94255fc3b9b6bac620e3c6e14caac40accec28264d19856140f71a97640e65adab6ce41ad694a79ea26035c4cf099bc502c023a75d550bbb968c870bb3b4a3eeae2a5c8b987870205617396cad01f5284d25f4a37be0fdf9fd148a57f6eaa0f72a8062f24110c0fb02c3a29af87e7a75502084c87b9fd772e523e520da8891a425199e8aaf732a82b072600fd1384ba75820fa205a991254069bbbec13bb8a4f3793d87d8cb504da2ada7b8b406be95b427e89bdf5d0cfff67b1b0edc2349b1b72905bc33fa7eb04de712b3ed92a040592fae559af68e1f575087a57a2ce8fc73220dfdead964dcb24a968ec3666d662e9c45805dd37826e0803f2f25ce9ebf6a4748ced03eb927c4531417b32c4b07cc0d607a6bedc1db8721d5ca5bdd5cc3fe15b9272468b2bd4c279f4a5a23f1a9426b62484c8bb4af39f31800d9f0bc1712d4d3f00fdf2df96d947483413ab719716b99ff4edae7ac407ba6e85c6086b71681319b3babc6d35d643aad59301978b3fa64a86ac7afd1d38e72e33f6da09f199fa36ea4bbec166d3f8c4103d7e7eb3ec3a1b2e746eaf739f1d378a649ca8dfa087058bf41d3ae0e7759870d839f0f51b1996d331514f229f4ea2cbfe6530fb70303e6d35e51119d0cef5e34aa733a5f3b8e7c9de0eeb473c9009754c3ffe4218b29c95a8effe25289b44e5826b6adab1fd1e07c484116b71e429c3c77b19c05cb3172cde0faa980bdd43ec8681dc4a82b2c3d32dd8dc576e96281802f3e579693d719a3adcdd9dc362ab0ef49426e7485d0fdabd2a592374b757143320f29515471045af4d7b603d3551befe6f49dc032c496a8c9771b77b23775d47201d35f124723873b659d0d59ec0b692aadfbdfaab15e93737363355389e7bc987c4e702b39a68145098621b27ff7a259d3db0191c13e5d7ed199944627ca7408478ce0800683b4e83a5c344e226ef0d2d7e7f9aeadff0be448da34eb237dc6215e4c22b604569cb482ba61300e010d115dbee781c9994a95f6d16574aea95fd4debec3f58344e6848209a759f433387682e090aa663314a738d2ffb794dd548d771be9d806796e512a3078eb0232073051c52bb2edc005295ad42449f09763a2620686b5443dbd34172b759c70322cfc94fea17df7c95c17386e5a2ab7abf598a67e3249726308a515b8d11ceea994d601df236a9b217e8dbc589cf0167667689bd63b778acb95a01f15120bceaec4ea685b5a333ad24b2db702fdb180ed8721f9350cac6134ed776bbc19c6667a252de021d6c45b61f69f935a50c67c68d6bb240479bc92c4df7038bc362dec5713dae59efa2ee5a11ff21ec7429899ef4028a8ef46c1a3cd00cbddfbc2c0a123be384ee1f745b332dc65efd9fda5e45488b997b4ee533007c7a6c740dc2ccf6780707a9182090cf33f0664b85f5b857c8e412c52a2e5d0cb159e92d21ca92d968369137b805b45bc87a5b9e243fd7e5a52ea74e7f4afc216bad145044c5bdc4d75ac20f89155aeb86eab3beb3e1da33f0695aa91b24c43c8ea4392afc18bc28cb605f1c305cecb50177da4e3cb1fb548c69a75929b698d48a33bf6254c7aa7c266b7419b10790b95b71f025fa086c5155d554e656ab08c033fa291de08a3294e814346259fad5e535c568f8a3c64c1c928131f62d863106356ec4c7cd4d224587aaacd60b9807a33d0851234e263e9f7860e8436069f42dac9469db2a3949d009c19e66b251c57a234a55f69b66fecd722058e1aaf7d636f99173a8fe470f289864a2bd0fbfc20e165b6b52078ac985913ee71f89c89ef36acd725d77bbcad1a89502438feebc8efa689537106cabffb6b416ee6258fcf0b8d484c34afb0b694e40d192fdd39551c61587e0015d9d257f84722c32047854de45d4715f90c75ea682efe216465c3ff533a5c5cc83db56dcf8d16e640dac2cd6bce39d72df296dcee2ff58760aba42e65f1d5a569571ae9b27f89b0eb1749616e3ba2bb476d633a1551726b1e718c7f08872fde8d4d4b1c2418cf593d5f56bd57dc6670c589da9c58d989807afd479a233b69db1f0335d96c437e20df37f11d630b0188e26e2f5f634de0dc267470058ca5e95bb56cf03e93391e1fd764c44b7f0ac1a4e45eba38b32369a174f8da11bf527bcfeeea86b490071ba4a3f6fb341dae77b810a3843d72d99cc0b02e11526fbb30dfcfc2a9f53fb835e30a30a942d2ef54eb04fc6625c976c8d4103f8b4e04433be45b5339ce25a74d54f4f0a602e567d56e17539733cde534b788063c48fa58e5e53127cd72e827141c92fe6f104307d542ee3e9c877ae53dc4473076f7a598c89b375fdf901091064301624b71de9afb264079ae61a56f9212d2e1cff10b883076b2622ad834c3f154fc58bd0419795ab48c98418cd9da89b994be457f2f4eef0ba08593dfce73d1a38c50e5d8a442b262c6318696ff72fc7b063b202695c9eed7cbbe9db9a7d8d7b65304471b640ac5d0d74965e2866713920689bb96dc305b3eb9054272c898e19c9c9c28543b1b982dcfc6857694abd43c4a0cae76ebe0ecd912b7453255eba3036c630a57b96e2bc9b2054d033972beb0d55b36ea5121aff386bdb97ab85195107d1a6adac92e9f312b9cdb3b3731df3d6c048e8372330c04d09debcc34b873e5c980c8f871da71c05115c88621c976dd5fc86b0c54d3f6052886e8ff365e10b0d14f50b1a5bf04f69ad11d8f3a5e67fad80cf66a1d1338cd1785a99b151a1d03e3dd101cd7ffc2fc7a993aaec570258576cdbefd63353aaa30cc01fc5d0d7d2795f82c928eb31570788f9d80101744a6a06f9d8a1b55638586baa75bbe60394af314a41e1a236534657be06d305667bde11c41255e1c5951ef7b847facb5dece9682f233ddbebdfd0b1452c40418322f5052047cf79fd59061ff658885934874cbc241f0aaeee9082acace5430c6722c36fd02006ab06975da0784eb52e52a3c6b2019734e8a13f3fd1a55855352070eaea7a47a82f883604b4d076780aa9c925b131d5e63f2876eb6a077eec539fed2e0cc0b19a9be09476f21ff99844d5ea08b894e084410f2b4eaca232bf92e42ae179f029a184b977d196d0249dd914f358af0398a3fb38c6c044f005cf5535b9889d290f4f387977268e4c67a5ade77d2f99b09dac61e93b344cb44e930ee9cd259611cb3fbf87035d5bb12d31b40da4838451695a9cbdcf28102581c246224d2db9edf8b77862c788d1ba12bfaa92abdd6d8320376386f25c48aa2b1488b090cc5b6b291a752c0b3b9619c011b7f726a30d987ae5cc193b171e25fc613ef23386fef6308c812afd016cb0fc71372858084670a1824dcd4abdbe165e68e20a4b23e1d13432e6c3ed66d77e95ec838342a58413a795ea4a563d37dd464713a8d33e31f3847eba2a1311bdb649791c4fc9802ba3a2e96b361dc6ad84b4b218ec87cd07e8158d59767f0a30195adf462380dcbfed355b53e99d6dcac17b05907a9ca66e71a19db74f514fd18095fb9294450da571b2ef61ddc2bca1aed6d3f37a3d3cafe901c8fa22dd1e4371c3298c10e5d6b65e850c743b76835471bb636cd442a03486bf76a803e198c26bf3509e46d9d98647839be1e84cc63ff2972c508f87858284f64bddbb1f2751987a3746d809fe149c36dbf701c4bb163cc67c572a961ca7c442d30df8da0f6aba250003090cd5fb119cb873d8a87020c0367806ad43db9a121a4c7132c0ba41f55ee2237193ada4d4bf2ad18741dcc98616dabeb9155af609d0d2abace268c88b2c808f5a270954b180168d7806caf2917742020a3e42c257a854dddc68534de1bc133d630d685d540542e9a4ab64f84ed76d9f76bb0ebd8264205d55e9128152eeb7ecb721e2d5402859b909dd55faab105889af8fe4dbc82c7c87612f857e86c4c54b3c71349b7b94e11c3c1c4fedd3feff99ef1f5b3f9e5a38b381d78b9cfad37aedc48651fc1dc709b52e888896f11a3f5c02b56fb7ab4bb8596eb178dd78029fb03bd03e3cacf9d0848d323a825811f78ffb3dfd0c3080ddf513074b6a46d45960d9cbbb2b620ef052b0c675429732219c4027299b7909f9d2a1d0512061a17e411830e71088845df85db774d39ce91e665e703182041fa626015567e1db0787225d1916e710d61dfc31fd7745b48ba90faa559c76e097ebdeca22427ca89cc0035336d472518c12db42fcfb177ac78be7d712fd5dd8944cfb32e8c1e044afae959e4e16c96f8371e13612cb670b9867f7819d5d0d0adcd0c37e30f4865f2ffaaced9923a1a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4d2f6e82836e72d59d554a60045c6889052d03cc21235b1354f7a47e7311dcc8bf294f5a78521af1b76148394a8d4773f8a77f3366d24fd0a01fb379a7a682f038990686645f434b8e8e0ba8028facf725bd9598f6937dfb2d5392138c7a7a9024dc60aebd54d2f9cdc85bfd0992e5a88dd93c6eaaf7f47317d0ea04abfa3a85e5930fd00efb13a6112944011513760049cd3f245b6ff81790b5ea24fe9f9a40d729332b99afc44d9a6afd21bf61ec977b4fda82667b7300bec6fb926c3d2effc4936ea7f7793c1bbb481c5b8b0c1298a3f0619aafe360997899326806429795980bc6d98df9e1b1bbf902f479efa4476f3533faa48b207c69bb4efcdd4b00128e5c1c9ad7f441c1fe5adf3a395f3a466e6aaf8884a06ac79e18399e999616e7f38c141589ef04b08c423dcab0dcba0723dd364b5d019588549243542710a815ca054fca07a3c72d49acb2fbcf10e9c9b03fca5219dd88985a572271d725539269aa9040f10d1a64d9eb26e8d9423df6f002bc4fd366b719a96310866cec9880f7cf43a0a55b7aa988b14b5a2b763b75f19032eb70e29303ef8427040cb9337efcea8a77d9a100982cb43dbba85a98927b3f5f1ba23a603a7f11b49a002418ac6e8cc959614c7786993ec3207051e79f1b5fa65e350f53fc80bcbda1b32bc2382ded8027c87babc5c80042ee6f5610f397b2a3a105f1f87138caacbba2cbb59577bf81e27e20a13132950c24d419362332fd986c9848c9accee8487aae0f995f934bbf0a8333d7b4d674c8855ccc701fdf0e17c7eeeb50c4dc2fb5a0335f22180a16cc700d8f4d189d8b0f28a1c5c88955b0faf8ffd0c6b0289551cb235f22bbee4f4f175e8e59efc988f030f35e3fdde4c1b4f3ade308a549d76071286aac6f5ce7d20fbadf2efd7129b3b97d3fc035d1eddeab3bbb9772d7b577eaeb553893d596feb446f635777053b039b495a8e0dbccda7743f7b2e81457f622533640f818d502ae1b25ef49b389b58d1b82bfcde1111ee9476f93ebe1ba6a7f75b082d4d713dca57bf152eb5f9053d016ac90aeb761b3193ddf7c7994a55dcaa1d2a00cbd729b8a4cff9f942810f2544242cf66965912fbba8b8410a686172162c030235f2a8239e25c0bbc765dd54d54bbcc99854be35de751714f4841773f1df01958a969f47f12d8be1520231d817ee1a9b32d4e61371de29def5642094d9798392526c50cb33df377405715900c43340e6d4df1a13c672ef63221725c982d540323b24f3609a30e4340da0e28f09a5b3b730690e8370642b6a2b871932d12fe2b843a3fbb3095a80bf9c095606e8549bd7ebc54dab9ea2900c015e0697537c161090fdad22b40188c3a928c3fa01d3151e809df0cdba107870de7b38648d91fd5955ca11e133ca8f0683a7e687f443850e7961304a17709700489a4ed34eaf18f9ffadf526f2491624ff4fd49b2a51856c4b0185392bca222c22e817db6d6fb7f94437415910f24dfcb8c59009ebc703fccc7d9878f767c4ef1729023ce6a754b0584a0a8b78e34ccb27ed2b6c85ca64760344b9b6825bdb704c5708037e1b8c0a8e52b4212898aa2184d8c212c8003c2f90b555a8985ee4b3b2b541c7e6c5b598a008b084e05cb6b2c39ccb06790e97fdfd1ab2fe40007a6ec5bc74ef39ba8f68e919760f3018408fe5ec21a313f9a60e0aa19201f3ade58fe46144f1623a532cae0a8150da92b251d65884b5223b49d316780345b000e3ed97a64cdf738b43ac2627e3ee53cc14c5cfdb423f8689f5140943d9383389517a34bb7b638dbf9239a3834bfa56e43eb5aa4d4500bd4c5c8017b0ed81f1511a971b710ab57d03510ed3ce91424ca6714811de62f6713cf2c743d37f1080f4606555fc464985055ef709bc2582388dea43e25daf653df3e5adbc45e672f3eb8b0d0a9da42c62eeb1b30c458b4f243a731e3ae36d51da9b97baa9983c30f98acb9abec9554952bee8a4d40e8befe7591c65ced1f7534c55162be077f66113684309c517ad36419915e8698860098bc415e13ca9ad1b6e27bd68a041503f27a2c5f28fd72faf9ebce7588a7abd6b5e7f0c47ba9e34269d4e92fad1f5937eb4196ee7080ca6e9ef9a5400934ae451057e7b453806060ac70accd011ab10120648b3bd3121fddceae294a9e634fc23f7db005fdbeafde6469bcf77d1677260336e5f4d1fa6abe461e2406be9aeeb62e194f92cd45295341dd6dc20fac4ed1450ba623712a5376a98b7e35fa58c51d1a703255891ca20002b1e05ced29618e5d5f5dc3e8f1e4fd50ad3fe7a11f08110bad90d5a4407d069a40cee41baf71a4532e15f490b5bf66de26ad25b13a2776007d6d2276ddbffabd335ee6e915c6f456647cf3e2c46562ddaadc3f7552266d02a76110084e0d1861569fc4377fc788bf04834d12cc8d16b5dffd694caafc3c232ebb8c0843663853bf14f763c53e41ea3d0c47982e4c690014d6a3e76f350996afa3841cd0d789854644d91eecad9ff53bcff10f01c5da661de8080d56ab73fd7b0650c9701d768a3187d7eafcb659f654c6477115436934b4e3e7826c3c026f665be722c9d1c0f2b87612831500903e96b2ff872b4281967b14a891f5524f6f24a7d13d1d8c6309257328195f6a10a7546b2b63af837c5c7f9110884752854e28bbcf94e9946f78d40a1c21f8643f7624338406bfcdd4271868b56990728507e86bf6321f914ebaf9a6c8dabe3e49a43ba3f0c77579e626f4fb9bf93447ba3442b8a7c0c4f8cfe927279029bb4ac115ec66fa3258970d89d5e24c3992e88ee815d4d0b890d35d36c772ee0a601979852846d83d44e2b0a8661ecf60efac0e36c5aa4750fa76eb86695463c90d9f3b2be6a82c4dc4b8019e44cdd5702c5c80b07d3e0e4a7df57bf0093fe7a2decc9d2273923ad4ec666ebbf6745b7def6d492819d7aa9007c3db3426c6c306352058ce3a56302014bba55d5e683b8bf2b3bb1d156edf2721c97fdc948717edb6026368c87f38842d5ebadf2677192c6fa507793915d64104714148cf0e0188197efc90d32af918587810827c6ca55fd73392d14f9ab35af81f67e962650af868708f46d27ccc6afca07bd73155f8dc0439704dcc937b6c1b99d7698033feb3f0949b6ae2ad123613e5228b04969c2fda04fa6713f5ec3929562a44055e7a9c365a8e01ee92211f7aaa6508680b1709a7b916298db481dac34d6756a032500b96ca99f87020d6d780a7530cc428dd4cbf61b65f43d79532ac72212f7cf1d186c2121d9cf66cadb2037bd6b22de0d120c63de79ee75c30136b5ae018110a8a133b4ad251178426defa098858bfd5fb1f16f86f821425371ba7ef07d4f76e02658bcd31d71fb671791dbef9894503bf448b88b939290265befb5bf3e68b8a3787aa788742e3a3083d74e8aa3a06d9bd68caa395c04481511ad7870ecf595d9a7e600268743e47ce1b5481b2332a99640d69df5b6f5a88c5de87e509ad549b55bcf57e3eee843d704bce67c7138a73a95699f62b5466bd2ea1e426d844ea8ed95a72aa52f05b0c9a70b27cac83a01e0aedd6a11ebb870ab5158f916a4db78d7636d29902d4ee187783716b666edfe3e86221a3321a1d95caebbccf9bc0ade07432f2d3ad6f68e5342075d56abae1e8181befa0e868bc5aec050a8c4200a3efc70cbb235865e6192bb0f23807e327b3ca123a093a087cc2a5725c224f2d58634270d5b0017f47ecbeedaae0aef4add1d505e1764b62f24a1f2b4c474a5b38fd6c2c2e074c83f76f30f0f620ef83d2c78236b5185aaa55adee2eb8b91ccf54b1d6edc56ce829cdf4388710f706a9bbb56bba3c9b298178c3bb36a36601e4afd5b6314ba5419e06c8b42a685f58bf52e556fb6c7f15e99b9908f628d6419242b2aa4049e6f58ba8ee04b4d74eccd5fc8f2351649a13824e0df237c2b4e179a18d59cf5f4e409f8db032a3b776c88d7d81dd4e4c39bf738ee836bc8b7ad318430507a5f2b77c0633046bd181bb7c60c7001949f9485717e2ac3a02e7aaf79e8f8ac1a7c4883d730811862c2c369c148760a78cc07db959f29775234d90a50109a4bd366364f2807c9d70ce12a07eb5a4e6bbbeeb0af93ad621223eeba1d0324a923554a2b1c4f0859fcbda876e0dc8bcf8d9f156980ffd959c0045436eeebe9c3ca71a1a96088159f48c660e78415ad8e51b887dd4561d2a73be40655721eb556263ae194d83538fa18218835eb5edcc1bcf49826d6175d70af63b60aa6886b4fa674f401f010961d04e73be3644941058270fbbb7cef3efac1a8ec5d17d66ae6a0e6468f2f06dec218ec270c5281f810e89151e2dda14c6e14606499c7d5d0ddcb30dc303a9bfead58e3da7a5474ad5add4374b7e41de58b5f4ea3e4178169080cd1c4f0e3333cb9991dffb3748aa4f8663a999c7d2caba129833de4b494c33d6dba929d1f2758d9af4471a344f1784425d1aa19e6ecd56c85ccbefb1309d1f95d1a7b9fc251038b9c94ac2516e38ec00d91c6cdba22fd30b9d716e0b889973ef0bfcaf477ba23c0664b002e0c8d17cc58f31e14d27e2381cbad793732935349050002a957d39b27d0e109637674bc440644167ad0961ae5427cfacee624cdd533a98266075f90c8a5d82346aba79d7bc5e29d824fcd021428a12ead963f4e535b835e1dc0779e749f5416aa1be66806c2e1da438dc110abf8999d6b4670f347726f02604b30a826fef48eadae8c2e68bab395b0c2e9527b32f9587659b367ed5d6db03f2dab3c6b4ccb4189bdbc34f1100e639cf2f51d2e17c4c8e80c123875ace05ff9b3142b484ab2b2d30ea256913a987bd0a528badf83c2cee5c7f43643b056c73c11e803f909d445ebf769a8ec8399142c2842129435936c7782bee287baa0c36d8a89b816ece67f1ed1ae598dd1d14f1860a2874b520780ee0ad50064214aee1d89bdf8ce9b74296ce47db709aa06234bd34bcfdaf88aec8d9c1c2d75554f22b253457738885803f487c3bbf08dd08dc6c11106c3a9e5bc2353d662198cd055b55dcad478c843f9672ee29ffcb39731f13a2bc97ffe0cd8c3599bf8b66bae3f2219965e32167eb3dd36eddf7499b4930ae2d54b097a866d01c3a8660abbb95dac7967fe739ff81cf5f8d67316ab5cab026858484bd3167b188f3ecf7c4adacc78f83df3d30e6917f86aaa183679d9b998005d37f1849ae9997498f033da6ccc5876a912dd80a3a0ca7f22078732958b66bf676c960a88fb5b035c49333374a7d3811da880b3dc5e78788050264997a5b3a251a28ef6bb5c344d0271dfad66fcca7559ee775bb1ca4863ab4350f0350c7426af0ec9f73b16a252217ed468e7a9d17ef28f1ddfa406a4478ddd3719e9e97d2974976a378bd0e270c7011ac09f5a760ba8ea558541fe5f09c06bb875fc21202953df70c0fecb46eb2770a9f64d2397855bea3a85c7634316b805d94ec31b13835ddcb71f2d0566b524bfe6de75b214c875d11d040898db93764da1c8c7bfec490e208fde48b4ff4f9630fee89c44e5fed4ead474c2cccfb5fe77b35a71dc973e95c77f3362365ba62f225093c78f246702ec659edf89b72b47426fc8aeff8cdc0f47f7e2354dd1b0e25ca3db77c53f17673d2e2241cb3dd1ad6c7f5b252518f1d1d9ed145650f158603874466e77e2e6e2bf4589f626af5f75b6617961cbfd49b3fd3609552910d52d311482f3880552074b9334a9eddc7e52560c2503d0aa987f4dda6daf7edbd81c093465fe982e32b487a1e3b6066c99de328526aa3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7d31f8afdab7630c04232a0e546ed60a322162ed5746ed17384332fce93ac56d415df465643dcc456077dff39da5381b0dd678fb4f82bd8303508b68870573f171dfb3ed3ff6e78954049eebef0a712374dba114246e8a1d774fbd6729a4d967da5b55cc905392356b13c56f87d3eb9f371bbe5cb1e03e6b6720a244c6f8d898aab23237daeb013f6a12ff08221e178eaa644a1c1207416b236101158f271c31d693ce606ddb66075c4c560f46b82ffc904c10208ba1bcca1298efd25d4be3afc1074b1c14a994fd8434d3311a3efb7a7bb1ad64d5da6c1caae47a935a2badb49268ddd19cb83a59a9629616dd7affbf1440bce0ba547aa856f563f309f828c617e231ee530c036df3513bf6d3b52c5146b879836c0f0d2c462461302a674230b3c4b32d02a74aca4792a5be57890fb0a7d7748b123dfd83d0f4049f99a694ac62e3791006728a877e3941bcb20a69b29966bd768bb820c3bd388ce55634e307ae7f957cfab7b0cf551eeeb65f6056c20589d99f1f226bdecd99fa229f3bf3a1655b756fdb1a80be44c4e8e4d1833dd055d41c2c477f594014224c65854204a878599b5507b6481e8d106720fc5ebe336347f8b6c1118ddc621f41871ff142fe4c6386885d325f26ca80409b280c267563e8af28bc72795ae2c6e759026f01f89d73be30ef3df82ffac454fd037a2f5936c3092e19390a070536132a373f614f75d3c3c9d0d9c8358d393085b7e833998202a62841080e3991cb37375224f23aa735357ccd0055b915f0ee1438f227b031f6f10a414c4450e0f03d41cd62c6b21017cd29024b24311ed1b8c79ac39cbe329f6a08d221d94b6b6fce06f3516b8bf11841b6bbc16f719a57aee43b991cd49fc68cf0fd54cca1115c884438d0e9ddfb9e0a77c2178c017ef506cd906fbbe475eaa10428867d7e30f462ff92757a8898046b8780ec79c82092cdb90416950cc60b4b5d2c44b903ba75686d180b75f83477e7421bed534131dd448a5caf35275662b11d595355878c6d70298fbb236c70b6b92407a6910a96262136a0333a2025b53735d46800b5ea3c2fe1993882c79b600c9b63f64067b86285a4a3eb6a292cf81235323a4376a6c0aa6f4ede8a23d3ac69d55e8f08f03b969d973a4404d193d7b812d65ce74eaa1c89087a9618b915b89047721c76775fda3f03ad8c38a65fec2f3aa1b403b196c1c862e54e2f9861de421baaf7c9b190ee0fe4b470827b8e003308388f66b9c7746384a39bc49d5ba97ae64cac6a72cbee0f1ad79a8b61d5b657c610ef817ea9dc481cbaae2e1f8f5546ff717ee7d0c76122e82f5910573c66c5ec0a1068f59a0fd8e30e904760b0d57e5dd52fdf8e8a1242f09f2735b300c6b1b175b024b691be6b21fc5078e43e99c9c1e30e7ea81dea6655d7c002abd542f9795c4715a67a9d7aba559137f053535be1b8bd08040f3d952691a11c8ead3494e35a283f0491fdc84b9e89c76577978a54c44e8d51b99e25181bd7dfd6cb26c749c1e7cdcd2acdbcc0f27fadad99884cfa5aefa9e632338551a027b2d83579bc95788aa424febdc61764203d84a7a1f21af186438e124c24f06a4f514703d8a40371d0d57327632c473137ce7eff97413775ab7ec6e4480abfdb2056e74a54fe7a1b5ac5e50d789c5d38872146b6021d870fd23aa3e0aa451b52099c5b806d8e4bec3516a7fbc7851ccaeb12195f73a90dee92c28336002c5301087ed15c2b408e74ed4ba298f266627d4992e4c352169bd3b7b05b8e930ccfd4e88cdb33ca37179835255bd8c663b679c2e476f624c110a66d538c105ed5b8d83a7b94ed64010c6aa7129474b39129f434dab9928540facd6e63fe404a7d5af6aa60010bdf4e6d843f497550e0d1dce4c48860593babb3b1f4f77ecf291c679338a5d7f9b6bc97898eec524731a0ae1fb7bd19c0fc91f5158a0cef7aa151ed73cf9181a9e11df5114e3de3d352f5e413eca05ba4e227a2979d6e675db3f56a915be578c0f76cca0ea376d2fc2ba654663ca447146595830d7c1475ad8afda0492cda4ce59dfce6d2130c3d4678735f43fdd3bd113198f36c98b07cd6fa9177898260b1909260750dbf453dba6e9eda76127ce99900e600cddb770a1dea5acc809752cdcee88119ccdddea736db477282fa192f5a9131f2cf8b35c2f9754db93f820a8b54fad4d0a580f691bf4fcfc09eda388aa4ddb99c91bc1846fb2e99fd4498d18918054c1b885e9512dfac7dc9116e5faca1b10d7b15b2e597beef497f1d45dd75df547b448253742adce62d1d2f8ea9e16ad3172d9eaa375e8c2630fb95b35d943795aaaba5b070bbbce553841632c288a79f982842f0dddd8ec0c4f87bc3a8f92aa799bdfbf050f3bd7ddc3e152a740bc04a7641b663bad7eedb6a03a13a8eb995453a31a718071f523428238ff8a3f93c6dda701f877672a098777e02c4195d17b00194cf3ab37e012658b8a9736af4ff2ece9960bad00b86aa5aa28c9cf16370dae91e5de7d44c8098626f05ed647ee864ae066ffc73997e916226b4191a7e14f0bab10ca3c3e87c6cca2189d45fe2790271713fa3a859d0b4a05fe5d1f1b8704b8b8de1d20b2d21347353576f5bb14782421f9035a0650bd7a62cc6e742d685ccdf8e1c328c9bc9d2d1eeba41e45d17f0914bf283fc22085e60479855c842453cc7c65dc86410b90009fe6c24ac634595f20b3a6e0f6539703510bcae3feadf02379d8e1006778329f6c010276b5b825c4544eeb8a196b00bbf6bf810550714e752ff87be97e2aec8e895d34c4f11c8a9e06ab66aa03aa449bf702ba0221f8b201f68975cdd635318f1a9f033ba203854eead5a818cec021621ff7bf293943656603992a744389ce676d5928e1ff4482df53cc4dad866ba23487936480b4f04eb394e79ac5defcec098fce7009254e3a062ce8178cdfaaabdad963f079d2c7ae6bc875704d8fe54483ab09a7e3048f5bc1518fa098ec0df1d21554d1f9653d7909b23007ef8307806631b01bb5cea37b8a03f4ace4a1a76eb68c9df7f386596b61f0c752c5228ee8f0a000d83c8a844fcfcc9985bd47151a26b5c6d2cf2240f26ac0efb89bb0af3eb85ea2de43f612a663f206a162680e6069030f79dc7349264b00a13a90b8fa0534dbce160ea5857c6c04c815527d747ebbd3b7e883038661447afeffd2718e24f66a906bc6b8566d1fecce193b822d9c3f859b3d8eb416a686d4ea6af9f3c3e4ff5f36fe929178da2242f79238cdb9ebf9c3b2b8ef35749343a02202bf950414f9c3ca8657d27596e461c54402ed6668127bafd30e207b4df1bfd39fd918edab055582e926f06507c222a7f0448c74598481d270c849304b957e7034cd0ff79a98a15f5c13a9159ee410151390062f7de3213b51ebc1cdb32f9fde768c2b1224ba34eb63f385e872f8f5453351bc2a8af4df282c30d50f4814f9a2a4bcab9b396c3533febf80afc898d76a465227baf33316f6a33efb955c9da94e2682e23bc92e97de846e8d9248f0e24ca98ce33d2bc6f48babaa20c656fca02dc1a39d3ba4165374748bea7a42c2d755e82340cac27fb2d975172538c15501341a548880df944e50322f89aa0606b7157194127500557cd4f65367dfa2a55488a79b4a13e3dca4cca4578019df9b87dd4b19795f10c713dd44b1d8f59708e9125ed11b4a3d7fff9978a9c1887d6f9b065d4e0e33e6b50e0676e38cdbaaf519cd0123788ffc455ff156a2394c46b5179cc3fe25f9b9cf4b627c3c2737e9e2f41e726381ae06381ca887d6907e9cc62cafa72946908cec3282c772594ad5cd5f59a303806e103d77b664604bc43a3e1ecc3dc13e458eed555d85c82910d9f5e2b19aacfae8717e1fc430c01b1e6410e1299745cedb30118be58d3b1b31b9501a658050ccec8a2c1993ef9c3a7ee63407f2c4fc8f37fd4041940c0b28a1654d3aefc0dad09e8a86d94991ca3310239a23194761fcadc5d34597f962b56b81567d290b6f396806891cbf1cf53e58c5d4b192402b85db3941c5ef08f61474fc3396f8a5b97307139b45c70871ff5a4359857afab203a6a4243e9c57985846f9082ed6284e331c60010e0401c2ac4fbedbe3a1a3444309f386e4ebdb3dc92da73b445efa2dffd24e99477ad2e0b59810925623d377d59efd872cd7a4f454d8f8227eb981d6b4c526dc9c462222a3559f674b4adbf17058d40aeacce7149e0d3d3014111d4d4bb365f929b5cd63b926c6daaf305d0fd1674a8c9c278fb6b6ca9a835bbddf4d4a3235bfa2784d259cad4170b74b6f0b80d9b3f1ac7b9f2e31643f739857dc083ac64157b501a100bec65d02a907c2d4cc8a1339440450cdcc712e45cbf731e7f175aaa6a78e8163c355896b1728d07ea90656139a7ee398eae117a6c88df2d902c5493b43e17317ea8b5e0bdacb36fa05822df7cfdfdf4586bd32468b351b9b9abaea219fd5316c405aaa9076bade456c840bf07f829510317c6c8fd2a1392a060fa922e59098a991555ec8cacb62db51e35fe55ae56f978a36a5acc8341cc55ffb0cd19c0d9389fbff18e7ab87564cf08b348e0f0d6239f30621c13540a57390a8760e75addea267c54ed08a6acf3935a60a8aadc5c9a8db243d94bb37242a531898b13205f81a9727ea1cf5c0ab752fb83caa72ec30ae9831ed3d942d26b88a2aefbbaa42c3d53850b30575de761a852dd14912d3c35754d6acc463dcc100bea4c99e832de7e6c5d0b4e0e9bdc8a6f644c0c804ca832c8161463fd930449ad7f8a2e1beb6970dcb456ad4882f5c805a2f5e7b091062b6460d0fb90d6e0520a320d33e8c03c88d5fd2b4ec2728e9a8af53274d622562e64a6ccfda930aa58d607ef7362670d86c26f1a8e1652a9f39ebada6c56c9ae057789a8cefa7b2573dec4a678c2dee70f3ab0b777ee197a2f9083e5f71aa4096e375c9119bef4831088832e2983a80e092f79e9bf67909e655bade3690d02899c180dfa607fa3e9b2def52ecd257d6d7950bb6e234c0149371aa9f33e08c7bf83716472b8b34603fc24d8aa38742e252905870e037ffbbd32249eb604687c91854b3dd245587fa4ef7d41a92ad327e2bc0f9bd4c5b125c963222e52f97bddd1eba93ef869316961f9cae0fb1fb543e9f722f11e9c68966774508fe6434cd7b5d53b902792c9dd811585990bbc6b407635b25992b5fbfe72737680e4798c698a2233951a7d373602423c4f5fffa90f966813910ab72eff3ca144d0fe675219bf2039c83530d0cf37ea4f950942d1c91bfa2495d4f5da13d842fe8176cd4fb60f7f4a045e400942e40f96c371c72415efb1811321937345a98f227fa7994af2cd7f8557d6f6ceb5228c0b3142476e88be299a1b1df4de0264dd177ed3b7a4f8873586f991051ccf8fcea62c9d4a8cf3bd428b8d6709ba90de21788e1069195c3ac26c03b502b6d25f83363a1a40b62a024756f98bcb64d2eb7f1b7b0a66febda6b320fe80994ddb4e97f4f087e22f1121a3cc34bfbca3f04b9b0fccca1b0a96f7a863f96a958a4d3bfbd34f6d79cefad1999dd7b8668dd9488b50d62c6c4ceed8bdd7e8cf21c5c3c50e19cddd57baa672a45477e642b224b798a5ad92ba406089a61509b3594514b1f0ee340987b5e10d5559f148b8ae26f5fd29c5f7a9bf03fd3e60397e7a1280ec56fb83cde2c76955a6b284853e527b993469c03022e3a1ec184d3abf51b68d525250e44bbf6143d211062a9605899e85d42af9b902d1acbc72af2a61817a64bf7812a3871352f79ba74483;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h39e048e124c43534abfb5e243b2f9fe9d4900259af6309953d54d95dbb602a83a3199446e498fb669c1d40a0a12bd54568149839f5c566bd8f24c34ca93e521f521a02a49ca9f0bd934ab0529219a268030966efff373bc10d7f4e23f4c15a950e40d9c4b2a3664140a5e90ca25aa9a7b672c0b349260663bfee470e6d4acdf592a365803d351b8857c16f434a6c16f0739a22cbde9e729d53f102822e2a875f6b9afa7fbdf485dff783060269bb617e7b13ac759220461fa12cece7e59208855cb74a194f93157a9ad989aa821de6463ac83a38e1a55a98755f2b48a4128d85fe5dc60b2f6db7d6356bd44fc30a23a051c7a903bc501ab1965964616398812443bbeb954247125c47b01a2af5c4d02e0949631f1ba225c2497506c3e89de1b4f6f62c7f76f3b1008368cbb731a055e9f9f18de530930801fdf60965aec8207d9eaf73dbb113264358c5abc5c9e870b455409eed22010223ee0a6e1bab4341815b222e1b2c8455f982fc56b6e252db7a65c45c8b6e791924b1eefd29ae0fc072b535c184df64c145433125e50dc75722e8a3e2b7d405739b3d2aca9bbd5f302faa3a99defa3a2745c262e2b02c3c0b421fb769f0c548b0e380e5c67c4d3d7f9917f390ef98c922107d5427a21bc05a5fd6ca9deff09a5a5e567be4f1cf4f265adc65087990228cf76a1ca8707ff64d7c364e0fea1fb2d47a709e16d091112199ac62f528321768061fe950d2e800eb0f0efc249e412f15c62a0eeaa5c3db9d09611d2556b7762135f8c10bca0cb86055eb0ee946d2f469bdeddf842766645662ffe25395c0bfd89db886ed075b515fe34fd9f10f8f032574d45cc613cdd6fddee6be034279d53d998b249dfb3e269ebf5d352225cccd103ad138fe4a8bc7fd1bb521a1a7c5ae81caf5b6e030fc65acd01ac43fd03d8eff9cc614a370f5b6813d9641ccdbc275537ac5d95c0c291b6477e00ffdada6377828aec9511e87666e6ba9f98de0448a88841cc3d1bd4f7fdaba9ac74d2d76edc214866ebd81024376700ac01ee58f2de56160bc0ecd93404161dc67076377a95832907b9e72b85b272684286c46de0fd904818b8b00bea89dc21fb604acd7d4c69ac172faca3ed126710da80b7ce344bbaaa9fac4f67a2e96783cfa4fbdd9b55fd5871719371b9661f34dd7556378e91b8219b8e5168a301aacf88fe6d1a86d1cd262c2f16e123ea60f8b214411ff315297f16d6cc7748968fa25ad93046403d012d6e4082fc0cb55eed26385623b18f0614386adab71be097a9f1be259a468da0ba7b526e9a6187462d05980acacdc7e1efc6a96f7a7ae984719ff3117b0451ec433a8f68919a9583d149e6f6299d0d94a0e7daddf909b6031b743c8bfe69aa21d004c2d256157cd356cf262fde8ff45969a6c87643d7683e0309919ba7ba611d8e9b6fb728e9c2880331e73be453851967106e06afb837a2d2a7175b32b56b6e1767d0d2872337bc46ce1ae75cf0b6bf673d259f71d7d5c2b85fc2b785615c983e9c2baf251d813338fde64add9de07143829e1ea5bcaa83348d3765c1637e1fa523562a6f22e9652ff1af874ea976b670b1d38e994c24f5ddef4e42ce93b030ba6d49b39e203bac3195ddd7b9f2939c3721ef3f28541fcce455201cd08f07893441581ec6dcff5d35ac4b141532b19272cac010c6e965329e5b26a74805add320113a99250f9f70a78f9a9d9d08824a8933eac14bd14477f3d003571e81565f61946b5d75db0849c4a7bd89a9ee14b1e8f2be57981fef14c535d1e371e1e3fccd405136a84c6f1b14bbe53c67b088ef9caf2b8e108fa206562672e71b05f8af119e604957a0f73907906ad6a20f049b71aa4cbb2567453c1b41a5c37e2a44ea0c49c7c7cc59dc776b6830af86be7f8c047059ec79b445f2c0a48b8469a4d09a8b8d2068ca96730641578116068c7349577fa0f4e07fc12efc87f5e69b9a54715106346f64c4197d486c95d44a50fc54e546b8199c72de42d792d01cd84d8d6ca77fc4a1ec16cfc6d992421eb49473bd139e7afef6ef727ef575934c69944f88cccf9865ccaae431a57cddfffa7405c6686947c32fc08e76d4ecef748dd775f1e576025371b35b5c2bb745b50432b18b826fa40d969ec288b28917cdfca1b12783ce595838c444dba5e4dc23c6aae2dd81e2d64b23c374b68fe22e57149a75bcfd6c82797bdd7f3a9ba344327482736e97f4f963ead8bebc054771ecbc625593c26a7224b3f7acf08d06edaf521fa7872d9e659988d274ba637cc5d73823ce7174fad457d8916bf2411f42515f22d414943c85cc6b9124b529078ab03911cdc5589b50e94a70baa90ed860a7fc0e4273a324e5e3d2205b70fcb0ba8761c10a0974c5b5abccb8f4d74678720ab31ce42400d81a94da67507d5b3403446d03201e58727c7c36bdec607d3e638679e4a09ee2379609d4bb05c0a3e34d7d8e09b54bb7f32b7dd0b4a0b589f970ab8addea983689d365b2ba0434839ff0852d9d0bc6b41c7386dc5adcbf5204879d5f62686f9cc646dcc729c97d270775df21da2d5b0ea31a533e00b86f8de666e34b8c6bff49c8cd8619de18a6d67427abd0e4d0b0b9f22ba394af35c0f70de76105d9a28c7c8625aae9cfce0db36e1ebfde9a5a7ed4d048896953302eecf55ec80016609c9b5077e508424aa5115c61ada7e110108f890e906f58bffbc0889a8fbca75d8f1d106467942ff5dfe63b33eef2533f7255ffa5bf6719e0861183c2cfdbec1359b8af58edec7e050580be89abdcb9310da01e02b8256ee0614bc51ace72f08d71e16431831fbeb5d92f877963de051fb38e6ad165f2c0e2221f2743a6003724af2b418ef9fe354e197a1cc201c2a3459ba259f449e6b5cdbb47fc6416ac96ec08c80f1197170c921af383285ea7f4222a2a045bbef25744e7a07e9f73dafcb8e509d5b851473aa28ef240a8b1a2cda2abe21df3e101e6d5623cd4693c5435a4adbea508ad589d6bb3ccfb22b4fb3f00ea745a7da3aff7e5a03ffead0e257d22fe706562108f6bf3d58b82169b87f276ed48cd042ccca4770f3bd1862c6e69c07b3bbfad2cd8b1baa86b0e1d33226ccec9b24762701d617d9f54bddcc168835d0bcf721765f4dd36f0834de58808aa42b800137b232ffa8d0496b673cb166460c47b388595b3325c263f054d6fee744ca8cee68383aa210089643dad33ca7f3c3e8bbe8bfeae4fada20d4fd7dd2fb1452163f43c11c07eac55d9c552c1663e3b64284e82fad415b1031f120d7e37a514d6e58adde93f2d3a5d6fb0840c2af9a75e2a10e1d82946f5817653852c740d1a8d6bde9197c681fa95c4ffc08777c1c1b5aa988f280f0270e5d51468c69a11b16fd5fe8f934ac49d49d17926cf621007f9c66b608669d8b132015f1f1a55b53d1af36b3a4d511975ef01f77ae394c6ab23c0e9a6b7c6f6ff75b0a07cfdbc711cd0b6a7da0b93bca76066cee9f6b53109991f94086b96f18e289366750bbb633e0a71966d563ce577f1f0dc16ac53ded4bedac7335d1e34b97f36fa345064126d49941c49a0ea281796a4da7d139c1b6e8898ee9267133f15fabf95a54c5168562457774c2ee5e8202ca8f1fdda50e2aa67d4730fd6f32a6c0201472b707d9e002d2f941e8e4da539155d8b079c66dd4844e10c6aeecd7b5f1fd936542edbfe7b5b0f2e4e1a1d8845ceb67a624bc5de99974237af9e7de6507c1904d377c9c599291f4f37c11dc2329d2500617588dae6f315636133ba604d17a1df36674e05f9889c6546f84095bb4bc4755452ad0b52ae87b88f6a4e0acb41ff389b5e59d68b161c68527ffe8580fe78ebd07849266d7ab2434c3c2b5db8107c3a3e47bcf4d15bdbeeaf1d4a510058eb96a5af24c8b7b6295d46c9863620d11edc7e8c565c9bb06f9944e9f879ed9fad340080a765b9b179b7276e0627bf3d743e7b57dbf6d936ddfbd2146f3eb6dfc20045a6d80a404343f31a5dd6d8b816ad12796079fdf8d1b8da79a2cf76e6d08ceaaa35b9c259a1fcbccdbea7be82d1d650c8de45b007d128ec648e93b6e626df9e0ad0271a413e4b83fdb62db31d5d4c1e3ea1a90ff768b17c221a46e029a0a792e35bf0dce8922de46bf3c82ee7bb0646f3dc9764c6d6b76e6698bf9550d08db25b92597dda1fdb7c2565fc0cc57615851d38bc654a6103e15dbe438a1455a9794c665b3ed906c0b03aa0d7197281f9724781aeb490d2613ab7c561c7ba1204284672a7d438ef8d8e3d1e478935b0ad26ff8d6022652d69647b750f446fc9709c1c29329a97f2453ac42cacb96251f339c496dfd7d4893510b3b8994e34f3cf17aedcc8c5394de6fa95349f47d0f61b5e511183edd8b5bb841e988726895a0f54e04fc71c088fb60ca872a9e60d31e5cd03bea2e8b02cd1e944e10dbd44e7357249979c8f960c83207e7d84d2882a273a1f7c3ef64a5610cbd32c77128261942b471cf00724003b809953631551d3790599101d381e2b3dcf2a41b232967a94538c290602eab21b63361eb9c4bb3697095a2ab23ab13db7cc1d90a32f15e291e8fc45f85826f939e119e8662f556ed40283b864b72c090ce741e203ace4aa555492da694a24d4b93d511f0d4a37d97af807db9cffd1bb52eade47bdb77437212855afa875176165ffab38dd5289d3e1e678cc644a0b6b5181ac92d67def8179e73f5c77793632e1a32f47c7030a5ef33a4abc11de1983f904fc1eba64dedf32cfeaf52c1a9866c982f3e11ea57e9e597c066498234ac52684586915bf70bf025e73f6877c933c55ff6cbbaa2775c44bec6a1daa12354cab21bcb4bacfe336189bf6d75a1ef9b911147e6791d01cce5f5c31d871d842df6329563f596715fdea00b826635d0aa7dca8c2eb1ee3df7943fd46c29e9d5b2abe035c5efc5e6ae58d8b7973a12baeada90f5eb919123c8ccabd0ea372974af3ac06d3ab7f0590375e55bcc7224784f1b4dd5206d7c72604e1783eaedd1c3dadab0f472f9cddbf32d41f200089b3a51b4cf44584c52cfecf0c4bb9cd79a79a7b0d0c1826a6eeb02cd37c1fc76f6d8ac2e2db8fb174347a3d722f9472b7b6ae7d004fbf2adea88f742ab6ab08007ee4ac92769b5e118e5b2ce43d005c99caa7c9cd27c2b905fddeb95fc5a1cdbc79c75fac20ccc433fa179063b6b7e0a2af1c8b88a893af4ce5d65fce987548b0be51db4a8dfdf739a19e054c8cb5ac0b43d91b92ed25cdf0a34f5d1f0f885ed0badd76a3a8ba1f1bc64f9c313a66d2c950e447ae321b793784bf875eab27e80bd8489afa5b303fa77916df37b41ddd4bbbce511fd79362bc0974bf752767bff308823c898399e939ced0a0b02b673a370ac46037cdfb1ad018a2e5e9c0437f80bf0db8bdec61f65c2c4fc07e04679d37bdfc5fe0977ad0d62d85ac05174d7f91c7824a892036a298d54b74b908b8cc0d54f180b44c3ae6a7971d01c906b421a608d64f62ac00a9a146c66aa2aa9564749259ae1f766996c13778fec6c48b6df96ed52c802fd0310f10eb21939ade59332fb1de6d577b5b3e44f05dd95e50b7868cb3b4804cb2689a3a4a46c6fa540431dc2bd9c85ffa0d9d30effe10f8031efc0d5bd7e5dd33825fee91a41f84aedb08fe17d8d18c0e02ae38793edb0a89dee541b11bf2d6335cbf9c16fbf03d708c13072e324c98fac921d5dbd9b14ff586d493fdf22fb2301cf697dd7c4a62223f6bd020232ee6d2163be3a0457a1e219fc5f093f5d3661d13a14ffb0943b980c6712b0aa44f2991b90c2239b84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1db734fed9c3b4e15c08433005acd1a503204da98af85b8a4cda475fb6cda30d027431391c27d02753cdd95350a034ee1175f510fc47e149f5610f1d70a1c83393531ca10d7d4a97bbbd16d7e43558603b97da309bba8abc216f882df2a6689c610fe356c9825de18599fe783880ca6aea5c5363fdf8e6bbeb773f86863b5b47837a5fe02748b8eb4846ebdafc58822fcc56c61f170a1e56dbe35b998edf0bf94504915b6ab0becf28d8deefdbc74927dad002c79497495c9f67f34e32a8bde8a53cf3957b176e3021030db5073979249fa3353912805f1bb2202b29f1b99df3f03a48894434dce533191f12a5f4dfeafc382d4109e1c4a7be250719a70b669cc88e19fbee025197f1e059a3f5fe56efaf5bf5cecae8170c1c307fa38eef2da063a439d8047f26ddedc81106396f17d2b67035e10772722270342f5af2f190071882e1fe30351f51aaa65ff1516de0cc11f244c9f717dc2ca857a54fb0620523bf959c89c64e2aa6a8c3b9d7d1342745db24ecd90bf5cc48ab0857231940753198ee511a48ad18f6a6b7b46ecc3408a3dceec13a28afccf9b0503311cf727f1c7c9cde03f41a5a8c40733c6df36d8ec8e6d6d1d1ab72cc421e522454525bb95f69860d79e1a4916b610eb8c0eb1de906ea952116197f8382ae0406a49338d77c8d268c4ade71c8a8cfefd9f2d5f2383c260d93be9551c2126cf8a45f9481d3a258f81e2c819890dee25ef0d28e911154a551d355bb7e9b3878d2b5200b0a2b440959b3df37383ad3648f08f9128aed3e6884fb313b6b164426fc09d133a7b5ba7a2f56e4ac42985c6bc7f2e9a7f93cd3df12e79a22bd113fbef79048937801f2097ad1c73d50f5123f3ccf3c9a8f6e1fa689e37ba895e1cebabe58257fdcb78bebebbade5e3532a7235885856e760ef2f286c3a3604a2c59236e766f674dc2143275ad66bf1c577c07b6a80aefb9b65d9990c958f649c7b271c77bbbba93dd50eaa571868a286160c7b612f7dbb9907476c17b28b30512dc7cdcfd66810d94de7382d7a38cde1677e6638cfde3ad1cff2a2ad5ff5c769d8e884c9d7d6f603158d525ab4d9729f174e708ce9e11dd610e36f405e6214dd4b064427fbf8372920f0ba05cdeac3dbf70dc069807507ff2608cf7581777b61e6502854e7371b490ea42fd9ed96ead403be2ad4f8426fe5521ec1a7a2e2fd670ce00c35a43513d85a7c9ab8b6e146a2566c7567d5de3fca02fe14a4efcd7f57e32ac01c20824d333113b5537c7cfd4126733b4177a6e87ed57a4ecdd6d94c0a3f23d8c0c5ae4a1ce22fbafe877cc4bb7f7692d6165f72becc38a5a51c37f17f176b9d1055cec531dde3d9ae91195160f820b6b86b2ebddf074e0929b212fed3d6bd8c277fab880cda11d380bfc70b963e393816242d653b74ea7ca1833e6329584dcef460f103864d3bde06226c7dd4572bd38193aca65ec23712c561be02dc4f4524c7ef0d298a1c236ac3fe438cc35d04289a9063345a4937a9707579873e5143b0e17be2a181fb47368a27b5ad7be4f7ce059d381a7d41c00d73ac9bfbefb95d06222ca06d223aeae939ef37ec82a34b420f806d97439cbe9ae06fa6a48827508d53a23d131cb4087c19dd16736d5242bd2c1cc5d7b59b415041f9840f7bb34afd5dfbf4b6dcf0d84d34542f48d0eb96c84cfda8f09393cc1cfc07e448526006f9af1049f9ab422007644c66c312b1c169194fa7333c77a91778d8355e51cdb7e0ca76ed50f6be4778208f76790a058895d80c78210721ff7064ea77cb81e90fbe37ac9013994c89411811a14f1e43f7d818914f5e1822281463a8dcdcc63e1d05025c94f3a03ac436bb06c9f647b1bdee96bcd9eb16230b1f619244dec86da356d074c216ec351f7de5384808773b8e0d288b51d6ff284c6e30f8f4c9ad5f863a54646351b37308dc17fafc3deb58698ae9625cf03187a097f0ae578b391e108c44ddaeff4454daed702916514021162588e7ea30e5d874aaae01a2299e37f0aae72decff6ee5db03d700705ed4bcd34cf8b27a2f39b0e876856a5e00f5a938715998f99314c3e7a68b87ef0cb878d11a0402a1356fafb13b377ff17bcdf068c68a24f77ba632f191d7234e0a1562b62196b41ede938cf0cfe82cc015d284f2e5fb75fa7e0e71153c3bd25b3c7f3d38880ba5fc316fe63894fc57b8e74290455c6d46439e721424f41b2674ca67f6f0647f7212fb0fffdc8e33f6aa5141971b0b155eec3893285e703f6bd429d25efd50be381f32af0a10355198b70bf7f111bcf557fb1a3d011fa3aca8a751b5984ee6d184c4f792ce28db36490bdd2993bc4e0732c3c7de49b0751586db68ea77aaf6e08b7f5578ca1210970b732781f9b6b3d21cd1f815d7184b96d40f545df6ed7de7bf62acaaa5bc611501a0f29266d5eb2d05ee39cf481cb9f2eb4ac36a8a8df7cff4693561f849da0d1c2d535fab2c96a7584e901fd388d310df419aa13744d785a8d630ab477ad0f949e55eb7e8e713e22cde9256301d39ed2b3b84f93d0a629802548861178fb6d0cbe004ce261246f526cfbf72234bca6af099d1371926eac0382f27978d2a00e2481f829830e3e5b2be0858c5d1bc3b7f6c92a276b4ea9b267d8789bec3088285fdc17ee3b449d7cac6916b20074ed82d125032f51619358f1015a5a52c08090c460f17cb8580881c261e5198e6328fa6db440594e0525f0223312a99c12e574e478df2581c74c8c5f1e510f684aa99c051d8bd38b2da1885d326ce23bb321abb6da08602e72a84013f0dec9b52dd6c3730a651f8e0b767217879dd857a6834ba85f30d278e0574ae48453adc09e36d2afa490dd20e4363a97e18c082a46f0d75cf9a055ff011e6858cc4f34b380251382ca780ca3e9cd0783ea792ea64cdddeafee26636f2e6b137b951bb4582c1600a1e4a37807d8b5bbc5ab1badc81fcc8e3c41e2fc794fa1a31ffddb52583fd73229c851960ff368667ba7ef0b8dca255aade9f2d09854d0f7d48dd697e8d00464bfc8480b59f983a71ce59df6e1273aa6a54b77b5448c38b6acd9391795c1763cb2c8b275865f70f06c1ba8a258739596908762bc60a909e5ff2b42982891ec3bf9e9fbdbe9ce3434a936aa3edf858d684ca304a3faf5cd13c2e0e138655dae88c5956d366e0bcac9772c8090e148d5100cf07237079fa708ba6ef0a272b7a351853d67e5325afc25761fc7eedbfc5a4dbb0cb125a18609efe3dfee39a708fca249afefc14f0eaa2bf79866baaf512d45d4c8a00645046c124013857e54e151d37e3a1ef1b52d547de8e5ff703164645551ade430002c6d0a3425fecd7a4770daeeb5bda662a7a2aa87e9d4335c06a9d84574a9785f874b9bae8316d779e76fed387fee0e318c9f353abfebbbc25d4fb527ac661221fe0f14b598c5f08bc5d507061c20172a49ba1ecda5f81e1e43f7f0e8086599b546cd6c56a39bc0cffd627beb43ed3c4355f5077c777c51a59b4f360826456befccb2446fbc24b562e7ec0ff61fe1c16d9043d3c41ab3bdb3392197ffb4d0d87ebc6fe560d965f49234e85189e29a06f326361b93c86d7cd4c3d944ed0f92bc97ab0c5650f32ed87f495a338a974cb8a6ff77ab1c369b1a18ef6765b898baa0894cfc3b6ab2dfa1ec65ca23ad1b75938a5bfce52f4436f3d57c11bb3658202a31b65b9eb61c571fd64ed6924965f9c204184963e66d10b2aef068a2129eb2ef60acc7b3f838e30953e0bbfb44dcf2924206438f95270bc7e2e112041a227f6f6d930e9ea667ed8c4d3dbb5c3344a152e3d82b398d2c00bb49ab3ff85935e0859c7c13c4fed7aa8b2e93033e78af5c96d1d1d7d7a9769eb53eaa6189748df9df0f85b902271e057b9aa82b2221d5829e0c9148ea949da532e4515f7654dcbaaa09411bc753b063b4247330ebe8a4890ec9e9d9053b977fee529ada4b9acb747fbb03f6342747624a08c315b7f2e8a0ec2bcffac8dc46334b41e555f665926ba89526d0e1086edf4ee4af2dd56bc0d32bc9f980915445766c12369cd1baf089129a122a7751363a3606e9c81693071b942e54fbcdfa06e0b8747afb0bf119fb4d994ebbb43c8389039330be5ad930eaf8fa8c32217c80241e25db39221581e0160136504a6682e1c6ddecb1ecd002976753709e7b57c3bbfc2c753a2fbe8f557276e75b70292523245b29d190326b222b609035e2a3afb80bee18f6bca078fd6dc6b04d8cb9b7ee9a938b9468a98b4655adbe0f19e4dfd05d3946b23994503eaa0d7c354aa36514dabac1eb45bb87383ea29bdddb25c9e3794c9b9c6d21ef17df23d437eb665981a0ee783d3d54f149e16508ee6b6b6a540c30af7011c75041ef41975a58d040f07bb4465bbcd0857a9ac7e2d385ac09a3d61095f975a332f7cfc622bb0acd4539ec117fadb7ad69bdf489fa44dca0d0ede8411b0f4fd0aa06d2d6d1a515e3b8c7d07020faf1df7d5ad77692e4124374f26e5e3e50dbc41ebf116bd31cd6fe5b9cac0a316b1d7c3d4d02b389b76cb66598457252f9f3334e357953f9c7cb55e783fa5092d5e6680195db6a314959bd45330a14a1204184c5446249f742a788620680aec12b4cfa564a5903a52aed2edf04130d83ffd274fd4d4b8a72d83f1dabd77f9361c8adb8680f38541e3a764406e5587c5c6e7f1cbb99a14f867e8a8d1f5146aeadc496324291e6e64b65cf0ce02133546d51ffdfebf54a4a0962e2705ce4d623574b5f0c95825216edac04563758b8ab630e2d433c3de18e7c544cdb951118bbd071572b29f941ac9a19655c5bb2d9e688379ae2a355f4d522f64a2346474a87e01249f7dd05b4c4ab6bec68977f34a816f6a27f070c859e6d0dacaf16db86ff23c64f6da2a15e6deae6928bcec44e463bbd0bc769207d2b4dce216eb6c8732046576848dbc89cf57e14cdf816cca3dee0d893232058daebf926920c802485406caa94baf6ea8223c637112b4b1959d0f780b3862677d64313ec11cbede26bbe8056beaf9b6fd9fa6ac0aed2fd9831f9d65c67aefcd1f7991fe60caed199a54b8b5e6dc7e76b7da633e94c939482ba97af8d45c6965409d31335c6ef889bc1cdd688c3a13604e41f0d72787d1e1bda84dc4d3adc9c22fbfbc7334dd30fd1d81e3acf3388be7faeade4e38d3f079528b57a4466e6c3a0b0b526a25ad1b05d9fc063877ea0aecf8cf1e61849d4d7e59a85b9ce8ec4e9c0dec14d7030e16ac2498634a21d2a58100fb6edfcaa4b263c8dae66d902c8b5782deaa68659ac5200920cad2f22757469619cba8204484c504127d49f5660343a3cc37a6267f0db20a365a2bd1ae70534aac05cdc44bb0100022e5734d8bbcf5c3498d400f5b10e85b23214fb5180b1fd18b9803d2d5fba0015f9821dba62c3e5b5755d965ba83f2737cc7248750cd5a79e0e5392281b6c97590f143b346ba3981fa78d8c4ca5d3c9c0e4d35dafcfa4ce156a958c60ceb6d28524d9340db5979f0da37b459df4a282f62799936be4c1341193def539d1fb10b30030e5a04a55c5ff54b73528177fc13d463ceac957bdba7c03e4002768a365531451dd3984e9aee423a2b6547565325a1a5903bf9014c2f92b1add047856621cc784270f12984f835f5457bce1088f19fac7c5cda465a5ca870890d3a7e489321e597c64e8126ac5a7b9904634065c9c7616e06cffb7a0c89b0d3b2c61644cdaae7c696fa85206ec9b37d59f03ef727c126e9f3f82072d1a398b25815f993c33392f07b8b02ca571300bb89ae9a6b445c4d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha79eb8de78be421fc8a9accf07c7e0ffe2573dce96bb5da81994ada29850249e85a44260a8b5fdc6d7482016b77ade7c302aba8ef8d03a8e7a5d0b5d315ba780886634fd9aebd8968d0ae9851e9fb3586b5b9a05cc1525d25e37423dba797004df6ffbf8d68cfc8e9413a2e216f993cc2090b001341e57cbc6a4417362d56f8f276fab8bffb99f9a13a94f01fba01aec474ef2656dc71becb9aecbaa17adca1ae0c9687f5b742c919b7bcff0ec9107a2c57b6a95e474004f93f11302c1f0911e572439a7a0a98908ae011d5167d2404c2b60c97aecf28e4382dff0e99f393bf0470c5022fe8529d576a1daec996504d6cded3fcd05aa703b5aea91edb1a37c4abe4e4bcbfbfa2fa068f6426abaf42fccebf672b74fb6bbba55920c060bc830ce441a32c9ca9b2b82b6d5bd2a3404f12f93ef549b644489ef31b5a9c3222c8d6a5eabfbaac3edebddcba0a0a6f5df39798999c0e45352c3207c322f0abf17c6d46f5cb6823fbeee8d4810863a6aa469cf5fd64bfa9153003e87fb93885da0d4aa6876f4572df3fd1f38f481b32f33e3beabf1d0eb5e38350ad86939f2b01ceeabf00a4748efd2c55bcd94cb6dc6349d6a345c73a00ac3335d98acaab1aebbe6b1f35685e9256c06eb3ecb7dc38596e57b508a7e68a8f5d757b08b6f0dc675b732d7749ffe6a720278d004c0d64bf8292fde0b02dcc04c29f1f9ca6529211191ea4c3766a1ff1cddc884deba03ab43652b43116a18147325b8175a547f8c7f85b2ccd225fc3ea9c21d43cc1517be02fece9bddf6ed3ab627c895ff6099a7b2837a51104eceae43dc2ee3e1dd0548202819ca4ac539818b0d0c2e200af06e317f5cbe5759e54a06d8267b294ad30cd9a43a9502a801707e5893d3fe5c42f18ae535f9c123502e9c41741486eca1e6356f05cf4a7d14449d02ff8bcadcd01757138213f5e82a7d934e47208f04c9fabdca0784ef24dccd5698b47bafe6ab13b84902e5b348ce9d5aad2cd66227adbc860b0d69a2df79c2c2aee9006b38e8722cb855f904c8f9556fe765ecba1a9d712a02638fca65e8269fde8126d55a4fc456c7878362a25918bf8025d370914e92fc6b9aa81a73ebeda263264848f2e51104c9fa0248be78dea03ff48ccce59513693dcbd161a66fff5eef60c7fa410feecfbd2a88a3d3cbfab6c775b6300c92382a3ef8567df0c9e53623e9ba8c0de6fc06fa8086462248e7f1d0bdd222cb54fc599ef5ebb137a505b24e70c3df8825f528d23f21c8bc459de7e269009ed532b5e715a6308928756a2261d52447b72f0f5a56e24d8e373a44505e30c9b77ed78adf87e15010f02814961378e842b85953553a142ec223c3209883b7c9d1a23bf0fc1a49c22a8c1c70fdd6879a32bdd1a11b9ca82f0908bd4856f826b1f664a6f9c3082ec3e9930955408c8862bd671f397b5cbec90b2ef4e6b202e2d6233bdf75cf08dcaf7ca58258de9c27302f68c9a0e502216fc2d07470374dcbaa10af1a47dab9c80a367bd7b368cb1c220a64f183a1c1ccdfad1f63c76fdb518d8cb214d7cae593d9a17612f4b369cbce702661cddfa2aae6fdb721a4c176538fa7a8cfcc4e62d98f4c61e726de124ddd606a906d42999a52c129cf411098ad58f1f2f78c830ca1f2343b568c8229e236f90a2223ced3af8a80cee50b3decc34ae254b5ed2e835d421a8679a10cdca90725bc3313f0ebdf2916ef916975e551422ec7fd9d5c982732051f0b436a3824529aa298b909d1bae1fcf8cdf4e80cc8a51523a958c7d3447149d3fecd5fc576fd6e59581d1119be5e48dcdbb33f26d2167511915654ec1f479d6cb272c6c9a0aa2e855a3a1b284bbe3513608dd573aa7d8c5817f3075d15cf8067ca4332c04787944fb3a18e9b7351fd8abc088dc7286fbb10bd1cc071669d144c0f9867fb186a9467affa05de86971f172e18cc4c741464564fffa2442b9953c45d89ef13bcacb91b4bb9d8aeb274fa174131594dd48dcef2d0202608dd9817b3182399f2a7edbac3dc91aede9884e07e40ffb773b34c95597567dcf292db9f3f3905fe7b2c2baa8ae315a7a88aef6498de4c5854af77362807bd2f5125405a79a329b812671965fcd08ed060b743e898aa3d7492b8432dfc827d0aebd5eb4ae287809d0ef3aa18e4ca262720b48a723afd8b602db606e3bcdc9d6015f6cc7e0c580648054ced8615c2500e12ea7474a1061f05ed332c46711c443b0a6e203e226f71a9003302bbba56e70e01f25e57501e2fafb65de7b793111a3a42df4636719823b8a703f589731a317e35423a467be1b33d4255c61f63c0c7f8a3d5ad12e78eae8a4fd1d4c5799f5f95d1cab284890e3ae5c70fce1000c07dc0a8d2a71bdf59301fed2ba5ba95f8461ccbcdea58eb7bef5c40610d2ef6c018d66ba4aa70d5b0f2534d37c685f7a10ccae7fcf35e5fe168c7947a73889166d1de1c8a910e4011674ef8c82b8f73b6d67b35d59040ba58a7ff7de54c338c262a92b2190fa2f244023b412cde790ef392d5c6518e8c5e879d582153dd737d10555145b73ea0611f8993f342871f606a0bdc5b7e1b5db8805af56d94a2bbdabb407549819fafc9a3fa07312455a359a100305344ba6e8bdf46a7066c423e586e307f7589c13930ddb8c63ff23871a7b82ba08af3cbf642c50878d1400e076957cc5865f5f69c915686b9e02f56df9cab5d054549bd810da86199a7d328a6635465d58e3ce593e2f1bf393591ac0d610e05a1bbb442324c8a3dfd6b5ce5099c6d46a966d16d03f1952571f4ef67791ac6d7668511d00cd7eae00bc55eb850c8ba8ac4a4880d71873c701015763da430354d29eb2a6ef046841c71e0d6d2061e8cae696ef04cbd75aa6747505ab4466ac8ab99f20d00c62d2f91f18b255c06a6df7628b5d3770f77fa125c014f5d9a1680aa42980202b5b72a26f035c79d1a45a0ded6bbba35f4db10a7afb6541e04ca2cea786e329e1f19d563e725eb802952faf3c08ffd48ff6c45b5540388e6c98a49bc18cd121ddb8a4234a6cab102ed4477b28cc08d22b88e8cc68d24143c1b73136bb4b554e316f66ad61326da14461db148ead21836f18bdb5dbfea386c3a1e2c821db1497b90f2051f7525a9b19a8a5d708176fc1e510d727ff042719ce472fa1a2fbd6c8cd2b969ee772fbb7339dfc843d6f4768703f749eb17cdfa1ba7ea6311a81feab29ad8e96ef5b30ba3c7736d4f7038e08a06a57f19c6d28025456ef5d9af9ad997476ef2cab760d3efed31cdff08819703fc758b9f7704ab61653a466af8db498b45a6e6f17cb0d90de2ca006e3ec6d315c89c47a16d930ed4d51c69f16a24ca43494ccf3eda3082ef6f1cecbdc0b4998803a1ff86be91cc225d41adfc76b6de9aa8825b57fa67b0d408b6f5cbd96e896b9bb7c1b396eb39f05dc4af30dd155fa9d0324bd28682d951ff64ccd12b3e2f46559ba9a6168d54c1ca26a2fcec5b5bde457620a377390a87640a2af128b9cafeaa7c29867005646966e25ae2c1897c6a7b6ac2a4983945f354b2b52484427eecf058031c98cef3a0ca84d3dcca031ec7f815f189703cefa529c20e3f7ffe5522dc1825e541de67cd4f3ef3a0b1b89a79dc21829d87bf0d6bcb84244638c07532308f5db875521b489affa43fa50213c8b43d9116bc03d3a1fb39fab4d0daadf670cbe98a8b469993b75c249eeb33c5e822cfdb3a9695c171fb3ce1a9ee703445d71ec6c9d5d97b3313100998d525d30b86964c15d993348ce6f3521abc7be32facf25fb139e6a6e4afab125a900628589aef851eb192d31f905e6e1317382885595487a602ed683f2539f967edf1befa96d625da12566a581b481a42f017d6aa8c98fff2be99d34afa717f6c16d5b787480d59d49fe21eb7d2492ea1947fdb87cdd84521658c8550e04d5a40021da1b77e0a7ae6a163d027f539c75ab9eb28098ec2b6ee354fda7321c9743259b965076a5b91cd1295b673ab488ad47a75ea700a708ed353a4ae9e1efa6eeaa1a97ad5d4a2e9ee6064277f10d40e804ed4787a66004d10379fdb69e17fe48e10cc85f7387a308b5def7b26fca5f9fe683fbc1b65b0995a4978ef5b79c5ef7c44b02d66a22eb116be57280b91b686866399d6bf175b18ad82a9428049e40bdc77c348937d74b9ed3d15afea2558a196349b04f2e4c32df135250f3debdd09254a2981f308c38a3264f52b2335cc37973ab76855f02b46a6aa459910621d8363ede9995460e93c81d9708fdc4b908061e1b3a7f6e97911c9bb19930fcac01b4ea5c1728e5221d43365a3257a651c85825ca2650cf775f9d790eadb99f623d6151aac0faa0efe07c1205832efc72240d1aa96a80cbd73d2b4210d32d8425db0a2ce2d6e956d912ded84877ae0f2aa3dc1630021e6d0e9ef9e9abb002cd31341259fbf6817471dea0cf78300c36f089ef7e16534cd252fcff42da7b85a4894a7b27bf0f0c94f64479d8e358470bfb39c1303cefe88cef375c9a12816ef6be5fae51342305d3728931f7ac7fcb9d9c94c21269bc391f55bae70e4d868db8fc2d1584eccb4238e858a44245a89571cb3c9cd2f82a03bcae2e0a62d5513f98b674f8ee2ea7fc31fa3fea8237ae67b98a912d18f102da03718ca144e910324932ad6c2a36ddfd322c93ba8cbc53879da12472259ff7722060d90061146715b5299eea252e33a089cd020c63d3004af2ff896ee020ba98c52a1df48eb4416fa53c350496e6780e52a611136490b6e11f8dcf0529681ec08505e6425b92741131ff734aa0733a86e2d6fc57c6bc76f78d29ed026674b36ee02d88794e33c16b267c35a86129b8f18344fc686595fbb9fe08c5412250a41ad5dd4e48024e00289f2cebd0afac074e7012d4507638ac053aaba5defbc4bf5ab90bc76eb0629c76496fec71dba34569c350b1bc6361aab45b84e78aa80d1c4ee143eb6e8993bad90564aaef83352730ead999cc02c101be4c224f5685e729422dfb61a31646c9b4af8dc42e66d3be4c39bd5c0c17e6905cd254784ffb33ec80902a11e746af757bd1fc9402dd00405d5e161bf0b0ed05b1c2560f296c82c1410184c39dea160c64064d42b73697b328bcab33e51fadbb68b61feed7982134cb604a0490093f487560f00b8f3c534bda9e85cc9db1e0473c623ed5564f2d9bd458baa69b4575ac82660a3ff0535e8ca8ad5d0e5882e407c5f19a4a391f01048317b21af093e888c19820d54a1c3bf50e0f02bc35bfcad3bffb02dfa68f20092ffeedd7c19bd24b16da95d83c888f31adc85888112fae18951c906b2fa1a6f2d0aecf9a723f558d53ce4598d4a9aeff1a260297f502b1d3d24123bc68ebbe119e8ccb952edc462a9dd51c43961ec0519fd6351b896830a41af60d07722e79e23d8d271194ce697d9191cf46b31c1dbe3680ebf8613619400fd24b163eea1732f779405797b9b0d1f8edc2c13a15e4a7c0b0da0303ad322fa4508ca0d8295e5c0436005912be2554f4c69f4fe8628004c333c97a2bc64f8a080282e1db9630e1ee839d7f1a5e8f1128d664fce51ad302388c2007403b60075a7df1404cba45a75a1542e485ebeb3c63976a8677481e56e00a1caa4e3891ab00c275eb2ff7b8d321a4987e33f5a3e4bd55627ae600e78cf7becbd7f66213c307893cee8704444f9ccc756f4e10cf8aab8ee17a6a5a20d60148a3e95f09d5ddf987e146236017bdd546717d4283167f7ab0909643b56666288ef81d96ca8d7419cee61eed654c95f59f72ce5caf97c885201a922b215863e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h885d436b9a8b88e11385889f7bde56add81882b070da313afe3bb750a4af7d3fb0e751654dab38b892a9638f9779da8281ae14d11f8f060a640745a3a188cac474de8d1d8d87d38fa6e7c071f86c86cf56364c9b1fbb329b9a65461677d46faeb26eff07309adb74d931239cb3cfca877a3c81ba9ced0e543dc0d83a9cfdf9a4b7e45058d1b192b310439f20293263177bdd1f8f6077a351d923cbd2378039286371142c649d2c0d3c732b854805079021b655f8e7df22983f74e7299b6b7c5b59de494ae543ea1d977358700f6052b221a3a46ee9a41e8989429bb2583d2de40d51a67bc949b819e694db18fd4ae4ff39f53b9c711388aeaa33f784e9629f7bcebac5ec56af74c6e1b9fcdec9b66d5e7a9af798fca8c6ebc93c65696dd25c78090f3c45b6f59f5ed3796c07f856186b098d568ea1ac36a16448c8bbca6ea917fd8b4c406ec2f28c9684065836372307ec87485e637273b2b27aec2c1c2ae87e0cccdd79258954accaf1d1a58b811214df52367a520e7ccc2bb3a59b1b9a311e69bd8671b6bc955a434c63b071cd3167a4e7426f0f09058313b42493e5731cdf7a3333b1f691d1230c7c3394d83b88d44b3830dea306401b0948698b56043e93853e00f1a78a3fd9ef932e0036665ea5bd2d6929e85c0212147fc8c187c4f881f3f6f2afa5ebc03e6cadb49985b8ff12eb58e84d71c061c210ea4d7e6dd500753d70b0b01bd09df27b3c8fa55d4cff01abb89b45335383f20893b5417d1c53e9e4afa6337c1d548c08a2cd4409b5cddc7c33049b3ab84d46bed065ff7f68d3ea3c0ba33ae14a9d6007a8d288f7d80a806cb0e1190a1090a8b8ad3d2346da73aaee981d86704ee0e9fbcb55f51fa997c6b916629107bc06312a70c17fd86ada3212a6477fd0dfb3d5ffce096c576bf1150e26673f197ef24f17d8677ac5f66a8c9dcd1f0247c8f3206f432a9ce6629e0c72695e92df87194e7e6c631d637be03f314d8b5e3f7bede6e9013b0d5b50b855a41dca68cad815edb17baa0f0471fcd62a4e4feffdc2d44eb4c8280fdb28c0994272b08b3052254b5c4e5af515c6a67ed95754feedd0e6fce65825d2944695edf74d1be56efcd32de2a4997c4721c1a3677a7dd6374469dd9b28cd2276241dd234a1ecd15e67a3255d5b2469c289e295220e827a8fcdb259d6961ec779e25e753903818692e620ea50a64ee66a57e5bddb3fd2dfcaa1ba9bbcc460c5ad5de780c42336b474f82d522a65456c917c7e6ee28383094aa8339e835deed81d704b4cf6e98e4dddf1820da8ffabbed453212d0f0aac8dcb2a1bf13b3a829ed3c013952c48a6d6da221bdfcd27b3b5dbe80245ff27ba4340951c0834e9a1dcdbcd880e9bfdfdf57531841ab1a979606a200bc2c0941b1c3ad67363983cdeed4a68c4fbdadbf310a86318028c24511f7d34797678d18bb8f96d513299ef3fbe6ff7d332d8ba75fc086023a9067b459f1fe3d56a420aac809f6e60ee5c710697aa48833b4f975017a32038c7d44d6ff057d1a11fe542c62e484edde7b123492e4dfe1e2e5c3b35ab0cca856e073841ad4e5839a5390c7607122951a4b31ddc493f5a8f9eebdb44b56d133589c464a818831ec1816d324ed4ef4cf16a3eb3c5376a1b70a6bc960eda39c487c9c768604f25cecbf93fd7b8b94fab4bd8d6e165edad16bd38623a76533ce6bee4cc1d45376d2352f217a6649e03ed33b188c4c633f151f20fb9a931d941eed69df151f8e6cc77519641678ec5a12394837985720ea83570acb7b2e2fd8aa13235f1effa29c50a1fdde7f1e80122a64a92d0edd03008e0a619745f0b5958aca84ce4a2d350259646e734b907c2cfc5dccf85ddf0cbf432e79e376f2e4ddbc29ef0a7db20d4eb1d5be121332814b06dd84e4f0233ea2e3fb12f449cbe45183282ed17c9a0b2c8e4f327b5998cda5a94ab51e84a5e1cf1ed9b74f0f1ef32d7adabf903620acfa227477bba18581c7fd362a417d5a03aca4e87d1ec0484d2caa3fb7832433c982695bc75ac968d89dbc4abf8f058bd94b08dc6d7f885bce38127798bcebe6f67541dfd79b1c04af62b491bb96635912146cbf6eb94c448b70970ed91562309f1d259b970c3557207d4fb5e79ce9541456017b657cd45cb37fab730772f2a76aa75007161d16f619dc03deb46eed1561a1445af1273aecb345ed8f696242dd235ac5981f386cb10f312acfda7d1bda70b9ee6d326dc35c7be848c389ef1cb61fbc06de12510c7ef55f188f80ca280da4dff21573be2a3badc9568de56f7c312347f0ccb3dd0ae9d38d7a754a6e92b8cb46bf780143e19caf65e9d121dbdb801ae30c596b8a428d75419f01bc8fd020b1df1dbac4786155a497ff0847a62a47ec743f1be5414580c2f39d21051bd5bb4687d04405827e94005d7882ac6868938b6ff911c71cbbfbf9a3186639212f573c679d0cac99cfd53fb9564f54aebb5d8946f61245926ef3299749d8174b4b7b8e60b0c140da18de45940516575cd3edc6478237ee3f42f0f24b9a0491a2c12d69a7ae8a3757558ca64ae2003eace7e8c2c6a5f809213d68177c7ddf4bc672a3b03be44fc4220b7131ac5bf90de3798c4336cffbd2f0e4bf9660fb8ba41f696b7e3f42a0887bebc14fcbe7e83d778b8f7c37871281c01b545a42fbb1cc7f95a266350edb8218292bb4df17f9517cb5973487435dda4230833bab4d093d5834e218eb16b3a991087b2de299a5003ecd5a3cd2ee05a02900b08156f1a7b75fd5e81e2d4ea1b52c5bb0cfad3016de3c8b400350e54a71cf53f547a0a9530c93a2b1779932181f8ff2c6ab91da15e24eecb90d60164f0d155075b80c495c08807dbb63224faaee65e3c0d470384743142475fe3f5bb9d45c261ab42402fcb09067df0c18d11966989ff94a12aa85104ff75bae16d87d5e3a530eb99c36961a66683a324060baae4a561f283bd06cd62d76b7c8e8fb4388cc00c8c820c5d951a8d139a95845c0ca401090a21fd087c728c21e6198afed6cec7586d19f15cc06d23a83970cd53d43fde1a6aa5f780f5092ac6e32f1c7f64572165dcc8cb73f1c4e5b762ff72d96a9cbb5a5a4d37bef969c86e8fdbbd76bf85ce8328483abf132e00795b85bc60776c1d08c883fa8c894e24aa7daa13ce61af87496d18895080d0d623ab3d7094bb271fae312f75761062149354c610eb2f4101ac4b92cbb28046720c0abff1666199b5d26a4dabe6d4b237809ac28d3520185c97d8f8f8905f0aaa9e75a0aebfcbce92ddc969a8a11a7898c7bee0bec07d79f567fd87dde63329e451966fffe7dc8c17c69ef7ce59a9e6d94c23f9fdbecaedb55e4cc6ec33dd4a7205b34f42c15bd6341d09b69a043a8a3afc44283bc9f52ffe69dbecf5494866c598e617f369fe7015ab29285f64cb39b04276f8a4233e8a46b8784dfd2b41e189b17d84be76ab40cbe79855315623dfa661ad79aa76ecbab89d0895f49315ab3de4f27bd99d62dea594a14106292a2153ee75f6896210018cd0a8dd6f56e24a082aa92e3ade273bb673ea9beb747b04ac7bdb17bdc22202696667663dc3ca0646d84e77d00cb588222080dcf8fa94200f86dfe052801a8f6273cc47d2c24f0ddb46547e7020d4b027567dcc3c598fb7f9fa711f5e7306758fc2f6998b79c4d86726301e996fde47fb38471b79b9cd280b7fd6e2a85d2acb7baf5df1ad003cd05ae8160e1f334a184847351f34c230fc1f148ec2597ce6fe86db7715ec67a326b586c185ee06f0efea78002ee6e714aa4b260e861a0ccada0a8d09734a5315f5687cb10d9cd4f9cddf442e99d948445898c1517b0e17c958d5bab6ec9c1bcfe69e500acc6d41919f1ae6954e357a133cc29a57d6dd056d85bc303ca931b29e7cfe4de3cc763f99758736b5d706cd6c0907499573ac9d80d19985a49c54a8a4b0f23fb500389ae70978acd8d0c14ef586d289222cedeadb1a163de391673f4870a4f1c5cdb1579cae9aaa5cdcf34a3d2085d1bcc341797209b61e302afa8159a82b4c268c72f390cd998de7073bf4fff72acabd479af38ed1832d463cb9d5b4fc8fc7c529c196a94cd1b804b5971098d61cb754d206b9c5716169177896547c90a7e9be0ace1887ea64280a8fa3b4fce6baf7635fcafa7d103e36c72cbc938c2edcd0c0df48db64cea2472262a7e8e32fc4d052db432d78e3bfad72ed2e30c84d766f5e4d43f0e03d914b79904ff108c76beb2c64adc5f7bfebbb41d6316007ad4eb69a0afc77aff8f55387532f8237b93226dd43586c1542e70a01c26fb6ff23573ca92e4ea19dfbb76d6e951e32914df7054fea93f7302c21aa4a1120ad39662758d449ef93e4d0ec85605c01023b5fc582e898b5ea2c8d11b9f6c48c50b1ae46c8e0b81e6b546316fab98ea0d4a361a782cbff8ad0c30db57e3425fd00c8acf69f50d70e394c28f81806b7dab981ae8fa0c050424d63ce4a6ad758d47e15fdf0ef510171bc6b10975be5c147b588bc26fa15a675445b3f1b3bed450573345f90f7e7360fd67d5636e559a84a83c61d7403d8fa14f7ab968bcc346f589f773af8a39c8f9540caed50d65824346effbf648f6506aec03716d8bf3a2650b0ba3a1474592a2a67812478c7b6e66c899443b0646b32461cf6a5831b6b33e1ce7a799123be443c2de3523f0c35d0a2f259248ec121a9afb8d766a55b898afbe25a882b785d257567bed71f01eb31a92f3ff23872b8dadabe6a00b0374e8d429a748c09babd17b101527cc76cf6dc85287344dda070a432270156ce70be023d432a0bb9afeaac725ebd73a04b59669d4e6446b786b0801aa4679162e11732fcbe056c2cd566d4607edfb73af2e168fd6bfd6eeae25dd8ca1eb21b467805e37960b504dbfe885ec633e119d824f7a5f5017915cb2adbb5e2c2f6649584310c8a7f4859125e33fb1ab1e4a190c45474d898bf5a7d82b32df01c920bae870a0c0f0d47117f860c0edc1f18457cd0a6f932e4f75c8d7b3b03bc8f61f7240addc1f2ec05eb778e7813c97d07a9be40e7e43a5ed4895d8d55d25088ea3fb120f857663e4bdb2b789426edd455bd92e0cf91d1259d54af81638fcba51550f08b227c41ce21dc5086d3c70a6eb558a753d07bc204378731da3446e9b7ca073b2776145b00e6380802a72b6f7c5f36f18320a9a329238a9643bc9fe01549427dbe122fe15a4d280533169f2f2458b17f6b3ef0626d61603b38660be3b061647564c68ac6ef4d5ef7be617ba4cd3cb75556eb9553c18ef3828974930bda82181f0f2c1358cabe2df7fe831334c4ef117b36fd47d862768c1682663b09a71ec7c57b9f8cdddd7cffb3dc7e35daf2ca0220a548b60374f5bd1eb1d58d42594e342983530c3db1715c84476fb4894865477b7d1d4b9135d1804b7c9d6b25555d60f6a0ca189ceb8f8276dcea206f378aff1b92e3464afcd76b64d795f01270e7776486c6a8ff7ea946f9d194bc04b01908a7aac1f53148632022c218dbb562183c2753a2c8c394634903432b6424b3c9997cc607ac60d54b1714461bc60f6ad168f98eb9fc2850cf71edf99f4399028841bef7ef0895c2b97f86c37d420191d8b7e155aa7340527949b2f2de338ad1d58362ec344c2a281110911082ebe43541fd40641f92a6c775b15491465032b9336697a6529b062b2e8e42295d0b8efd1a08ade3ca20920e804aad2e940e63acc31b026a7e2c152ab03b9f0b889ef8c40dc1564cdf42b62074846347a1f5ccb15c79a6f95d1619ea3fc48af0cc88352f601a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h21b2abdbbed349a0266d269fd272e0bcf6040796cea24cb7f2fc2f43342287d4609e64a3c2642a368b22a32bfc8724c6f769bc66d4398789e2f2f3454da59369033c77b3635e9cb3040ab9985a9921eef9677adf5ef638ebfbf745a0a9dc82a7c4bc5aaa4d44be5569c12700c2bf3ae85397388ed9071f6ca8989df84370ab1d48ea6c6f8f54df9f7be962e3c1306f139c854dd31302d0286ead51c29d3109af152918e9baada042efec003e577b9991630113cf256f213283f48dcb6ddbc1b4a79b32e3fd131681e83dc476f2365e63d145e4c40ffa70792631159ebefc6bd88a14368721307c32387e59ccddc468c3a6cbc79ef9acb1b55a660180fe5117d3f45e350060d4454c02d531fa4647184a4c3f22059b8c6a6e39375bdaaf8da4dabfcd803d0daf703d0d76b30d8f1d717fb63d552f41852ea265cded041972527195a56ffc0fa4949fa5ed423b9bce3fc024876a37daa4474c6d6650c7a29df3d75179b57acb4e0a6d28cf9d2b18b138fafc9ef390e53e3cc05969c830dffde3643e2f1bf598d684a42910cafadae873b83cdcda49a7b9dae947aa92fa52891ee23d28af7629cf0d4f2229dd136fa2525cef3da1763fc8b1b8681679163f50af2f689d349e675dba8a9259d1028a0cbef1abb35c04ebf2a5834cafd1133ebe0ebb331329decfbf6236b9d236ce0d656280c8dc7da27ec7ec292f4e6521ef58b2508d3d4021ea4ca76a013dbbd052a231329a69491327eb1cd190e831854016a58da5d7f6e576d33ff7d04cd8c48eb94f1312307f2ce35249cd5e1b25ecc85d6f47fc53e9a36ae2c768fcff011f7afbb73356184dde8afc4b55e0eed57d4ddf67b9eaf04afa629884e70806f9724f5c8ab1c5d063b4b4dfdeb8983d76b380ec0daa88a0e910a9548f826c81a17ea91c3c01296a2e8eb47c8a7e0bf520aef7557440ef29b930359beebb34913f42861d4e36af1637c8987b7f0820028f6183030744a50a5578f5eb3dac99c19bef7f2ae35f85bd8772bff072f02da5a8e3d0e6cecac3927f093d31723bcc395813fa74aade4eccc0de92ceed3453902ccf4495951ad60a556cfe093d8b7a1a2ca6ebe6eaa6b7aa67721bef6d998041aac8638c043e7aa43bc43314720bb1fa928bad89bd6378902a393d262604036bde6cefb43d53fdf6956c81e2b312cfc4ab6c7c50efbb84a9f2b8d672f1c7bcd561a80105459cc7c5da2d650d84bff6393ae1c332e181915a6f2728d5e093ba6ea9bcc32341f6a254fc4673802f538f49a7c76b7b86aef6e6922a3537d324500dfc06acba87d5f9d443bc8f24d8601ef73e03a5941c593cdc479970cae573665044953e8a14e4b4724aa1c9f866524a209feae4171701d3e89bb43afbcc3ad5524fc6a57b27157fbc0768e07ad8642e8a9298e62aaf617c5b19fecba324ff392dd784135fc4118972daf094d767a1301953f3c8d6416fd97c2f6c25b24e9300eb2ffde7f30a3779607f9cbc171678f9456a1974ffbeccab1b404c7d5b0e57371fd93425a48e622b5892b6c386c75747dbad4ea0c092b0b07b4fd2c29a2d2df1a47f9f46ff6fbc33cb90e9c5cf1401fa55fd7ee1814f99468b48158e01711fe56a0192f2a0b38887563c5b33b7c2da80d35357435e25f4b017f6720feed41e40494799790787530ed46c77425d551289e38c83b588932435358655a8a866ee98a51d6f0d0af1f61e96401fcbeba002c15ee2d66e52e26b7d98731ba67a60ae2ada11aa37f2e6443853cd80ffd9aa0379886c4e0c65de5b37b439b95a385c78e34ce6b69720b76d264f53998a5e3f6e929a4bcc2b549a09a564f83f46569cf0fc9541f606020ea8651d90b2e7a733d1998563a2f88aad4bd8cdddd10344dcb6918a8b56da85516449940d495b23fc2bd4a0584cee36851ece44d343c2268e8a91696222df222531596de57fba8a3508bba533d2bc9956e7298ca18fa6332dfb2643ccfa3d81f6b0b901f599eddf682e3286d7bdd50b9b6aebba4f482acb258377bd8d01bdd6e5b0359879b98dc57283874ae208704c5d77a3576a30ac47962a5fec64a6300b0942a2c646e0e336d4204c16c9cc97f948a2774505884410fd135991ce8c64edb9641c8311d3543a90f5ec3f02af50478bee697895a5bf93384029a83b9337f2676421342e8cf2c71437f973fdb9f108c6e766bf64f4ff6fe8b99906f5d91bbefebefd475ed469ee51a9f0f270494d7c1522f83bc5615966006a2a0f65d1194ef08c14e4ed777992bec245541e9dd90f27c1f31302828df996b11c9a7b55c3eaf90be2fea3c717844e82462ae6befbb029db467b5d191296322bb915bd66a7adf81ba1dd6b47cda08f6be0cfd1e7d0bfaddc1230d20fe3249588dda3b54efc32d4dc7484a2b996601f5491172f9bf67efb1a21cb2b0f8f6db7ddc94c374093095bcab9a683a28e1124471be2f937cc35d3f60d9c293d12c7df42573c9dd05057b601604125c19ebd050a6bed35a28031dc1ecf2e3a88bcf240dde0bd2961149326770106e4c38fff716d9bba21813f8e7b71d80192c8e0a6cd8509b728c24320d3c3475e2e09a787569e98152e04d46d724283581c4353c2444777a8dd4575276a23e9aa3dc7c1c2487dc2b7de654d612e99edc657990384a726a58719812bfbb874d2db0d742fd041e36df54976de52e8070a54e954013d02e588da82542d7071c7510dbdef3450c458cda1bf7e2a17aabce7977dd4d99054f75198bb4fc616337a9afef6243263b457f01c44a124a5cc3b3bea8b83002f0de2c0399c6f3e26b4ff0a78501856d8a139067c4bdd63348fd7e14b74d03cf535ad895fba465dba8edbaf58f601e910f69b5ecdf37e19f389995d0f30cca3e5b7c61c96b0acb861cbce2f9a359ed7125b16d77f8bdae416cc892097073a63d908598941320f31a609f52ee11bac5d1722894ffac564a1d91848f0b3768c04c12832d184041c9500f81ca703d93b7f4f699c3cf041f0d2f0e48697819c1b574af92194b0b9df7edac3b807d53c1873e8e4fdaf10e394eaff1203d56a81a6479520dfdcb7d38b6a126bbfd7ecd972f1984aae49b84d9bb713bff99876dbe1de4dd9b2861b3d7663195ef679b62cbd2b4cf32d789b57c4662aabb886ded604d4bca0fa31991be4bfe2afbc7e842a44b40bf8815f40c9a5ccd5c528aa91eeeb67d948501b2d97590543c430ade43ed0be6e8a19e2a0cff2358827546895c3f98ce12e6a5694c69f766666dafef18196f504ae1d20b4db450092f1dab63b230c5e25f70b1a820a37f814d6c2e74f240fee555e238aec956518994baad5e9f22160db32cfca4bb4762c37dbd83525755cfe1f6038bf45478b5cd3de8f9cdc2ffd3892026d653012b98683a36750062ca46110fc0b3f8052f31adfd8cd434e5bb05837cc23f89c0007ee0dd4921906f7548db5d13d310025da3c383b20d6505c6c7fdd742c3d1b044ac51a62bc241bc8ceed901a39522122c92769319b22028034a08cdc7ffdfcf5b33ba630ccdb08b6496170a90f0858bb6f004affe00837868d40dc9299936f829e32519e181cba31364c51f03867ce14155ed27160d77c0df26f45b6839368ff2ee5669858ff086951534f20ea04d70867451c56a8078b7ce8ddbb00e6fa465d287ee2f7d86fe4def23da5cb9151edf32a8d45faec876d1032c8ac5865652502553f7046884c12d9c15684226087e6c171d9bdd75414936fb89490d0a59666915afdda429d47f81944b8b1e8eeb8df9e0ac5d3a802bfaa5c919ed8d399220a84115d0c87d6a046bc5710b3911f240c999d358690dbd202abde4b3ae07d0fc0cdf08645f4a7901a2c5388b8e991b332a3da5c695497cbc957b398424721d0195064d2e2cff4e0a0256a3c10c2dd6603e52dc51833074bda873f35e4ff6ad803f4c273242de48edb40964354e9c1f318afd9ffb8f9f516ceb6d21e044aa061138693960810f3cdd617b271625919f7456b51a9a1e8ea50fd63ded8979828a9096b0b712d36d722fac20839de350a3093dfbe4a4cbcbf1c28f91bb325f94ac32a54859d617c10aded4c99c58df9afa6ef9fb9c88dd5d63854e94b8cedf0d5bb50635d29c0adb60dfdc8b379d35e0eaea2e74d20fd20548b67f2edba61fcc498a42fdbda634555e0a4fedf3a26d8726c492fca6aba4053791886e98735c06ef59b974e432b2908a6c35d7367dae0adc1ffabf91fe938686454dbb79a8d0e47ed385ed68f44aa1f2be71bf173d0f54ddaf49c3958ea8f78b488ee45a95c70772f37b5f332f063c0db91771cbf009f5308d27d51a96184d8be5102b510fa7882aad2257809f575a5df67fc103779a9f7f61e9ee879b6ef6a05a16c7be67ebbd28f7939762cf1c7c2f1691b82d021fe5446aed323c8e503babfc0057aed884b5ed9806a0b072a235220c32adc8bb9f8e090ef2e501909be1813c89be6283358090c6d5bcb005d48ea148827512c5491e10808c3eaf5b17b036a4f2a58256a4615e412a9cc44fccae5f08c128af3aebfb55400468146e00e860fe11de01c48d6bd422dd956ef50999b52ea37c3e245511c705a93ff63c04ecaafdeadedaf40713d036389f0d110c71f8cfcca17a821d4172a4a6ef327588b71deccdf00ab80d8c6f4b901d40c92d7922ecf22b7272b1c590b25e577ee56fe779a46fcba3132ac25976b85fc3dc11a67637338df3825c83dd95b14d1eaaf0bc3135124e83801d68f9b4832e43ddda0c3203e602e2a4dc91b47c7517c3795dda8aecd242faf514187702a22609895f50b81c9cfbd0f8d2111d38e99ea63e840c834b44f576d45f4f2398fc628e6095f197d20c27f224d9a0d00292b463952f07378faa31a4cba4b559b089f93dc58c36c644369c6d9f6e332ed5006f1fba0d61ab93f4bc512c137433e65e49de54877647e390870561330fbbb9283419a641ef82c6767bb8daf513306b54a882e47ba08b4a62112fcb656eccd1f98a46715bdcf0b517e2f9392cb5852b510a13cab9558f0a556e49dea066630c080b049f4234edf6ca2efc732b18d7cfed7750ed1dd79cfce858ab07e200625accc75f19f88ff8b3e63ef8b4ffcd3e9aadd23860a46dc778d199b485b7820cabbb28fd5148c582be5521f36a5e153483aa397cee5237d0595d01364831f0140189b133ee263e2538408baef4a6c59832ffe4bc008ce7c2cf407597bfc43af11c3ca4e7237b16b339134da17011e47cc8618627e45305362670e8e227df571c6e1a987724e3d0ef0df46ba9390719e97ab63162b5fdd1cc541723f6d874ff9ee489a7f7bfad5b34da49f262d8d5a0bd2157dcc0eb99338f3ec6e4a2d3b886a46b208326e1b3526a1d7d791da916add6c89c51eace45ce989568bc179da6dd2d6bfbdf0041ed6c1c0cdb03c618eecf810446494418c51ed8d05bf046aabe363308b923cb520753c455846caccf375bf58f50ef2110f3744f239b9714ebcf3104d8ad5af8b12c353fb410aefe091d404d79173c75907839f0fd778cfc03c95415e1981af8b01d9db4aaaa516e3e3d3f192209ef555cfb4a1c22adc1484fd61f475b181cfdb434144458209289c1ced1ca2bdf2b4ad62f6e38ffaab459be44aea87daed9fadfddefefb1604aafee8544189520b36c794b288108e98b80d5dd72706ba907aedc3e854b864f030ca7e3547cfe1f4b2bf9a190a1ad896ad31331d1dcb3882574d638e19d0d858cfab170f22f98da3d7ef285be071459bc6ac7ada69ce2b799c803639ba1277a9541b82a83c2b640671af6244;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h309d08507ded6bdbddec9229ed37950b4c77af80e1407bec63b84c5245ec80f37766a80bddab69551bc25a10d4e34ffb9850f1eadfcdec8673e7f090b063cf20881209aabd0c7fd04ef1b5550861612288e4f9b6f97a9ec2e47cfdc424b15bf277c560c899a42c62160085ba1dc4a7df214a4e6297eb58fc5905df923906c0ef1f0b813f6e18268de88e59b790a02785b6f8d7c8f7116bd4f1e50404dbb3e8520f67df70955d1ef18bd21a87f1bec7211b8886651282156790752bce89f4f4cef73596734043778c253d6deddf05119607e513c32970293ecadc5e14bd83da1e806f4b8cb267e935684ba6f25cfa0ddc7140fd9c350220e73a1cc83b0d6b79f9017c23d64639e3c3402dae3f2d4d42531ea2ce8650de8030f9d412049019a14325bf9eaaed8a186642bd517d258883b06db95e42368e3a2a499284409613cb50d71dbed82415e0f2d1e6d1582943cf52342b5cd0d856347795b55aabc911b79d1f219535327728444071148a53e3de304c723208ba372b0eb0d9f3ce153396c3284a41deb063c7e137268e8391ea7377bd28fa00b6e71d54ea12e1a1141d00ebaa72a403099d39c5615c6d8782d5d32f87081f68469b33dccda30e2a5043e76f6e6b2871fbe932496eee04a191d8adcf6450763bafd36194002ab80e5fbf54ee646ed64996c6c7ae08e7d9c95cb32ddc5c21c321b285457d4db49e2dbf8e6d670af001307a613dca716373a574ee2aca3f497ed804f93341929dfe70d84c5b870f95a55e02fb8dca4cef5e1d1bf19be1a30b54adde45b89a14c36a5b8d144d50af7d427d1a2be31c421f7641b0d175b8c8a8484ecb58d512482af676cdd6be1e71db05c7fb7f45a2df9f27a61940e07cc0b9b77fd64657a43514c9dec67527ccd6dd433b2fea477254064dd7efb5c596ba2afe212fdc408e6c1b54048aadaf88c068efe81593b2ce643565fcccc5908201f2a796bcfa59a0bd3f162bf123410b15bda90881de0774cad4e21c39fcb79e4c2d17c6115e40f9fac1359a723f777d488ffb7c9301c227a15f355b90f6013680a11fb5756fcbe8554b619da4aa2659dc031eb607ce9892cbc0095af706014516b1c12d952756f680ba96826f3d5a8f4b120821b15c568151179d8b5f1bc8286390293150fac1c18f17d54694a9c35ff7de8035cbfb2fffcc6b1d19b26819f91e6511122215d5905eef0fc82c22af76405617aa7c3653041c933f8bcf97c7e5b7b647c9e5af08b1975b7809f85492243f7e990432303ceb04113e06c5024595fc9a2b19e535a714e4f564dcba13f58ba58605427552334bcd55d362f7d37e54cd0900cf905f09ef2b2040e7bb59f9b4b3fa3cb2d23190b4b6d640275b694c207293f4af11fc0bd044d09d3c13b2d22d68f7a4fefbe0925d48b956a4b516053d29f1cc43f2098ea9f98ab8608b6bc35e5fa96e665d4245c606eb69e81400caaa776d183f621d992d35c2d4c1b3fa13a83168df5b1f31f709bcf2361f1ffc246a888f239d7d3a58a1dac28af62eb0ac1e580758cedcf6227f8a1862058e5c1007751f69296bf05ac790c6976e4e655a53a038d2d41d1f50574f8cda2e393287342956d554e18727110b0b819d298d7ba8e7f8f087d2c487b02ea89e91636894fc03b284ec0d6bbef11afbc62ad87528d252d94ffa9b239965d579792cd510a274405a76dc59c3845639af82474f7b072e05861975955fad058ed44a2ef272984fb23aa8de3b2fd3a1a3902a3d69fd90e936c30bb360fa0bf7c82267642eb73842fc8131c6bff93c7909777dfc27bada12c6092714bb686de21b13a8838dc1086921de76fcc0fd498683a896a3f81d5fb837cb49e5782e62a9fd05065e35f87f3585a765d68311ed46e659b9738447dd4fa9e1aa2228142100d489c3bbf37a5dc181eb74a5eda7b5caba7c048328f2ddc23cec20a1c305859b6189f68d4a208037e692e4deddf9473eb33c332899ff9346fdc04bf8fae0a76451831d3d0c59bbfb4858ca3671a06af91d6a763593e9a7416c051fd3dd14f129eaf4447e9a95eb6788579fd8862c912db9c43020a8b8b09cdea3378eb2bfe0bbdae669f742795c4eb0d5fd68f5a5cad9dbd335c505e9b4f6ced1b223c28cccef7fe5006cadca69c3aa0cf173890667109d5248135dbc99031c0539db2a99162006e717ef38ee3db6494d583c750708b499ee834a66708d812c046c4176392d5ea2e495a4bd127cf3fdb9d61d320157f074e7d05c213a4497aca2e95a865ee03cd4305b1557b1f693fb20f1d9b3952abc8e7763f785341bd25b236c07eb06e6be89fd6dc7401e8d72e615a114d2006404bfd83012a079933e7e6e910584cf18e8a8fffa80090f8a3fcccabc083d35de933b076b74d7aa82fdf752c3d4b99e5c2215f3527fbc9ac6750bb0ff9fe3a51b03bd6deafe83ac8e602b2a9a32c94a7606c43c60dd9c0e87f2192caa30d81652fd4199b739d54b077d1fc36ee56691d943d6833ba6b46489fffb37d2159e02f7cfd1e3c65689a2c9311afcef2fbb855508423707b86ed96742a229ad77f6850f04f6f54442478290382ee8c96dc6ff482a207a77a95d2a27e65004b1fc4021a9d9ffaf6fded2271b7b20c5ffce2144f7edf40f45ac8fa128283d142c115d858dc746afc6e5f23bba11dc43d5caf5d10110b80eaaf2f32e935d0064178a27f2e69934e3e2d11dee869af823ec6a164a3dee3d9783956e16e094d0734a82e7b21e484222e5cb3012fe5ab182f27fbe6ecc3a6d8639f7c7979292c503823147d34122e84f92605ed133a8c72e9a21a4e80a563483f24c014c231695e912001fcc43f9cc9ae8f54aa012cbb993d39e409f5599823101bb89f3b5e218531069799295707e909066fea6450def5a3c05425264e123e43d0518fc55767583313f8f62eada68ac9f3a09eb6e59bbaa6b1fef1cce6d515883c7826d1bd5832171093cf47d08d2b11fb8b81bd75516cacb30f4b044311e14a4f502108b3de163234c890d3803bf0492569614e675a7db4fb4bb3ce4ff97b71030367469e2c02f40f134bb1b04c2eb65c4febd5c12d9807c28db0df0b3f4b20d9b63104448c5b2d598d91774ff92223b31aec088e1852fe72a6ad37ffa47160638db2df09c3963fcc4a9ba606f71b21d5abb891195dd5d71cadc2c59dad1bc0392d6be006918f9d29401236becdad3b9cfd2db0d9d1c1a9ae7398b79cf312c28861a2a17f6c779a4c882974d128acca7055fbdd97109f773a9e5913897f715de67a4137a710b3e964960da5bbf7343b0ecbc59c0dc65223f53493b688252e82cbdde3672a07f639c6dff9214a758f3b6636a0610517e15e2988f573efc866c97f62155ae1eea6bdc30f68966d32c1a2a81d355348f95707a27934f545880fca0e36b289e2c4ceac51bceea55acceca5c17e8f09e79fc2aafeefeba8627794b8eda18386d34b711ea8815594ca971b0ebd2cf54cfa9346daca62cf6f63e77ddaf88b226cd437d4ecd419c3ad51895794bd1950c66072ce7b295254cf4458a37e64221ee555f0a91a5081226d2cfa16b93b69faada9c6cd5114280f1b91f0c0de9c82ff9f1d5b944623023db2a474521a61cb571fce7cc53da24b6ce5e2cb555c1b097e67565737798f194068ffd6a1466ac7c851731c148fb291b1590758ca4c6f0bf77d034f38ebf76d95fc15cb0e399c072c45d1f8ab35b619ffeba90dc6ef8b1a8518054cd67a8fa9f426d32650b8ff9b40febfa877f2e7db10f28e95aa090b80a739e642c02bd918c216439bbdd3297c67a48d1b7faf89b32953f848e38628d67505e34cedd38461b932191544f3ce7deb2fa6103497f9b5d1ea3f592c84ddb4709b24dc66841b44308c23928af4d1bef834fbe5849509b1742196fad9acb5d123bca4ce4620f9d30a3f311651338abe4de495c3a4d2c1c62ed4fd2dc44c0ed3d98745f420f35aa8b8c6c8e7545d84e8951d6df8ce8dbf5a93c91d91f6dd3ec23a1f67090aecde90083302d1ba796834c0f43277452f2eb0d73df6d49d1912707bd0cbe260bddbbe237c18c4068a38a6841e9283d9a349153f2f1880cf58134b72856337f720ca9a1780743cf963982e32111e14c9c749cdce9159e1ea61ad6e1782ea5549571e4b7a8c2e54a259856cbd5040e6818c2de15e87c9adb0e331b25524a64c84403640cf32012bd579e894444c34a9a1cb94de81ddde6915f9e6a0f2bb278af2922f01217d62f5731b86d58f381fef851baf0362d34c11ea57386e1a1ec0a4710551f0398029096f2d0126c0b576203433bb1684402834b375c551478f2b7cba2e6a109b0dc00f41a8431573e2daa6a563882fe676ff4eac8b6c8f7cb4a2249036e74af0c2b221e8ebbcd8785f4732b5b42cc96c1fc83cfbbca3859c6bd0b085cd0486e705134ea11da18b555454449987ca80ec43a76780f81847b55462bc9afb08bcb321f686afc40421486bf39ec6bbcbba27b058f95322ae02e840dd4d86ed451ea8ae3ae7828623f2eb7ee0f5c38b63901303e3ef1f9c4688e040da4c51eac04d4ac2913fe595e1183af812dd3a9d915af015bc3e7a22736c98e610a43696a128bebcbc161440cdac727b85dc975a679eecb9f5acd9230067a046bade6211977547696dc220ae7041c23526451ea5923e1154c8c3d85936559c4115f3c76069290ee71861d7a2882a8c1c045b926552f0024ee7ed6584afd7a78f757cdd95bf708ad23825a985945a83ed62f054472e0c05301d493a20235b012b4ed60a9e2be7e7d0261e3102d5e615604187019edb3e6fe017047134202c7101a9845a02274c4300965d5bbc41e4282223f03489684cb4d008dae281d21cd6193b53cb73823897f5a799655330f8dea9c62d3e431b34fc3cd98517edc24cdd31d4f783c56f6f93f3616c99fc5146c62e833cc2b7766d09e6b6b867fbf3c0c6456a5fc0f558240eb16c6678cb38acc544c3c1dad34e92e0305fe9aa83a78d88563d416ea8bd08d8f24d14e0b8b9071dc8e9b5c3420e459d2f49e0365f515e3dad1b216cd5c38c30f2416e28f300c561b2781bd4253a1273009deccd843a3aa864b3a99847ff01ba0e9393a04a67bfea2a520ec04505a62b0c41e46b9c5c9aff222a5078f70b6882e85cd7e4424ff6cbe7c5c7ec57b0d9fbb458f7c1abee972a60cfc590adfed7d132caa98156eb98ebd82b89ecaf0f8ab1bf65b12d03fef6fbc5ececbf14826edcb609155ebfafb93f12a27f77b59d3bdbbf0cb085b130c265826d6a1d576259185dc3209c8d4768c129f7da7af3f9e7360d8d5d45ce93565c21847f23cc490925506b6ed085546667c97ab176ae1d0aef18bc74655bb47e7c03b57f77af9fc22252d06c697fc32d57a124c8881045c1d50fbe9da8f4acb06303e1c575798eb5d7898a42535bd0b2387fb585196a3287f8d9c995c37ab44481439edf76859df947aaffd4eb825dbbe0dd35ca42342836831443d5d10b0560f4ec41b46bbe1149cf96805460ea7b530e959d34241333785e264d04cb06b0f92dfc2f1f8fd76b9a4201d4e5fc8bb99ccb8cb5161d1a9d5dcd81c362e83aa89970bd279f4b89d58449d0c455cf57690b1e2eab1f2c6d3cd16a3d5c53287661c1c83262ecbb24be8eef1055a95b97c5ca891b2545c30aa57f0acccace07472b4bf5ce13cfccda5d89e7c2391b8aaf36357893d314ca80d2c3713f885dd6b0cbd566289ad38fd2e2e573297290d9b4eb17da8fb6d70cd1b36b626389fcfbe711eb12ea836d3064a6af343cc255c19152aa18f444e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha3400532d8c4e016c40edccf3e88688ea16d93fdf9f0d7cfa87345a5b3eac8f8b1dcd3fbe8da3ac0058fd85c8cde03c97697907258532600e31eaa4a855d41c43b1437856cffd08fe7466cdd163276a4dceb8d830616fdee9d83f34736fc771e49553a5ed0791fbb694b6384f9e89a1358a8c34045d90e1d523496ca749f53e6c8716c5c6dc8b18271fb8be53e8955ef860638f4ed4c4241af4aa2395659f0a5ebe0c082f74f61d8adc9599fd75a513db4d369b9a8ec7f5df7c7590b0e1b54c89948703a500889e162f67c5e25a9f6926c1fa74916232c5e1570eafd93095e8c9b9f31e0134475493be5621d23d1573120aaa008fcba5cbdad3765e976225301a10a5fdb6228a1f1325801ddb47eb928021e44d15b4d2c416d48b3b159483d7722f781b8ce46bf5519adcee1b8cea6094d5d32c7ad491594c923a83d789ca1ae5f9ab909d41d25301f544e96ca534b1db179b7007521499f148aa369846abcafd8bcb668ae59d40037ee18c5ff5eed4ab35fa8bd18ca1bda96282567e6fad05c0fb1102a48b7b20923ee0737d3e504eefcbd24d5fd8253699d7b6367618422b44ac3a59946a2a656363bf9192523b3beda0f6a38ec25077eba1de19bb6b2db5150e7004547d1e7ae37a2e41870c5adbdbe106a053bfb05dd0482031eb8294b2c6a59b1eb48f7bd43744f11f56a7b90c9d41388699fab477b9a117af823e5ed728007488dc2b086fc2dd37f71b21b120e1cec37bf627d9a31047aaf820ad8920dd9140b30e42c5ab08ce9fdff987926ab430858d59d228050323e06e5f3abb8f0f0360a94c17ba573e688a961cf7c819835ad03986999523c75d798bf882ea68c1bafbc07bda118a3f14188d01c1a335fea19d73a8d9fb9489ce0f444d3f5ab214cc63d0be8fc47ade1d291eaa3db003745dd03c523187d6d8e8b08a6c77ec2627fc3bb8d4b78f5e017d3de8440b2d16fcdbcf67082b3f8fdace40738d405a342630eb9ef6ade84ee2c895b84abb34bf0881e3504fde1beec160e8cf6d9b591fe07bb5eb86d41c02475398cd0cd8b8970800e5b4421d8e2e0d3ae26022c0878fde49739f7e9b7f5cc26ee4fb3711461e9bfdd7ec180c5e3f973cc219c0084d03735450dd2543433e622c8137555b8faa47b2eb3eb1c019ef72f7b9442a0aa27c1a7d3aa36bd3a55a10584eec0804258f5d8a5e6100a6f4afb8837d08a8cb703ecd65f895b8449819dbc27c7b249123a9ca19bff5e609dec06d5924660bb959ce7361927521b6ef51f47556905fca4b651b5de31fea3df4ea32a4b315b2e04b676d61b73873939da76e0003c38bb9450d66422f3cd403567b22b9527c6313c823d7f055c26a20ee410c224dc5bc8f2a33526b382494bbcac90f61e40abdfcb5bef05bd0f5dfc63bd177090623994d75202a437d94a246e2c78e84542bc223eb7931f32b4864556a736e3c7b6adcda373025b0a514f3258dad4f6070fe801d5393e645241388ab0ddb6f2fa469ac8dedf199e117e267a9e8bb1be31670fca58d67b54e27f3ef7a633b3903176a78700417343db670081f2703862bfd4127e56e5f07f0761bd492c3790d41d401ac41443aef6022c2b66982cf04e613c090d9ea7470666d9439b7bb3e8e5e1451220184af27ee3943bb5215986085c6f468c90411e96deea0b0c6fc8038219dd03f56dc96eb393a39281b3ac47f5af1157f6cf326c2ebd7d586759507f6262a3c1643e99e614945d57b3bad0b5e31c277994792fe2adb46cab43b9a84ec1ef3f67b619673321ee6ef47177ab34e804b24508486b076e513c8fab2f7b437c4ebd5568d5c99f9297c7329346faa59fb52cb86b38817b4422df12590beb6dae463a90a5c5c0b7ad0cef64e4c6fe0fafd7a77198f4d6224cb972f4abe522ba00c6efe73a4a5cbd8aa945784d88e374b2aeac285c64953faf90e8428033645ae3e68b5bca68c5c9389f168dddbc8cc6c1090188cb7c064da1553fcb0caa5125cf3f1c66f305f27cd40183073c2a4655cab85d8a11c4636fa95d6816dd4b9bab5a7ddd7da49eaad37937de39aa097f41adc37b7c9397ba65ccf74931db86aaebf21430ff081e9622eab9eb2693f6e1d8431a85fb3fb01628c099018e9286272ac7acef14fe876ae7f0068ab59a40d3a5a3be3806d04f79d9dadfaf377c2fc9aed4391be412291269c665649e10f2e582841ff069b3a291079ed4ff5dedb769d554d5031e522a31903f2b2ebe8c0b6baef1f9a1f2d5acb9f4fc21ce1988e50a9c54bfecd4c7f4804551e1890392a1b5051357d48ecae458be10f63cd75abeaf8cf96bd39c5225eb8e5fc9a4053f9e824bc1c699a63087cb804a50996384a716c3a9712f160188119dfead7c7d3834ae66393d698b25e14fcdbc21d320f25ceb912cfb22deec49ea1a51f05c51ddfa022419a54145d271f61ece29ed102f0bb40de66cba7283050a3b085766615a895bed350a5a1adb6fec78bb40824481bfdea50c647c867859ce049f7ea863b2e63bdaa381f20a4d3027660d8570d585291ccc7f6fe63ab8d26330a27a558b4f0186303004144019610beed61d8fbee8c05a740de02a6b9a31b0d1a069856d8d7e9aa2f6ffe9e9542e2a91de6d9e2fff5cb02e1ff579699d18371d0e3186546546ac12412f81d092d0f2b807a35f46ff2948f4dc5eff5e92a64a5992a543d81839247f22ac6215ee5988c35267f271e4dd30acf969ce8b48686c1be17dce623185d8823ffa534e112d8a7d6e1f86a9b0ea56e1de8a38c0a5c4a78e22b5d6a01db322bc2349b4b8b3c3d5a8246f8438014ee4a40fb7bfe04b9a92b847123039e726d3cba22d9fcf9270c81c432581157db781ee33ff9a9171c3a0f9ae733d720cb94509ec823c03adada1d62391ce1a9ade4c6e8e00bfee52ef4c7c2737283b2405176bfe2ef5f56f73e86861f0bfbeb5003f9c9c2a64f45dabdbb91bb4ad687313f99df352c1ea1f025196387a3cc6d20fbebcbe9198a11d5b5b349ee03e53b75c282bb18aa167f2081b59b0140d9e4b62ab7c78c0854d028cd273aee48f4f93f769489a0dd573154a594497b9443265c957b5ab236d2b16b9d350b0d87c5a2aec866bcd74715113255de1fd3e626cbdb730af052ceaa372093aa05087c162712cf31c525d57af505e131c9695c9e80c4727b1633598defcad4dc982c83a2ad78e05e742473a089b9f734b2984e8a377cf2f062be714e35f223dfd03fd83fe1714d31451e4a7706c09d504b06ba161d32d6d53f5768417f03be54cc55578e136c09bf73607be13eb4fc90f744589d9193427fdae9fd0723c4a6aaea1e5317438e7d9b0b5266e1ea54fd12b2212a82c7b99d76e091b1a2af6adee5125aa1605b8b13b4e81bcb5bc8a33ea95f39e7380806fbfa46c34fc9f34a6fc185fe3cc16310611baf4eafe5d0a73f3527c554e118b099b41a4d5e9372be9903ff4fd490a248494b2ac7057744921149868f1c8160bf389c735d7b883028c168bf1678d6d85730e50f6bb7007bc308f0276a819d9d466f234775b3d3dd29de01f8d00b5070c2d053872885dfc8c7b9868b2d748dffffeaaede257f33c7af131e967428e3f71104941ddfa6ff00df4e2c657a7347e16966b5ee2132c9db1a3e12ccf18cf745d902a14da43bec6ce578cc572477a6b08da7a6465d020f7b37eb90369cc1b169ba46ea69a48868a0acd1ef511e6ae96a4fe03b528430b6905cfb90171661f06a9694685e006de3b1b367866d71d9691ec713dd847ff612de04321f9a44606e9b52b980129b5e1a3971998613ba102d17dda2707525b8329db80eb98e0a9b76cfbef23339b1f514eecb3d87056e3edcfb82fd4476b19934c461538b2ac836c97a21ccfa2fa52c2774b37212dc03b2dfab97cdd51c21f1b6ec648ec6d357036299be21114f60538da8b275998f74082acf2d895fe7fc7d7faac59c6a503ba51bcc07b07b2aa31332111019843621dc01ab2915e9b66c594e19fe2eca8e8220c2c28899ff49aab2bfba999febe0d5e18545b4c734a7f020b5d757806872ea63f7ac82fb8de3ab480c0f29b2d5e8daa1c1374cb7f6203dccf558a096200594c4a65f7a497d79d3511dec6d595529ad0d9048419ee581dc75380645c605106905aea53cf3b6da6f4cac09817baa306425bbb0dca699bcba5a9c0e10c9f1ae22e90af4e40ff589e6f3baba54ff908291df5e72d9094d78310bec98b0a70110ab9a4baa6528d6c589a2a753d28332fb52975f739b32cda43e793bd9ca8612bc2e3d96f76007153aa4dc42e39d8737c88b665ac6f8d85f302dbd9c3baf25b893aece491b861dbf082501052cafccfcfc520d019a819e1cdc1a48693f22253d96ba31904bea52b3b8b50df1f968fa3c7c167c2b88baa118eed93fb2c76b4dc7c90573a796d1640e050b54e50725c7d3785f22059136b7c8cd9276d1f35fc83dbb5e186c0c1af423a23ef6af2e382ab105ca71ba24c7d2ca86d6b1bff0c9a61174a2e800a58e6376885a57f30763faca513596292b1209761f5889fe330be3e36730ad63a6c595a86568c20329134f4e1a19b396b015e711f3b1fe1517b8ab61366733b5fea553096c96b5e0c0f598194061521781e916374043b95c7ebc96cd50056a6ffe10c84907f6eed0bf5de5e7446757d2c05e2444752e4944e9052534a1e0190619cabb78363b071de06ce63d9ae2e7f89e48da5ca9e45f9c5a06654161580cdb9f159e4d596d17a2f1ef8bf24f179eb165d74c1d4b73ec081761f8ba680fb3f1978cdf206c8588dcd5b2ab045e099c4bf10c53664cf5d9084f616a7f658e80effafae65c73e1df77dfb2e774206ea7338a50163fbcafa8e63e565f2c4818ea54f821cbd31404128f763e4f6b2087290980a33188c4835032d115ceea54c80bba4696e16683962d6f21df646f762e32258ad0d0aa9714cde7b91a0cb6bafd66cfe3868e55e6e54bd3e9bff346d6a2d7300d052085d5f327678e9ea19138fe45d28f73e94b87bdedaaa14d089a933742fcd4d436597a46d438e5b78de1412c40cc8739dfc12354525be61f5d4ca818657336ec20afc3e8721717a7258779821fd35a13d7c2e126d6da48f14a71501961e19e3161f9483e9cbf2f56c22505df6d8245249af225e01563f675c49f49e1b4615a2ca24adc8e26b274074a146f8a0982d2c303404f5b1f6f691cd82b31a49a68721e6d8ead2049fafb73d4ebb60032cc22a07468c693b73fb0b4a87fbcf406a7e61e07c19c2f4f257c9d62d31aca16981a8b6be13a8f0c9324a4d11928fccb270a5d28c39ef65814a6efe4fa75732c0bddf1d72d23246504b4802a0f6993fb4ba05c4c44f7ca654742f81c692aecd043c66f911a98b572b53153325286333680edca1e2a02ea3df71d4b4ea4ba3f5b732c74a498a37c06df6c072974c73a3187186164633e9bab31d87718c120ae586297cdebae4f7253db0b3945ef26e958d1e08fe49e076653c1243b92c95a7251467e84abab67fe2ad74ef5f3e67b95fe127de631d75b75e0ebb78227499bc5c4c202c980603a74ee16dadf225ae8ac140718a29c3694495f87664c958049924d5a6134d86e781ff45a5b3643619030e573e7b4fbcf708ecf9cda7a7f3e8049895a4de5393af0c0bafa9fcc0d7314fa0cb3a27643eec67f915b2d1f63ba3414428369345d61974cf7f9e181db9af261e2d9d83270719c24f14a675442af83fccf8d0d698991f1898f734264a2d35c35606e5926036df29f09a212d5df1a97cc65e8026a1a5c58ec90b5affdbd4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc790f9cc2af29017039099d04653aac3afba86ac117c47cbf962ec828a82dc22d086ebdfc4e7fca79bbb901979c00c8892122041f9ede9dbccef907bce58de10cf046136fa33d1332800a15c1964e68e0e301658b03fd52c8cbcdf5ffb32099f22fc5aea5adbfb91e21e217f4744321e016f6c462f92dad061a55b95c7776436aa693846d23944d7c4cc0ede66f294a739ddb2e655dffe63fe7ba1603ef4186a232438e0e04adad35010920c83acb0fe96a1dca66747c0cd4a785a1f8e705fac626a07234b047be6d312ea8b5cedffcc038b404904ba8cebfc21451701f06b3f5a42b2d01856707559833f5b5ca9fdc6f2da28561703fe78de0badbf793b89a6e4d1437eb3ffe9347b3bcad3d72afc8fc1ead0287f169a2c73515f60cd9db3254fb152720e76c7e1aef30c2bc4b0e82609be9f461828fbc9488d1155388356bdf9127bc42b1fad6f4082a6c655e872a3d71eb0d8a41707bcda3bcc2a87c176d31f55af8d56b937bee6996252b41f61e22292d6cffbd59b1378621203e12c778856fbf03955ec3f84a5c113f05a2d8592864d8594c00ab2f9469ab42e2cce0b52616005e095ddcc330ad00a7e2edd5f6696ecbd31c54ab80494a5fe32cd61eea56482ff31ce60ba61c1ac7814871b36cc77b8fe99260f5c294a1a4ad3d400e2e0acb94576befb701afed2454bc69be3a85573729ec962b66e499337483b28b83f9875241f8bfb094b7884248bf4a4d09b277653dcdc591367508f78fd51885a71fb5fe3bcd46a1d21083cc1199d94b44b87a01412100080e657a8b504c80f766addc77169b1dbf4ac3f5e02c79644b0097a4ba3c1fa543a9d135be4cb203128a660769e733cf827ae6f47c4c1b673a15177f40270b444fb7d1187d3d3080d29041d0cd5671ad684fd3ce558f35e1ec3460b082ab0b9f1e3be690cc70af584a35a259a904e24e0a4325e45d9c6862ce2e42403ccd507cbf1d94156cc7331ab546fcb95d3d55b75b6085511943d24aabb7faadcbce6de7a40c67ce33ea09d029afc8985a57d8b17860658f6323a5a3309955dab3dfe870abc60cc7cf657c6306221f8411a889e44668b280fe0a80c80fbf71dc58ac2c9d52f95f4530e04d8c8eef9de033bee023cbbcc580e9df826111e7ad55b0f1198f1645424c9ce72b28ee8975d3020e90c4abb8cdb748cc840a0728288bf87b5cbc2d548bea008746301f2c3444ff3da3103b34c48c1c2c88dbf65e360d6e35f5508eb56ba2d475551eaa6d940c35933d31388770e0f6df5384f6a4b84ab975211194bf0cdb7337650449d9354be94a855f8dd205b9eabe5fd2d1650166faabf481bd3108c8464a8612988fdf5701b2c5ff7ff90958a8f1d0b29eebd3c584390e855e764b28ae430485277ae8a70575fe2e6498dea485e8ef09487e42aa3f3edf1910df798bf3a479048e3d07e2c79e60d6fd4fcd8c6b32aa62a42cd65541887391a5e7fc7e52220498e309e41e405c56a023ceb1a6f9ec5f840c81e6022f817ebbbf82c4815cbd51c46677b79be282fb0e490b4987dbf88f1dc4e60c2f5bc19b647045a72e4eeffec98bab861d1004509c4588c8ad3a8b226e2e0887d2d85a876446b8a4f903c326df8f8f7b9540f8e219b8dab35d24e49904db0b9c991de18622fd41d75f101ff2c04004a9f3f25974899d2af457e401ae535b17612720ff5f8df219e94337fd9d422ff6cf58cd06e5f2edf442cee8d91be170bf90e7a1ab16d29ae32066fccabbcf3bde51418574dcace0d629b34d042f85ceee7e324c2c3a77f8b0607d15be42d39789b784699fe791c77a79e0ae776918cc044c5aa1c74d8e636d0a23492a9428b57a89f087199702b363d15a2ac427e4f47a035b21503d9a4b717fa3d44d5d4bf2d8a7898e7ac0d4e3993330fede99ad767bf929faeb115eb3003068bb8ec77305a849b71d810a6e77c489077584a8f06767de764a98abaf71b2cf6637acc3f666ca87d3f293c92939913ee165aa1b9a53687a3bd12863ddeb9d0f208e3d7618d5c432a382f26ee0dd6a8bd4678637a76d89c56b8913e8fa4caa7b361199f5c1d56930906e309f795b4f4ed1336daa0e4ca49efd5a215ce21446e67dd6fb5a8574750aa3e08a3183deae1325891eac0479d97cb7c9b60e622844fffa3792f5f5b746d089d9188871729f5c740a2023a50faaee8a79641de57b91d36cfb8892741a6340ea95b26d607fb66c3c2a9a951b72097e83b8fa00040b81455753ebf1166c88aa350c189c209c9e68332c750b41d885d085ff4ae7f5550c98de59b8fd30a0e2c242adfb2085a391e0b9862d0f609d87edfbf3b1e3b730fbef7157e2dd45af7574dc677c36eb9d2bfc7d8216177c0d3a7f358120b8aca328179cd15b3a97cfc7672564a70608c2e9f341b3ec2cf28684cd237c9102d041cf850dad093609e91a74097118bfe0e53e55d28e8b44763cd774b3ed1bf086fa3a66b18bf76bf72bed23acac09f164686d4082b7ed0cab11749949168fd8e6c1fabb6e5a3351c477796873c1963b54809b9c1269964dfc5fef6f50d49be414e9205b2d36a81d5c62afb89c90b441c3abda143a67a86551f00b2d3f10c2440e936db46589e4e2b6758c687b70c95811d7afd9b43a607b512633e896d0145bf2fa35d3bbc8c7486e9d5185aa3117380ac3395a69ea6b9f4d2e9347efbfd35d3b5b7cb09a4d581bd532adb865d2f46fb0371737b0afa2fc1dbac405261a4fdf384943a0f03e03dae496d7d2a3987304dee89b25b3d805108a7eec73d13a709e542c447960ff74b9d9f4464034cea6ea507052420760597672adf6ebfe2ee85f1c5871f3b3e478c0442c5fac8accacbaa95cd58bfce0d0861609d1b3f25aa046cbdd9e713d0650b1a0a8fd08adc6be89d6aee0169c408fbbd46d3be62a715110e6286f37924d3bf07ba6186f1b4f2fa6c5bad68277e01875c92a563e87e599df18aba63783dd9434f9997d2a3e7f77926489414f83fec09f2c5645cbdc4cd3d6ad444b66bfeff84e74f7b1a4d4189cb6d1f4d1ef9a7896eec1caba7085d995a008df00c39f5febe8463daa2ed197ca46a295af3aa3b7a13e21d6050c5720ec45da7569191b00036a6dc0406fdd5d87b63ce569b6d230bccd0bb610804866a7ca1a017c4ad946a18a4813efd3faa6dde6bf893867bca6695b821926eed4755e7aae83fb1636be9b4f380105540384b660d18b27f551a3ab9159764c815b0ee6261080bc0746987026d0a15fffac1e5873b461f2e9f43cda0fabbec3449f31ee21dd5a7edf24e736e660a52aa75c01d0182462f0258ad83f71d14680003f6c656798495c88f6682d802e799f305b6a5bd87be7175b84f7adac25b882c968916c27b4c51287cb13f24c426b160ee87f9efd459754307c4b1fcf492927fb1e4326c2a12bfd17d8706a509f5bc0738de3fa267a06534b36732279c0633e636690454c611f259318412080f3221f2ca224c4ae465aa835c87ad559bba8e5049c16312c33d703ba81e8189fc9b174750141e227d5530d025b537f5b32fc6d942a0649dad249ec0649f7d344004ff594c6e6cee3d13e214160c5ee0742147ec46ec410868fc25e4bfdbba96fbc8a060676be6297f125a9e1f6c965115ba8f33378bf422f0a16621f32a51546ab1590579a654adc707e9042340549e8aa12e16ff62eb7988f8b21a6e734afd0e68ebac50d39fb0b12f40719a8eba345dff43a77db829acbdb42cd5c4084403594f391de1298464b55c6e4238e2dcb204cf537ab86ccbb0eb11da5d22fde0f1ee064a5c31e2a7ecb5cf42fa419214069d0077393393d78d2d5fcb807d507f4cd514df24eef682296cca85722639b9facced34682e6d5c5d2993a697aa17d2aea3ba76bcf53e5da0215151d0bdb146611961496ae37065ad1feadb93611539ca7799af2df2cd33183dc1261f01995c5945f076e6a6a1a1a6009bee55d8ea5a47cb816a8a587d681111fffad124b3357f299ce76a389f6651e62f42615ed7fc6c31c936b059d2df53d1c60c3851af2b13fb3ddfb3c66d9f9a8d4693a737dba019c1ae932b84bf2c7f21b2953fb579a537657156c7ec4132d1411e57ab3980f464ba33cd8994d60f706e1edbfca43a7f99e6def1faa39811dfb129b47d4f9d5a5a32a6ba0d3530619238f8f63285053d48401c80eb517843001059dccc880d46ec9ce9d3e1311e83ba28f79df278eb6e0f524b4d661f4ba2d923cf224414a9fb091f1bb90d8c90d89c648aebaabafa28f158d5e8e5650e43f1df622621ab1cb9041e0c5b572a0f78d581bb4f4c1043a1c221508a88d591372b603353e1c1ead01553c857b011e5df1e9adc21da230d15f69b2b9467a24727ca950a4fa472b5b58087b9fdac0260cad596dfd00a36ef93af63cfb10d7934d6cbf067019c0d7b23f4eb250fe6e371278f7a67ee1dfbbbe50b3862f027575c165806488ccecb9a5ea3aa8ac094e4a6a8e0e0bc0708294fd249423f631175745db1809828235a2c13aaf4fdbc79965ce14f361d70cc52ab41ffd0a035459e66e7cbbc328a2c7a2f2f9f3b682b1aac3349e9a219e05f622fb3fb145385be8f0ea2718c42e2230acebe46bb0ad34ff329c357364003329c3952209fdb69d132861bab4ca6b0f037fe3373f15e7b06cafb061155136f411dbe194b7fde586a75ce587e971a32990422bc1d387eb118f7314303dbcdcab05e3b83bab249b6a94e1732bcdf25677ace6a24ba91b582357962c960e4632809d8a5a6a8dc182a4ec83107fd7fe95783d871e813b21d2c8f4d33c9d013e7fcb97933d0856ae9bb5ed1c479f0f28c9a59af2985919b057c25f4963d3aa46d7d5c520d1a050d0c21261ec4d67e67f4909b6ec45bf02d5db2d1c04036e5f0f2186f28e55cf2e0a40bf31c547b527ef6e2773d0e1918545076002ee51746d536a22ab6985c75dadb05a3feae03aefaa6c29e9dcda93e0fa64f4cf38d52f538b095ac1ceacfdcd31560acb2d1943b11a0655bf781b6a72e52c8a2a87514d019556655320fe41cd6d0489f91008f3fcad1e8de9c141cc5e9ee58a04c38186ff39c0015a9f40c542d20d15507490884803830f9ca4d95d81f822c1750e7dad807253946e51c00ca718e0a8065b344768d0de759559b74e1b461a77064f9f8d4de808a9e6d8ef15a394306784e01f51017b92914df91c1d179e5e5c6af71e64bd50ab8585d967a0a5ce8b3935c5a5d572621542e6adf2b6077a79629e8c14f24985eddd7c91133cb02cf36ede7816635222dd7d8edd2aa497d87f1b74c0fc2baf666905869078a34ab29fa3859900480a72cf49804380f1f03af861a4473a6ffa057220d4c0209e969c5533c4026df559bdd866fa6bd6f21f41da16f47b39aaa1953a958191f1d49eed7f543e184d7e6bfb9eb2b386f6e0dc0cd307950a3add7e46b705847fe72a5e4c957f5cc527eb753e4f79669a6f8076daea73b7e45196f6b1a94ed9fdb18beedc7ecadc3fc2ca0069087f2818bb360abf18aafce7df84c246c51f165502472fcde1c34eface75495cf46ff201d53ff4e238cc0be319b9fbe0f8d3468e3b72b72e4fd8cdb8954cdcee1c29012db949ee44f1be432c989d1c3d9362f3f009023eacd63b23582ad2330eef315c06fc20ad428bf76630d863574cf877262a732acb68643aa361824316ef8f488a29c132d0a7f440f07b2f891dacb7e3e565b1230678a34dc3e32c68acdd7bda789d899563005dee485ce3ceb9ac4df79eeb016573c7c1c13f7ac993fb921a614b9be626b4c20de17;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6f907f7ef50904cd80d460a6f6981adc605768bee81ef628c2475d513a3a1601ccd5337d388f02d0903e5557c9c3d6e13129cd853f7cf0d0f1f8c7b9b7314d04875d9722f72944884b84c1b7349b752ac16b279623374d908028d21d22133b4405e84ab759ef4f71ae726d43190286532102999da0430d88308617e36677f24781e18c7d956f4dfdd9aa33ab756fc726e2cd5c09da594364d35ddfb061fe68e71635da7cae6ca30ba6c4c27781d88e24ac46a8d2a6aa6d5b92fa227c6700930e301bb15c8dca138daa3400f298f743c8640eae1dc23e83e05b579bb0fe4a0b64961f51759622068b3001f21604a62a860e4cd3b75384a679a6280fb87548a15a7157e5692e67dc3af2a1165b903b34b776a83f03cc1ed8bd836dcd20ab4abe01a134778dfe33e26a8a1213693d58387c7dad211eec7ec029e3bb3a15b83af051d294f9656a175433cc2875b9a3c17fdca0a8435e5781f40814303d5f1b0720412addbf04a0a85d205d58caaad31b8eed6aa00a65e3085aa8944f964f071d4006eb5788351e783ce89dedb4ac3a3fc30fe3b0cac39613fc4c6db81c19eaba3bdabfea70d92c2da011ffcd1ef7ba76e8adcda90e0fe478f7e7b9138e63cdf2dfdec53cb92c369a8a7d71c349d262766c9ceb61b2b4c7dd9f4416f1c32ee8c33e3fe800377a0a7564d23d03ad5219505236616c9946732b9eeb57574cb7caa89e9d75c15a802c1672afebfaa412fbe0467ee77fe3a65a982795b28da204c189bc87fae0388ec6ada45e8cd4f80abd672665506b109c749bcb3c0123be8c24fa3299e39858dae5eb6de8854093e8d358bd75204a7eb78ac4ad0b9d15d30fa33730e434503b64ddf87ae91166ca419ab036081c6f2d13814d1622a7f15786db120869a14e8b63a22f12befe0d31ba90e3d4de22c58197b0ae2fc305c485e4283b3141e77250016d1a6e29cdf37d34503d3dbf951da2499fe6cb4c57a048731f677146f468c4c1f26dde30b2ef737acb28c4f2f30fc71f3b725d7b192d8c396ed6919dc254e9659a00b828b1d36db90d1fd1090dbe79dc1ed890c2d54a0f2d543bb507979b850d5eb97540313ed45cb86dfae3fb51440612ed6ffacd899087dcfd7e290c692c0d33cad47412e5c2d313476e7c328867a94239655357f1f0467583170a424ede89e2ad7e40241f089a1456e8049c6e527ed956716da9ce49ef2d0638a783ca4c43107483eb27df1ebbce156155ac287f8df13744d64d943a668e1d21a5f471a03877918326254e411c2ccfd390743c06190cdf7a3251300efee6769fec4fac4ee85d86f58dfa038be3bef743a1d7c3a2e087e76d468a3dcc254d272c83c2edfab079a2a168b3d5c5c21c2e52db41305d42b75860cd8d7f9c90028ddc698a73297098f74bce6dab29ab27d69850bb7c4f38f0a237aeafda28099abe9a94d19e9c0210d5da290a8081d508dacba9d5c7cee62860dfc45cb00502ed93054627d9b8c412718916993d1b61047d24cccb390f0adf0912f28fed470c45989b5e4c760eb837a9edbd38281361b953e15035bc433efe541d4b6371cefa2847fa3f468ddeb2bc5d67682c20b72411dfd5a6c78689b6ef5d0f71010a88637686d80a93497521ec4c007a6576357313eb51409464d111f0e2bc5fbb12a3c3992a79b8585777bec7df7cbe157f9d1d5b7134bfbf1ea3d3938dc14995b44a20dc1a839bd253e367754586d28ff1c1eacfd861b0157379afd1c299bb89befabfd2edbf509ab820aa0d39a179a8336262656bb4343801cecec52f52e9e90fa708eb50a8d368cbfa2835af386aa91cf7ecb767bad5d8e25fe76da2b5f4a22830cc78c74e53c57750314dc33a6c887dd04b58fdcda1ae841f969c9d2d2f95892ab8c5ee67c570fcd3000d2063fa3345d23490b48afc88764161eb77b31fa648e363bd019219c03f4f3d23df2836ccbd3f56c13910766f59f88f1e12d1942f837ff7f36fcb3dbf2d0f9a387d3e6a7a8f846f0e7bf3f2a7deaee552d180a52126ba54f554925dc0a196fabb247f7ed0b3e2ef5dfe32094dfe613c41d6558fded3f25a491845b15d990cc73f4b48ddf38bcbcdbcd1c05ff71f3f4c9e0402c3ea57d97ef6de8fc79da29dab1f10970a549db813b5980cb998777fe7a0ab355e33975194091380599e735578171e389434365424a1799e57d648d2ff83c96f48a7ed9bf1936fef4d7188ff5691df566524dd1ab01345e7e65ca077dc62403404bd48ae7f948117fddf92583d84c44f7c568f8eef34aed9280709d3538cf200d4ceab0db744550515ab6a373648fa5e5c96c89dab04550dcab4620bcb929ee3b8687b3b274276ef6fb9ab51a05cb133684c11dd2c6974e4470b77cca01d423c08d7514406189f41a6668ed0c58032e46d874dac800fa2803393bfa5319921337ad791b608c5de57777dd63c35a95cc95c83f7e90629bd1cb0f581a528145ebe8b7875db5d765b2bf5682f91e4fdb817da69bd15abb751b2bff368ce6629ce8a2fcf8e11d445888290fcd7925992dcafa9d6f0fcabc608134bdbd16faeb9adc7c0ff793999dd9b21f3ee922ff12e9eef1cac8c55e75eece75239a8b9d38a214e49773a4777ba25380ef3224c7a299bae8b47940222a51d9cebeb771117d8cb2a09d8f62e586aec1e1f910d9667535bc0e991df5fa4d353b8d4383a7b8e8b369e4cd43b7183d16a750606796806a7ca755f8954434aefe8750a0715dd6dc446bd55d226945f3d7771840ecaa86d49afe3f35e35f5194fa474326e90562f00ba70a6d62603efd45d893daaecffde31fbe6f2aa03dd57d015fb5d0872e79084502817712e453ca5b09d438e7a8e0057a8851f673e096bae2f58a1587ed16426681f15d7caa1139e07f54809192ea23a4baad2c7ec489b1682a41957ef07bb0954dc3459c5ab7336f94c97a6a2660000ee678c88fcd01612d952efd5d5d33e56175fc26535ea546f39fd43c1af671e85d403c46868c80b8929d2cdd1e865f0ae253f0a78fc12e511f036fc4cd242880d67dd41875dfc6cca52514b8eb19d4c989dfcff5a5cf2ad1a93731b46a361c396f594b609200008d362a65184b304830724baef58f16eee65c6fd875bcb9098f39da2fc2d782c5e8a03b9cb8db33a9e793eca5aa6e8de1a93fb74aef03cec42a6db1e4f423b486649226b646b03e1a51e6c98322445cca3508f60c75b4dd53ab74830f6ccb9814119e0ea0f2514843c04da2892c533e03e1c6966ce3b0ee310d4f79c831573ea36d32cf1acb0f8b46c18198d431b43a4d8f3d3b129451c8d80df6a53ded7ef4e1cce898a37a74a6b9082e6d130adf0193b624bf845f04c0f6bcf86464e8a6496347a13d336b9d5bd732de3d6042557349a94abf0de8bd03082cca7081b45fdc76293045cdbf79ec63b3e5e39ba64236724d90d60772e9e97aae1f682f34243043258c3553ffd332cc09a1d1029f5cdaffdeaa2e47f4c31d2a7bfa95ad358e35ab13c6a09daf3505d7fa403bdc677902314dfb0950c0fc65fc3c424d0a41b68b54a56fe01997f691582b22c79c045ecc1b0603090256dfc2caab3a357b44ec5df558a4e3c0b40467a981395ad7800b00bc1f7175a0e7ded5cf0a1d6be7d54a8ba3e8428d615f0ebf34be8abe5e25507f5507631c1dd508a0c79d16877e8a51aa58d36a9d7f442d4115caa4a183df3e7a535500c45b65326e0b83b493769bbda0e4346475f331b054fc00cf0a7e6bdd00699bb049b1757384cf4198d690e1d1cd01e729517c1cfe8d1d34343ccfa0e726ec529aeb4d721865fbc040031c360ef2c9db9d690151d5c85abefa8c84ccb9bf9d3c667d8dfbbfe2bc57c1e59746ed0b53ae00e181dc7827fa4e542d8e6153f078224f8b1a0d6f85969c1b7f5c402aee2c40a494037cfa4d55960b0885b55ee1d59ec7ce3595e5846f3c7a95ae50a4a51dda294b6e7d7ae2d61bfa165189ac9f4b2cb68ecc522cfce2abf1ee2a5bde7c8816275c2a3f3fc78b58d4377988d42140d05170aece890f23e826265b6f2bb71fce008940436601a6ba949ffe8684948c6f0effcf0b54fc21298d3f430c4395803730391db5cb9c6668cfbf7fb5818b3d449004129da8ba1f8ea7b071497163f02b887c1846e4ada9fe9b7aa47a36bec476266e7fdda6fdc540f9ab8b4d0beda5d54c3adc81d15a5478f0c5f76c9fe5012f6142501655f017b5654ff910ee1d1c01eec91cc1cca50c1111126f8d6f423ca8f0dd4fbe91e1c24f79a511c94f4c818dfb22c0ea710041584f0ec8ebf26b985c85c349776c1605dac36341584980991e9666d3a758fbd94e92f825cc90c40c17015d1ab5387424163d3cd81d922aad823add041f064afebe9d910ec97add6d1101a0058d6c6f4eafe209243f92d9773c809f328305ff7af06422ec2907c6b1757b6869f53d7f645dcadd4bf82104ddd890417a0ee2122303a668384d907cc438a31ddd958ae269cb60a303ad1477c6b1c285c3e8ea54d71f1ea89d69c90cc1063f49bccf7e6678d0f35318c468720eb286a6eb1cdea64ec0ceb9f1aac3b9dfe5c2e7546018ce807802a9cbd37cc7b8f55a2bdf9007e0870cf9bd78376e060face0affe1886b68bdbfb0416959a415afbe8de5160025e747d8f51a26fdb576e76aef8ba271a6f65809329fef435d03550f81f164e0a1ef0152694bebe839ac2c6277e817b7cfb3343533f8cf97e6a45b522890864c35d9222af0b46d1f505d90b9be70497342bcc585771ffc3bc48cbe9995598fa817f26a7c6dc22150bc50d7d1fc41379089331278f7bdf5758e23b871c80474e5aeb3cb2f021d4009358227c55ce31114887e8815a077be26d9266ef4a84e96b222dd13846915067a39ac87fae18164f1f1df6940a291a22f74a1b714415fd6b4a60b445478327fec0decb052fe90749958e531e68806b07824ff4af97527b9ef6f86f48f91ac533176f587dafe8907c737e737f5fff10e5fa36f695a7b56839ae259bec4aa27559e4b2cfe6d63df8a92b4463df9ef64a53f917a9dd997df3816dc578f35508930616beb168bbc9d8757db2653e24f1bd1668aa5d61990eb8bea096402e134e6ebdedd7ca32eafc8dde7f444e6338419b4217eb23f5d6c58e6776d0c4c9b269f0b57c844f6b9a984fe98eadde9230c444e54d61f5698cfed71a35bfcc9bd2e29b928470aa7ea3aa76a833774c9f6a67b316997c2918be2ee4b9f1c7a6a646f1971288c4fba96901b4c2260769957ea8ac39c0002b96d27173d672071b4ca5d94959b24dae820c9fb97ba2127b4beb8dbd15f7ed5773d26f7b831230148d1802ce03f63ec56cfa0c5ce9fc1cfbff42f9a021cf061933281bff2aaf089504ce3c68235088107cfac07375b9e9dba0b95ec745ca7164696180e48846437013106df862f1b26f8aeecb78ed8c5521e73a9b5e087e777adea0deea0054d5d16ba32b33546d15ecb6e7ffc94cabfd15e3d661d62319cc7e0c64a5e9bdbca027466218bda3674b485da65cef5d11ea49b59475fd11ad7a16e88331f00e77f99e1a0011d32f75a9c1b6396e5ea2eeb3ec2a8d02ea0946fd96a803b952618526991df4b96d10930fd6a9664792ddba517fbf172bbfa6dba7d359a4410fd9f7b1a24792df6780559431e3b91d2d75089b394a8fce61e9f1788b167fecc63f1b7c71ea6699d64079c748abe29444ffef03983fa5781092c692207045dabf1d9c2d8c0fff8610a7083899f790646bad8754bfdcd8e9ff2532dec45a431bda5a49909793c0f2d917c1fd41c01268c36;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h35ccf13501f3b414603fa994c8eabd8bdae12ccbbdbba67f16af48ac5f5655203cd9b7df7bc81ef1be59ff546058aa9340042dc78075c76bee3e1d0b3aaeb9a754d49228717c21af0e5d75a9eb1afcc1756b4806bccc53438e082c3b52b3b09ae2d459e545b48dfa232bf57ed8495e1d3641135d701c88898d596056cae322a424b1e29b8688b8ae0d872978ee32d2bcb7bf0c6365192148fa83731881a420e3b3c04e08f5ae34f5305057383e707405a8252ac1d69c8a0a28e611188e353f6ace1e601ef8b71c07eb8f3d35ae757d72c78b168d90dc1d1cef0cccc40caddff7bf7f80ed045551c2ac8b84e8e79f0752bf35dbde1d4077a763033cfa0bbb73cdfa07791ea90f48c69f66c614e1687220a19705eb311d729540aba530b1c0185df13e0bc58bfc48b4b02929e452e5fae087dd122fe6301869edbb8ef8186238020c48f928227eed16ef0cba4f32ae8a23c64d734a0984cd08222a67b31afb4454460b9edb67c491ded636482f24dc25ca00bbcb4131a8778e5b03745636a7279e1b8b583022f1bad52c242f57254123c145dab36ec48b65f1bcf07b8e514f5018c860aab87931435b71af1f34291e3b521b86c3b80715222a46fae22e255a3fe785d1ef04507a60c44a02ced42023b60f9951e517fc05e20ff13ba796dfa9f20586eaa53466cf01324a11deb64fd18e7c7814e3dbd23bb52c15fb019eeb966850d62524727c404cfbb27b9c296b6104979eba9f456a187e74099cfe7a8d298d4792d7097dcca19d31a0eda47993ddada936695b2f270c705e0a925e3b662e4cb8b3248184a4e5704c3b90bb2a79efcaf728c183263149bef44ce4e62d68559ab6162865ab68b126efc139bedc4b307d1e09ff255b46e74f396befa47c5df8c60353ce10526607bc958590240be45a20b5e82fb0dc10b79171a28c6e3ff17d0f68948fd426a28bcaa88a17daecfc0c80717b8da8c3672ee19949c8b727205535e1fcb381437ccdccd44d2c310071a0cc3b7937592e42949e0d5f3eebf9619c960244cacd7aef483fd33bd62e485526936bf32798589140e3feaf7198e2b6e026bf75a41b5cdaa084a58fdc2368d71e9e022af36704647a19006c392b5775e3c64d1092824310d885b95c33c944288e2816d6939bbbd2ac839b6d4ee657572ce0099d64c919ceeb47a93609659ee53e4eb5f35a2288262e8a755f5df02c4c44b9aa860bb73f0d91d795ad83d1a45163d86ee5b2d142c342af662ba20fd86b8273b2db8bbcd7a287476431405c519ac3a940d69bdf57872590e027ef9a237ea1f1c4ed5ceb7ecd24b37cffa2ade73d568ffacfa8654ecc3b5d1143d34ceb64438d90ec741c5b7f7f32c608b3c99dec0f648400553609722a1fe3ebf23d9bb34e9714967ab2de52785e955efd6912413a6026b1c4d80138b2518a3f7cd269596d15e73f9da8c6d23b63f031d9a0bb8008626ce4113285de16423c8769dacb41a6f01897223ccbf5dce2a7b089ec67bac75f86fac2fe9253b3630a051cf149b59169b5c299dc5951ad9a01c8159c10a82d4239c1756e2d7d0c37185c76247ac8e5dffc8bdc142f82da218f3a934f5207313038cd0744931b9029df9fd53ef6c933438bcd443e03cd8386477e92ad60440a8dbb87bb492e5ada9ea0eca6b56277f7a124609d960c250e05b7ca74c38d40d1b0a3dad857e51a448a5146fcd125fe8e76eeefd22fac95084b18c6e11103e5dbe8ee1765de92931fa632e378f05d42fb6f5ee786911aa73ad20fbf1de046c25f34792369ba83075cc583ad6c5307f63a940e6bf486d0eb96a79ebef3e94bb94b0740077613f916002f4abc056a09701833a07e5bb0cdc93de84fb95ebc6daa42e0a41ae6848529b5e21e6ed8cdb1264c1c69aea131ad5df78813589bf85d999f93b5ad70e7f7efe4b47b0f4d6b5e8d217f9482c22f9ac31b496f82b1ce3424c5dc129893f26a9f5b9ac0b0e26bcec1f797042ba337252b44998a55279163fabe738e8d6926e807d6afd88f731e8363dc1acd3bc35d5df551713f4b4f1d0e099904e6bdf6e1786617546ac59dcf8c3fa60dd0e6ce5aef686153463dfd253812a6b20055eee5de4d591a519a8b7e65512541d2dc82cf5c9ae7531c10ac1485c449c41644b0f7575e01859031450da037890b6b9d5afd61139370d5ba78753ca50c42c300017ffa8d324e86d839428420eeea87593ba90578049e738aef4e275bf4373b7cdf365ce6608db3869db97085e297043de7e93a6155caffd76a5e3ae6700935f2fdfff3edf1999d048623d5c0c138d3694c7a6580dd2b0ba7040104c3a4bfe217cd21f9c1ecec633d6ae4c06d8b32ac6ba993ec932a9787a37561d9571a829827c04cb8df0bed43dca2f8f980a5136e00d521c770ca6c44d5be70a7030ba7761ed4eee160a2e620137206b3dea344a783b1c46437a09257cae75ce326e9e82cf242613cf15a1219e451574e4ae4b37c625d330d1e0befeb7569f9af76635c6ec5d1df1b956cc4c7c765c0b8dc60292334f962983c5d1797c2f3b9256407ba3135c6da029baeb001d90558acca2459c8419ea174c124cdf857a9fd605d8f57a5b9e19577b4d771e1f00e006f9a00b7668613cfb3379ca802008e4bf3c5c574d2e4bed2e597fdafd39a0e64d86d451c0bdb591b53287db0171a8b26dab400a6b0ab0bfda2cb630b004bd42c6e3eee28b691a57aa6f73759945729d25bd30c2cddede4539df3a96e4baa331693b1bbf910cceab50d7c529c1d1c66d212773e1dd83590e4d201c47c3ed82da284d44bb907862dba82ad6ba46b755130535d6b6911a19f37bfe2a8ab3c28d012e12bd72926e619107315c6c19eb077feea8e721ccd35ce5cfc6c524335dda6c6a5c3020f7a7bdc16d203330f9d20ba22af39f4df2c55c35dfa41c8d82dd93729b227991c02be387e092fd4587e67c3e16026c23d69bf1999fb49bd80a4bb93ac1ea71920ec0b1cd2d537c8a005e39a96e1b90ce9b63149b17cffde2f450b48cf2fc1f34f067d0425837a1c607ec19081349e665dd80a7963d22643432f5818e6448efa1fa5f21b62fe4aa96a9f8fe94d95067626cff444a09545b9108e97757903a6e7a8eba8baaad109ec9c41a918dfda3f0422f586da5e6a1c52cf4164017c4e6a84ce0acc82abca19b0618f4178dc405f81507e586d5fc100c1b60151b1437a0219a1e30ee2c9433c804e65a879bcdc44a93bbddfea5f5239699fc74112391700dbbd62a4d9897253e55b10c7709ef652b4d5317c83858781549c5f187e3529a367fef3eebcf6e1fefc2469dfc7012738050d40efdbb55d9e5bf0bb694f50bfb08a3778898311a991b7c92ac1d2b08c63c901b62db95301f58461ab60a4271a01c2697e96a807b97be88313db9eef12bcc57b98c226b0cae1f4ec154181791111181bbbb623d762a5e432df8f94ae5fe566547013e1a461534b5f7cc5937f35edad4b032b0323a545f25466641ecbed31cddb0ceae685ceec00b0cc6e95b5e3a23c7de3b0afeb0a2f91db120575b31d333b7ff0bac2a4411151ac309e001f671b7c3453f1f1d1a052ca539a212d4f7f425a6309f3b4ef1f27f964567f92df1fad4e63f5050efe1a8eaf791621c1eab0a6068ca4f70ddba3db416ca72343a6e67b7767be6742ab1e15a6305e512425a9243ba17eadec67a42d793a30ca267938ec8f319154485a9a7a76015ca136ad8e650880ab8dcae8e929b3463dce229a84a43726017cd5344d8b5bd25157ac7257d50747e1b458d933aafaa8ba5fd4e302586f295e44eeb30e8219158f05892161f774619a138668864687c75cdd9044a2218bf7eed8f79a2445e7619bb355b2aaa819f1aebafcf4f527ddb2cdc0d1d4fa4609854f37f8d8740a868a96d5490cb1df43c67e911adfa71392feaa99b11597b6179abf0a440ca17c724453a4843726edb1bcd4098b338aa43b5696a2d234771fa3913e94109a80311d90a660260f1ffb94fd9735c533c75269c5eba2e0ba7d098c451eb9cf4b0df7e7bc1583e4a83ac7ac9f3512f6e1bddad3a0efda3a4c9c9da4086826b38036b65ca03e3097a9850438c3e001dd7fe6016acc2d231036b4beb379161d35121bbefeb2f40a5cbda0400792c68a16bbd0f6d77d5a0f9d78f2cbbe67ab0e42e1e09c6931242b204e4e973b0171c09fb4ee0e5655e5df75f1a159c29cabff73edc3b2a4ee604a39dcf3e704af8f8e6cd3d7411267a0e7b98fd02f7c686b33da79c53b10a9f060a32d1b486d3638d9ebe056655e68a842ed831bb4b0333d67d2c1cc8fceea3bbe74f1f74e9632bdbd445bd3d6325f0e0035edf615e3b1220d77807cf2dc6f36a743fa466111a85e373f21e9a5307a3d226fa100fdf0d7a48d5f2ea6e37683583c4c70557040764a19ed3c159bab0107608f561c89d73ea5bfa413a7b5b4dd27bf3e5c1cdd2c0c1cd20d903f54ec11f4c209c7462475eb9b5c7960dc72b8c6ab5c611ac0f19264dc4846bf336d77ec317b7aa277f181e3ec2f4962972df5a02957bfd3a111e81b7aba3c0aa08f1aa4c14d45fe11d94e5354bdf4e46bc2768b45b0b04f5c56d3d40a9a3d704dba74ddfa651f7d523014a64180250f8319f1a840b95cf6fe4d66d5268e85ebebdbdf7ebaf3637822a7c0395635b687db72f57f2e50216daf0465abb8f5c141921a62f86fce7cffbc3fbba15177ec7585e6870595d339c49de0975c92af7078866b4df4e4d840e08c314b6945cd59bf79682517aa5f0ddd7e03417d7bdc17c725fe4dd76150aafd2e3f1fbf5ff8b1fdc178f09bf9e9c602d9fe3f8cefaddf72100a6e374913a1883759395c11d1e4788cbcc68a948f0719c68a17ee80b44d054332b105d9d08fda83d0d290fe3715d3631a409caabb4acdeb495232d89fce922b7d42ed1c4be27d143817a477046dd0cdcd1f2f3fbe0ac1e5c43e0de61da2ecba0439195158b654640f99c6192584ecd4187ef1d4a12546b816dfc349fad753a9c94adae3285d79f05a2834a21d096a1cd81627028d0a33a093c40f1e0ac7b0ee02b3264046f210106d12ed3fb337bda9cf7b28cb1defe6a66af2c27b5864bf45c319575746525d71a1c03262bb9d5e981b40667e18d4dd5697a1be2be7a26dd4a43d34b8c7e7a6e71e505f812e39d95563ed95debede08a9f6c7846bd71597e7da062e1264e0582b7c6afb6caf8317f3a72cb57d949febee363e24fc5d011f7688c0116b9f43a3c59bd6cbbc5bd3c09d07658b5980b2f9e6ebc9c3908095e3ca0d447637e37476ae82df3fc3c74b0d49bfa71f9541a75131779620f373d3002d08b188edf1dabb3aa6aba4541c8d1e4fb5e453c5a84409087bc6290e9185c10b779199808de8ce1d4c969fe8d2e7a7013996513a12fd204bfbf5e341f5d2c5c7b4e1aef01c695453f78a9dd4d37129352d1d92c07c6d1a12b8f83f232e731b7d8ea6b8396758f4f9052e73b06a95dab401447fdafa3cd57c3749a6f548127a21ac67c3344fdcd0d0232c42fb6e82f05835313e9eb0c1208c82411f213166291e44b6553f814ea10a793734075f4552515a79577ec9e4c220c56340674c4ecd5ff2efd0717079581d9bc5a9d2f197cc95a30accd809ece85c19d71e23ba250b33403ad341197d7402cb8c59dbe3a531a40b002aded7b29f1574336c81372a263e5fc0f05e9a0ee077e7134d79700a7ec069cd5178ce9a298518e9e88c4c1fd24a60a6eb8830755d23799cfe0fd960c9d3480cef31ad60d7ca69706152315783529a9817e48c36137541d6a01d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h79fe3ec1920874e78dbdf0370ce7150b2d64b47419ad789a1d34db350175a7d15afd580312680df98aaeba1883c031cef3f6fe2a7d7a2f48fcf4302266246572987d9f7b62a77b868a7b856c29b39cc963417c9fefa18216eeeeafeb9b5d4f95e1a984e91bab1573f0b9e18f064e73774f90900f4151de14651cd7bc5289ec3e9931c60725a6bcb30f17fabd08a3abf2e680ba0b9248353264fd93f5cf00aa083f1c42dd343f9a687d1903826941cb2a019e64a33c783f56f46eaeee17fa41831143495bda9b5c86f2751f56b3182d3b58c891071ab4c6226cc31b6c73e9154b30b74099cbd27a4913cdc07cd38466a98900e21d4259eef734418a7ff3750ef1ba9332f19736616d30192a5d9a46c49e5f5e03ee2cd144760aea1ecacaa1693b925703203102d7e74441b7892a9f494f52d1bbc2013c8b7d000f0899c150c06d92ae1ccbd075c6fa8c14a92469cac7fa4349dea476498b9e01d57a997b7c9767146675aec613cd7a30d0c0183ed8419c3780657ecd9a6d98a246a8113ce1f7ef9c8ded6a2b71c4b9d9f9cea7b42d6bec2d5a79579663fdb005723c72f7760e85b14bf3d0106e6fad726848505670bacebb37619cbb1e6b58ebdb32b502984beb62946de0dcfb9830642eedcc54ff3ae1ce6aee0b210e514bfd559d455a904fa71be4302b592fe93addab193a52ff35782e8a2f53fb246b5ae05070e3530755ca80def837de389e33cbc4c47ce86026326d3a479cfffb3d65bb3ef7457317734b5d3c8721ff15a617bea0364b9e0c66d43f05535cc793cfc81195eb391f7f64241061d6178a9771e038f89f64fb10fb80b4916846d638aec16a2b3a656e2a069ad3ecefc6def88a52db4e65061f2ad10cb9cc8e764ee6f791daeb5a215b809c0f1fc141e0bf82efeb2192d402280edc85ad00690a7f0db89914a3710779cd6e3023859a36452bd9a2ccac063e3a64b7c97675969f17f10c9f7973fd4fcd480d813b4db09430994a599d2cb9faf2704eac10ff910141f213abb79efe68a582387237fa1390a2e208321afbba09509c8f359249ac0b22fd986950ab790d753ce4e0bbd3bd883a9cf00bed6163f0315e017bc16b8b2fda97e8abe157a5f16aa8ff60185b6d4d57e2c4e5747dd41dc4085f11b884cf240c677d9bb061e6412e730d133fd335d05bdbc465046705f633821fc48bc8aa2ddd2c26f5654a1a92af1addcb16733481dc7ce2265855e22c25158f9e35d00316d5fb7d373c819e4b4242076af119802519a8561ced2308601bfbe77ae2774325a0cfd797aa342db0bd713da1b7ea519710f1044649168a123e445cea2e0227060f8fcbd9f7b7437de628c5d5ddb852a57c00cbe0c31bd11909dfb817fbfa64eb7b6fc7b998545b7fa5079f3b2001a8f1b5441348d82b5075cd72b26c0066a100271e8ee2e6089a7aaa2a712b93c58465f36102796453fa9e5f4a192ba8c0af4561419f96ce473a18fe68cc96a6123e212ee54a9e7dc1f6b411ea68f49705b1b6ffd6f6090ed3e1fd7a0df6d3acc5940f93e9df876e2c8a9a0a8f2f12bccde8f8aec94c31af0e4b3fcb7fed32e8af3102af61d9166556bdcb20be9cb11701634cb298a2c925f95588a5a25ec4096576806728c3c88e57268404df49693f426c4e934f2218fd77840c6781451c531e0a03010cc332c80ad7b11dc04aa77b8f40811ff84488dfe266529e3769b01c71a96083a0f452298c87674d99e063f72dcee71211ad39191f57ef50b685cf37603f5ef8df400aa26cd48db7c6d7719e0c83c01fb91e4cb97384c8ce54ce272761ab3e846c639e26e2d614fe7b1357fcda40ba7bb23380a98189e9555b73b55832a6295ef0da8530394fab7e05e775d1cee4494d79767dff5de4c02b81b09f14a095cf7816c5ef71274b3d38fc74d7fb38375e82fd244f15075066a8841672b7631247dc9f265ffe116529dfde0fe631c64a3fa17d452b850e73d5038d53cc61fa2d92d680a1aed694e448a9eb36bb4f90016316f595d647265becb66794f40132ee9fd4f523a1876abd8e278c4234fef5f1f3f62526aa8047503e9144e98b513f73500a3a6f0f2ec59a9f11fd09c11ba01a64859ae624bd97b8d0d2e2d80cd68c3cc53169a7bec9a8ae8eabe1cbcf0bba023564bdcd872641296bebb795f8d3ce6a6aceb544a81e71e1262b73cf5d060d3942b5667eeec41bc5930d41332e51ad9543169c76bef84431647647b793c17f1488d2661be5a3d87ccbf57fcb02471fdf366f7d49887d58caf10b055298517ff0dc13c325a299d089441be7d3ec86bf706edb6a4e8120e66361da706f06c6cf8cc802d9a61b8e8a4273f8f1d951ce24c1e8fb8ffee92f49d31ce43329c79aa40d983dff1e6735a11206e006c3127d21189b481fa3a6586c1dcfbe0bf67ffad3c20a579a1f363622b7c1900c6a3892aeb13fccac857517359645a1b97baafcd15d505c0cec7367c1cc9d5a61e8a24f9c501309009b202e113c7aee62fb9da862566866ee33f263ddbd4ab2f1cf72e64ce0bacf7c277a5d840d48bdb124b42c4fd176438e9a7f57695f24e31b3ea613d9d51e5f2c615496a48ef82764b6414f3af4ae80da708b3e52b6a650d96fea4e943e20e61e1d93b410971a47fa9eafba4e0f2acc7d40a9964e1119a810c7e8798289fb37b65d34a6b31f619333b71a68154370f142017112b43679ab7138bce2c21e89b2cef42a906d6eb6de8df221779b4e07321d51e327b32b07f67a32840c9539b2f0a526ffe189ed16065d6f6dc0302b5d8df222904df51560c39cd4c93740e485a675abce8a33a95831dd16eacd426b8164e377a9ea58b0800d1f9464debc9239c9a5116f8de21c33bbde07ddfc9d28dac8972e08f4e5adf2e2ef7cfff5a142b6e6e22546d8c8a0489c9584944f34803bfc87081dffdb6b4d25b4440042d0fff7f438de557dd5bcc1661f35d9fd4ec8804bad46010fe64449eaeb03af3e4c451cee8d8fa8e818010467fde324483dff3de25b07923b5a5a2be25df956d71fec95f28328936662159c13a3430ef1e964b9b7c0095e5502d223d6472e26bd433329ef064611ab45f33289afd5b19062a4a3130506e9796868ab337dcae4309d8bd725f33354fec63c877b0c2f92b26fd9f1e3df408b66cc58ca5179fae3aa8620cbfd58775fbeb0cc998f6d1b2ee2d5d532b2d40bdab14ff463f398f3007c0aedbb0f30eab3bd0441424a53266b3b120c0da75642dcd1cffba51e0c63f1c9805d4e7ea5fca4a17b4901aaa992d62ff6e32b89138215f69e1dab7330a68cbee3a6822ffd836210d9ea5b9a51c405b965b1f27bc2e75b0933f724e6a236e9383dce866b1541f4978364eafe4d54212c287f12bfe8e544969d7f17ce3811fc3dac1232d070a5223343d8e51856184698c83f1e7aaae557e1832e91018a317bec0debd9a8671b24601deae6e96454f75cc389472cca6187a3fe9d229db7ea972e5e023a91b45ca25b691158dcd6892a5f46ec57c45b5dab3a310629e2e2e3dfc1023efa147bc7f53d78a640411f9be73365f2f223cdb2f7a4cb6e16dfa44f6750303ec69169efdaa0845dfcfb23a84ad3eba5d23880a14c71cc652801a365f200632bfe98fb288c632184d7581d036dca79e812731ee2c7c62496f3ef407337e00cbe915e1e220e7e76c6b6f69ca4a16dab75503085b61472015bbfc2c15fd40f624986a7210da742cce0060885a37c82c7cea812adfa717c499419318cdf4bec342dac3830ffee1e31b1789273adb4a33d4423a6d51337e542981a50510cf2c5e062bd9560e5c8dc2b171bfc3256bcaa927cfb5c3760a84f2281859eeadefd7652f0f6abea5f3a2eb0acd063a1060a5675b86c73fd2cb702acd7d12ba54aec552502a7823b923c729b9788f2d98fae239c29ebefee67ea18c43962bffbfaa8b29f66ac3f7ecc1276f87bbb7633141a36476e1e1c4b9fd3ab1069bef7ef4ab065893266f366e3e1ea486140d45d792ce239fb9ada370dbdcbbd10a08893854a0345ebb8263e4b014d9a0388e706588ae038bb2d2e326d14dc5be17203c94df29cbb2dfc7543873a3c63afc42ab3a27b71f926f64c100339b195d78c991d79397d6de0c2ef8e31b025ae20e116a0a6e7ebc28b1312578ac7b601cfe1120832590d1ab7e8bd157c2b970ca9b0a8584800027cde30531e7985a34c858f8d151ed0276dc024df1bf21cd65202b784d3779b72b544c17979de2d51d2b42a77afd5e8b4c8025552a3587709b146613801feff58fb862f7966f1669e32792b635af536f32f6861dc5af2172faa119b8cf6a121fe2cddfe302433a0fbc58a5b3bfd809d83419551609cac171069b36a0262e227d742db1053eceafe8f45d0b8c0644e8cff73f6b29e6fd061a1881e8a81454d62ac060cf1d345fafe66a1731143a5064aa121135d212d46e91e3fb33bd3b2e0057e814257a868167697c38a8f35d34ecd63137bba6308c5105366449153fe3541cedb2e92307d2e9744e6d4436fbbdd5387a19c91a729350cc1f2e9eedd597f92b22ff9351bd9815e9101f946b1a7301353383d3f0f5a2de20568d44e3314232d5300e22f3e069fc8fbedfe2a96b4725152b9a694eb2c19ab9d4b2244ee7fba40ffa1d5d316d3bfad66b3df1195348193dc732c4981dd7552575fe763f63b59f233b1c8410b6c79540decc96652f427fcdfe72517843dc53141f836ff3211e3dc1c2ee91eae95be6400d5f052e14fc2638026d888c0949f578ee20774c93b4197fad81fe409e1c3e4140a4d250a0c3567291d8d61ac8c8b581e0b2bf770575c37ecf34cb7930265848e709bd72dcdfd183daddbde728767f4ca912fb76d5b8c70829dd058d4020089e6131715d15c18f1da75052f6aa6b4e9fb79c98b9fda5296ac42cfe2dac53dc420ab3ac5952183151b7dc395649cf51a415af40cab24d628a7721076737c0b1de375715799e6fe558780bbe15740e19e7f7336eb5a0c8acf29aac2db8eadbd871c4d507198200f37cff8f593c5fcaabdb03b89bafa3964ae37d065277672c729ac0c6c8a9bc74e36547bfac7644c0581e7fe36231b1f2c85059c77df85af3f8ce3195b8ac4a7953ce8e8204fe5861814e132e1e62db0867dbf83fd822d6a834a1150766a194ea390b8cf2ec8bf5ce28d4e3b28d6160a2b64c0536b85aa77f39a8676f49f30db901123f2c3b858b3ad1f47798503cd3e0ea1c10339a1c7ccb823ba031c6c40de9a794cf18b3f22380f9d0c48d77092bb4b6737a28736fab2ae1bb41897d9f2b2b66c5f56a029d1f25e1f5e996cf2e5a3b6804e7e43a89108a9582b9693476333e92607e4dc961adb3dbe33cde3900d1a20ba75c4b3db26351b4ef08ea689c8ca2348a97bea6a9d3009fe066f7b00937f39c2aef15fbc10e25b969c9bbc209d1e0670c6c9d7fad5484e6452bcea8dba17d0e882470582874701e03b40faf17cd70a67d29a22c467aeda222422c6957ff86307d5a46bdd65f96148717b6b2c79e395588a7360bec2626b6107e552f15454640902ece398905c7af5d1dff9e5308056a4b4b38cc37afaae40c595779a7ed67539c16f2d8e796d31f5c68bf802f22c0c50584f5fb3db0a11639d9a837adc4ab06f81446c747d0419d6dc052491e570a636823f8d9e04bc561def04755ec55290d012811d5763e99a654b10592c8cb6f04327cfa9172b0afacfac81f08b6e38296a29c9c7d4abe20bdefe68a8626e40d67f94cc4c9f35a5616b17a800363cf823cc69fa9bf21f01f8ed629865a16c944006;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd73a85fade02c3c6a2f586b13f605243378249a09f4f403a244f7fe8cd0370eea4493383bf985194a581fa9b07e589dea0afa843e0e2e6459e52cbe1b63fb5e0fc3e805bd1bca9881bfb8a48131fcdc02df41d96e60ad14df6e0883861210b8cd37fc9f53b24cbe9489876c46d54f52ba32a71425ce9656a9118bb0097c2a0c5a407f5f63dd9b35173b57434fd49517de2fa2ede76eaaaf365567821929383160eb44ac76a433ac6c38ca60fa1a2519263880483439d24baf37da42a1b6669273dcb85c3693afdec2306e18852a409296a5add2b72bf6bb1e1a31717d0300f9d31d2442bb55eb880513f391c9984158117f2cfc705a6e1d1683f0c2dd64dfdbe0010c4299af89b59a38066b99dcb12d96bf1384d5f9f780c1b4d609e0a6d62b5283d08883fc0288c7ea39a8c139495a97fc0bfa63399ed8c920fdb6ed19f381cf3f4cad1d06e19ae4346b1978ee379a856ed3e8eb442795306ffb976f9dc9775a5554b66b3ec2a85a9de22d5466dc16edf69e6711401cd774023c8d9bc8a078649947a8289c3b69f1ae68d356faebdf70343e6a574d82d927361f8f77387598be805a855f1d43ad3504ad7c3bb5522b490e958b6bd7a1002b2d85b7b99a23e8d7a69fc8719b1263ee3ebe01f7c5f7859ed4fc25df51923461e507803c064740c45497d0c8f6f6f078169ab86217b3f2dcc804f6beaff5357181456f125276faa79aca7523e4bd45ed522b1f2904f7f054173952decdf2cd5cff75c8035521ee2b384113240866fe8dce83a5389b0e658bf698e28829a7a99d07f5e005f456677781b346bc557abe87cc4015393c15a8608981c85050dd98f3901bd8b51d13abdd9d27d748f128b5b613eba0e28f83ecafc44187fb036b00645d417d03298c4521b5b1b6cc0b71f1cce8530615ba0017d5108d0a9bd29af0459be208970972305ccdf73ed50b5c02e70f82a0c0c76dddcda7972cf50a1e1a3eb427c15b6687a82d5aa59f2eca961406208d1be5f5200bf6058aa2707b11e9fe8ee9879a6b66f74c7c8d1d37f469dadc67efad0df6312816d29fcb590d0e8f270414d4b5ef314039691070475d4bd3f1feb77d084c00c73d8183d2e2350a4e3116af0d50e090014a44a08fb47f9f0de22a4e3665cd2ee45ea25c790317a18bafa4f63ecaaea7df53714a931d2428e252fbeb3e4e52ad7020b3b3ce68e2c01ad262795c3d341c02aa37b91e5dea616ca4b7123a4faeed4f51d038558230c204465e386db489367e7949d3907c7a4cf2cac614763487ce7cd32afbbecbd23da0417320d6e219b85485243235c1ef9300ac16e4210ce1ccb5bb6ec6b6d50c608144b469a7e7a10ce261e021d00f290676db97d40f3837dcf9905bfeab230e30ef29eda8761e0f12ee8d2440f19e114c4d8c4f66f986331df831417ec0f887ce39c4a377c28426fc838da07d3cd32a77beb9005ec441348ce1a69541e7403876845b62a3410f6ba4e4e155eb77eff4d31e388b58dbf22fd1521f69b4ba3ff87d8b1ef8f75773d1e911197b307995e7d3a607c8b9668c108dcb6fd82b38c18ae5d85b106b7b9bd15e768600aa947d3edb84427fe1bdb4db0694c957b76c2878be37741c967301466229c47042da13b9d8fbdc2891ec989b78c09c09d727ae9e9bdc65d9aaf1393559661803132814b0939da177db2fcb45835ffa07c81ac9d8a8ef49c5401e4928f54cd1770d5221c55f9d38159348a3f8c463e0e95e62ae90a878301faf5a26edec13f389f18b9a56c73bb0948998acb0d819389e09fb5db2fd2b070595de9357ce7ad613f543f6802dd5764348053ea43cb77a48b9f621c86d7fd750f2f0444aa31cb2012bbaa7d997bf5e67920240470bc2ebd40fc80801c803dfeb8dbafc937690fa85d5e2f64f39943a2b1bdde91884f573306cfecb29a33e2b106f719db604ddb2896279db266f35614b8044a1ec4f13e46ea2cf1d1a88583d1a229a6c1fdbff13620d910556adca95814db72b0c0c64f693b90b03e384556c3e65505fc5dbc6ccbd914a7a40268748c6ad29f228bee17c9345650f0e6c434014e135803af8768e09ff32367e0ae8ed91b481885f9f0d78d5ed668e6ee9ac97c0379ed112afc902c5a2eb54d434e8fc487438df460288dd2008a13c827e21243c2c76725edf106656cfa41db59aae56d6b7c034c3ed2d92ca3275b80d76154664ea9646fcfc4a9fc6b5aafea988611a5ed36be83d54a9b26a9aaf658d77f56e451503485fca7525fbb92228155b94e9d98435881d06da12b3014ef2932cb774e3c460c7112b479c24d83ad1a2d151055d3d2c8b0422c81d7471bed8e49f90f10ebe4414fcaacfdbdfca1b1e5fd997d5f1425df1b8de6c7be82228cfc1f8287449418f4950d3e6034ffea8cc1af4ce141c34a57411738b0eaa11a022a65852c370cb899aec7047e352703c59c4300987c1986ea5efd3b92d65d0723b9d0d8d9b1085a97b48f6ae08c53188df6f187ba24b31a7e7e795ebec2bab39ac9ac89349d0cec938fd97200ab0715850050d1a1467ab772c7cb6af478380705daf955f24488e2bf1b613176c30d75f69e1342cdf887e2e0e875ac23973e70985360c669e57f1c12573371e2ccafbe6e2dc8effb44f84bb1b113c290592fb42857207c5e4ab12a86d3144fcc80df88deae44cc6c3e16eb10e17b173b8aeabc4b1ab06e7eda9750f9c6ef4bbfcd80335a3594496db0e7e8da6a32ca1ef1f4cc68458d8deb05dbf92109b467cf73854e435f5dd87274db0a933ad0f7b6af7056d6b97492f78c690539c8bfe35f292016e614e59ca4339248cbe81804fa1417242eeca468929c5f036905317f17797d3159b5ec3d845bdb8ac197aa14e9e7baf635a708ced035f223cfbce2f342feae5a79f50577214124ebeb03059d87b57ddd612b7efb6e1eab97d47fe57b191c6dfd86008ff429c95d2cbbfb53ee2d32c353aed3a588c257bb841e3008006f42e5fb4085b8374a5aacaebdf1ea4e4386eaa77a0b0d8c54817c4d304f570d49fde93a105deddd31828f985c8eda5e43894385e557be756b891b5e6f3a25069555f44729e76b0ff106ee66e224d71759e110831f9b475d949de2cfb6a33e8dc49c72a6152ba484240cd1326ef1d8d2784b802dae933822e2a3a637841a913f7cd1966a3a7f6d3f92857dd127cd3ffa514f1ea2ca53d151c25928b3983dea50d0af5bfcddac969625bbf54e1d3770c360d436f7166248c975ba0471bf7c00ec8b8ede034eb024cb91972f8903ed877967c3f4115379c46f0de863a5b955a32ac0d339d3bac15eab3c1b6ae9b27754f79a331b22de9c48d6bb60cfc14ab459968fa6b02426ca718f3e6024e54fec8c19c36b693d7ac338866fbd7916cb9fda234bc6c985229e11754565d505901d764b7d7b10489d4e7fcd8817de7dd6e28680072ccc20eec9c4458b84b6e66b7e56e7bdcb64ab4e5ba9f43f4a88fc60982d1ba8dd02ffdb6c5414df6094edc5df58c84d350a3bb54ef3ced2f33b89b3db9a5fabbe3d4b1f2f5b9ec4009b7047223df053462f73d2b8b267b2af7a299519b068646088c96a02c5450dd25abd07e99732e2df49c7280b1ab62c2f94c6704e23c23eb22cfa7ef2de3b5c504d74a07cc4a44f17f80363cd743867283a714d107c9154d2ab256c4f8adbb246ae280e24f2c379b99518dc6ca8a831063d887c1214937a1b2974c600a8f951a5d5948d40f45bbcc19b39b593b5d9769cab74f82396518cc0264f2e0bcd3a1928d76d7b5218c07a9cb340eeeb3b5ada88ff5f573a8560b92cb9f420c65454c9c54d4522477dfdece9e16d4f82fda7bec72c53a12b9df68b04c14627cca84db57cdc34f26c137a7859fa145c37fa389c06bf8f23f20542006ca15edd3343fe1ac45e93392799a8ec262a91c7c0bb1816620e5c8aa294767934e35b2720d380c225295f306dc3830032a2ff80ff6a968cb81e3c49ac0525e3b95ee7b1474e2b5cfbfccaf5437ca9371e26db33a67c275f1c16b8b1a563689ecf1c14b26aecf91a51673c4da721e569ad5cc3cb0ce3dda6ee13a2f1dcaf052b7bc9133e3a678b2acf7ea37aecc72619aadb2623d54aefb8f30f3670f28c006f84889add05b5cea882fb907e5ec692ac89f9b7a5767140f872f11413f078655db181119e21d0c5a4a4c5439ca1c3a5eb6ec5a7d2760105304f9b0b960c6c04aa05a8f1c5f4959bdd4e4e7f688d4b85d8a03c417dc198e27b9db08357addacffabd15dc325933e88871dfe8b0d50633d4f1ae6c0d34a5bb28b13438b9b25df8da6dd39fcf642993c26c370ef2959ffb96b272d6f994e776ebc443b5720542554afc64629caa6140b8caed7b1f536a42ba8245314fe64696aa5a284fc1c7f09d57222c2c93e21c8633bf706988cfc51ed7dc5058b7c709966fb8b83be61774b616f57a79dabe348b4ed61c7a5064a97c5b297fba2884dde4958a4402dad224d16033c2394e892d2efa67ab17283017f0fdc57171c12c756ea1ce351453e008b319e44d1b925901e65d6627174a36c8312bc3e6c270748c4403015be39c05257029dd372f4c6e7cea3b3657a5d19ac667d05e549b04df950c579e3e6544d42930029f8b1fafa6b31879cf698bedeef490ab4cb967b4c8bcc0b7290488a241f61ac49bff2f6abb5fffb19c36145b527000a239b6523c7fea9995a361961f5e1f5f35e3afa968c5da0e3a94d90d0c6e8683f636c766dcadd42fed258d6eb24f4c1b77dfcba0dde7298e052c5db1b954bb58732a9066a345c7fccfe5ea573703faacb238530b8882e68dd77672da027d117717a016d2651c4fd4d62711a209bb5f9f33b7dbe8a2c3338b3843e4d949a635f76ea9d368354c6ae956bb4d93086517a1ed05515800da1761e20dc1c5295447e4b9899bd520ce3697584a7f379c73f65ca6db909abdc12aafa4961897b394486a1d0dd2da94785d015edbb32dfebcf7fd924e21ce263b6f8dd31dc879cd6832da0a5f8102ff26351e72ed9151fd96757b599444f9e4786963f8ed7316b43aadb1c0d7865b0e040d2690e73217acc239630ef890f70d1bdfc215fa464617c33285b132292ec9c6a0c7b57286ae146ee43aa7edfedd363e6cb46541e5c94c1525f885bcbda220d2490f4475f465a12a316ac00fe08130034206f69db5224a740869f913fc5f3c5a47167c30690caaded5c35d6045910e8dfc3dee005b8ba567d38848fa00515e0578317535ac86094cd715bb850cd34fcd27ccdf9671bd6a76801b95377957886058f53a9250137aae9375e0a30c607aa736e4e76ef57c4f7898471647aab526d4b76996e8af0a7d9b7bf9748e0cd31a3efe339a32de9764791390403f78fd744b2de1dfa26830ec7f67670bf109b1eb9cc48a1d28b4f680cacfeea3ffa122a384448213bffb430bd5540e0a6bf80a9b5a669502bc20b254ace8722757ba2de21b5892e779f84ab81badc0e39803aebbf4239f0e67961894b391716488ad108a7a7fb8b2ae614c07e3058ffde73653e51cac97af43cb42dce8b06112952bd69332d7e21a84c86a1459a6f7c78bedf7b10058284efee088a181df1f7f395be6581f30100c7041cb0857e04523c341c3fd922eade775ca9619503b750ab4af837df6ab1ee127a21904490da15688a4b7a49aac274f8f4848ba8f7ffda637525bca7216d64c9ebb814a03816716e76e9212859da2fe07ef2cc0374cfef2f3b5d519ca3a9666d8d8d94270ce617c917570ddf1e3922e9a4b0bb41f1061744a127a628bd48b8297e78161e178d27e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he4a61e12da23f340d938ce8791e0b7557bd2094b87f925322dce8d033185d29535c640bb335edaec4af4246fac547d01f6682970ddde11d2334e1d5ade4d516d85317341fc55a9f23dd3742d0899e3597c74a397271cae06f56f509edbfdd6a2a6147add23bad676a3d0c9a7f80753d6a6c6dbbd850fb02d92763aceee38861db2b39836f0068e17002f4ee985886a6a9368214df8f8626e51bc3d9cfeda88cb123c036d13295a90c2ed2fc0832b8d602abf60056bfbf875fdf48ab5883f04c3713d7e107f52f107411c91f5ef5cd4c1cc6cd508b1ec9d8f13c04afce5b1974d1bb9a1b88cd7711f230c80e4f41ea6c87aed227bd7cfbe7568856f809dd3955ab0e2704ee8ac80ccb7bb06fbb2918cf91862c20cf92e32ddcdde1914bf58236d48e31c53719fc1f1973baa1faa44b81a4612631311ac4a5e0be2e65fbf0959c805d3c132972c32bbbf78342daa88c5d37a4cfa6af4bca27407e1d1dd72d4b8cfeb22fba8b75108519fbad32cfe12ff42f2e4ce42f9f5e0416cb2f9680f509d877b32fb27a3340a1739af25a16f733728b9e3d4711eb0e982da56964a6a0c0e7073ff01457875136e12efd4584fd02a6defa6e142383bbcfa2afeec76dd23156f447db3930ec215ce883945c9a669adb0deeee75b21db91714f0771cb147456e783f11c6cec8019b1cc970aa7cc279d8fc217f1573fc1475cbf5f520157b21ebc5310bdbf772b69fe25d0f6eb8d2bda0f775d69bc387c861652d7832989b5e5750747dc5142a9a8734a6ed546366e623d4615c5175863d7edc69d5416c930f5ed1cdaa44a8c7daefe9c0711d3f211fe36151e74c52f79c4568ae1df8c31ffc155985eb1a2f2f2323a0296ff28857ebc16f63a8b0ee67653f89c145421f56015da390d7e4e59e0b36ec49ef5ce5c80a06ac517f9be302d78a701f1e39c1fd8878534e005fe3fd5e790ab1d9ecd74c8e6faca5814fdc57dbcb609c5f32ff775c9befc7e1457b5d90c30d66b4ef538cf06f80e23cd1787a4967a5cbfc22995f1534ce7da88ab325cabd61fcb3ea52cb9741e0c515e9f0a5a33e2f603cd014c05ec1c9036bdac38e0fdc86b2ef1fae803e1931e8abf42ac416fc50a11b1c3041b99ef1d356f73d9f2ab651ae51d4ded31bc8d9d22bf07e92cf7170e8eac02bc8668c2bf36bbbd40cdf34dd3e5a5cb64e7002937d535af3693e26cae996a1a7ef1df4a66586256745631c397215a317dc127e5cb2717261474f7be1522387aeca91ef3ee5a6e9bed4b70378c5cae75dc4abb672c9a2ec94cd22120b151b8950392f1ea52cf5bf0b87bcab4a734ad37d1720591d8a7a9b9d195547d98d458a6c832ba8575c3d875f709ca630e55e9892c8fefc360bc75598a7437a4595ef1aa95af3341369ba9ba197d1b7e5bf8869dcf029ad2e5c69f16ec0c151f5d6cc46a929227c1c39f20e78647db2879f6e0883a643e3a18c1aae11507cf3a91336fd6d75cce6ca86169ad3bb044498385354b9730165e3b272a8efd0994696fdc58e5d511b8dac2c79ca714a4830c26d49d2722990c355d3a3c2d4f7fe94d30279085f9be0ace8873420a3da8c8410980b9f5816bc460fc119f8550532f3ee6578230e697ce5fc7a7db6f62db408ccf8355590ecb449ff63807216d5ea7843a73d48b8e39d7c18b78933406d94d5916ddfe1e85ad3e8d9f7073c896f30de59914b706b061a9b6b30b689a547ee4e7f61349f2a6a206ad66e47c00a19047dac56e92e0b814d179eabd3706a9238fb5f05c443e770a9fd13054b1e350a57fd058218683a47c4ae72e5bfd2a19ff037459e9df229f947c7d4931bda81b0d49cbb07a5fe4f1bd670187c125f78e86703d425b694023a5c69ce6576148b302ab9b96e09d9ef14c4b96bd103969cc6ddaccf911bc22ef59091f3004212e29e1a682bd4ac6e8e273a8292587e11b2a34832af1aa22f8d22162eee5f42e360cc341e50e3d60a0b1f1753a17198372a061541ceecb2ac398c113fae32e19f722a7f1eb4e7321b6602f984ec6f4840520550f7daddee5d6c514e891670504d3fb33291153d09dae6186359c5266d4c2873ce0fc84e1edfdfc0fe30753e307e5885dab3736e4c47033b9dc405a6aca7910efbec301486b045f43d0fcfef34e43a4e03fe5d2cca67026cf084c3b65c9e1af74a8186d81cd8fbed42cb9445e5f4daa1826c0a8b5d0fbb7ee4ed09f3c8e385020a07560ece07fc254d38c7510cc4de370cdc40dfeeff9ccc53e77be3be886df062362ac2c61a5828cf59d1e97aaad7215ad4c29915f51019d0f8795d0ef55c443285d16a568709f9d49c0dceee54e6582a4cb36620afec9913a57e639316f50d9dce9accc960bf0c14725df19d4d3e46a3626ded1c7c599e809d9a9651bca98ae00cec8b3c47f06c3ac7ee62b34d2987a51bdbd111020f9dbd5336579066cab4538531d31b5934ff244db564778956e2f5ebd9478b8d454425b05b477081453b2fac6ca8b9585726d11d6ce9ff2925afa6da3d7d7b6d67f237bc84fa9b6a74901afa18cdf38726b1b2c249d81cd5c290baad441d367aaed998c2f61423dc9a3096603dd10d0c71e3514d2027a6cd39658d93ebe0d5e1a38cd5a20ef6060ecac5731f29680fea7a142d347018e399446a8e4e1c8e2bdf81a1ef36bf8a0ebbdddd5c5e3ef8d4a5fae52cc1afffda9ebfa70e8bb1ed5d55f3c6af43a0c9425c303586d4e80b0b4c33cb85c801307a5cc56811cdcc9e4f90e0d5b702d9e564a36491fb455fb87a6a66894f4447a8e0b4f101a671a0eee1e70ddc83907ae47a7bff8b97e2ee2da86d94c5a0d30ede3457a3ccb3bf23b9ed76c671d73f82626e203e2e4d2bfb6bc96aabfe9e7b8804042687243d08a6bb57f1917f76760c430df49f74e85c0957d6cd9c1df259c0c0bb2cfab1ccf0e02a9fb10afa4c373037db8ef9821c6e07b956ceec7b5e28892ec2aecbd7b6ab67ddb26bb9f6d43396498785a5a2094c9a0b5c998ba734d41a460caa5ceb4b8a285195c2cf6cafbba2f7a0d364618dc81b45e79f28d84ef445e84597e353fc43fa2630905ba01a03b1da34ba56e6b071f20d2e3da6563ed3fdb71fa4cc3459598636448a1e91c112658990afd31b26b60f9bdb83ee1b2a9f1fba2edc3e34081b3063724ad5e6419f6bb9f761cf615665a8bfea350ad47936684c5eab4d343600337f3847eb283991a4dd878851cad92a2b2e40a2fe4e6122bb49b0288e36e1567089fa3825a598e7c878bdc64f761ce7990af06636212453859d64dc4359ec7e85bcb92d32ffd39b84290973cd8d163b37de10e06d78399ddf2c48876084fa4b4a35fa4e129723db3206f3971652da8101a398041c03fc21687033ffce7c66bdab311bf360a5e9fdd5e2755d2834bdf0c546b51a1c5e3edca067ac64d7907ad04c3f50239bfd6aca1bf046d7a99fda89aee614c06ce099ea88b00d90c078d0b48a19de0e18358fda805e8e24833048fe0a9011d734c2f281886b8ff96bf02b3c6e40834f552b708312d260b9585be8e4720dd8cfc72c283c12945f5dd4f140c71bb7c904292ce5fbd59dbcdb2eec85ca7441520182994b2b03fbc0bbc07a7e5386f908333e5725e148e94a694ee9de4f5cdd8bc721620935a84351c258ae340631cc3be5f6ba4c76e1f068dbefed4093896a1bae5bc052452ac9820684afe52f928698d44fc90edc4ebaf27f7882e51ab6b2489edba01fad89411185c7b7a8af3f4fa4883163c1deea257263dc11a6bf59a87435059de8b8d58b09216c81c3c5c6f1e4668cbd754ffacc51051a9019f13666f07bc3a107af38fca012511b4d63089d1da8ebda8c1b27663d3ceb9f4a274ae1b62c0b54ce2b508a0c02835a12e4d15c0dc4d0a3b8caa11354c5c4b8dffee0c0dde05dcbfef8a7cc51dc97b365bd54f7deffb0e40290b9d3ad559cba9f57b2ebcc43f370f5a302e2595c168f2eb03ba2852f3a2053507d99bf9e7cdcf717b94d676209897733c6441ce758fec104bfa2036bc79d26b13546eb56f6612ff601dba6ef4dca396af4f9ba1f5a4612c8655b830f9100ce877d4a676462c9563b20aafd525fd5f9e18ff4f4281faf478283bed1623bb9ca16a47b973203e92185593487fbf90ff146221ff184c4b9b75c98072c28daa6ea8028f6c84f8857d0ea4fbc516c296fa74145ca36f40e56ca493cb43a392e6657d66cd75e1fa59fd50c2aabd987cb52aef71ff1ed865596ec7ff27329c8e80d04bc49d1285d589d1155c612f65141d28a6054b433b20b555fc3ce74a13a025b25145e4445a15dd1cf4d5af551eac93993db97a44b7cd6365d35c34e27bf07275f9ff65d2bf1e5f839a046b839484c2c439fa38a8c3fc58445189444725683951d5754dfa148c4edd91176299eea17751882add78d77674c6fee0c66b24c1f6125a86b301b2d9f4c3876e018560cb20c38f90a05e2ab2983a90b5a58a6a8de420d6240eb619f4962fd6bc67767dc04c618f51f6fbaaee0c6fb160a14b1cc8ea34d7f3ffc76d6d29af3da6d95114bb50040eec75de5413f2d40cb1b4831060e0729f7ae7e7800337dbfc8f0373c1e25b980596453673e6d22d7da58a1207ce848f54cad4627553f2961eac82c695f47503f047152ead4671def6a1542a72ff79b9658eae63ca9b45881a4d3c163cdd71dcf0e20ea5cd751d71de1af4b08c478cec15860a5f6463cbc19af82dd2bb52117340d1a549fdd09e61ea3568a7e7199525a240d9358e8bd015bede8d0fe6ae6786f13f49e057a43ad55c92ba33a8a7aa9be56b018ef8c2292dc2b0a7cdf5a57a159948c30f75ca1206d3132d9c2f7d05aca153d86627c4794ddfe47beece5345b0e679e47104574a85c95acedd7db89fc32a4667aeb454e98bb45ee31dad9428fcc299a942609ad16b961e3fc531ce7b3768fa2926ceb1c114fccdfa2552eb6a3900138699a941ae261c497f0fbad71a502bc87c90184c6107fe5331612bf07e9869e1ffcba8c372962c27108a3b5b4038f8345243009053484b3fd954b366cfbc550a6278d7940a98160374760bffa2bc1fdc808a107fb24d3e3703a0c14adba58fc3c3fe0a4e57bc72fbf24183d8e1f25bc7323795aa6d8b9cee92148e0ad176cbf7705d5d484030a5e15bfd128672490bc9f0f4ff416cd80ec58d6349766f1e6dbe56807f66d11a3a396d1d57cf1dd3aa7947d14f970da9be691da1832df648aeff8916118eb98d69f5441242321ae32ba13cfcea3480504474951f098aac0a3ef21251e72bc42337e23e6941292fd863fd478a86b5513baf7dc24a9e1ce316975fbe685173699f087b2aa86b149fbe795926c38186774b37e315e0f2b8ed6850439afad299da318e73cd2c51269ead969fc59b03896900c9b807c5065b82703ff8c86f2dda4407af72664f9f470822272fb2c55987e6d6c6cce40ce707148f2509a1ab2ff999686d3cfd7e930a239fe6b652a7d1bb9af66a60283cc51bd6df0bf56190d6d18740e9dfd3c2c8ec5d4ba94276ca63d84e023dee9f0c4c874b38cf3830e3481e85acc731cc43aa661b2e344097cd692ccd00e1cdb68064e5b51201be994e58bc9eadb5bafd0d5ba6be776a0a78b52bb2b4e299f7ff3a52a3d1adfb44e99c348297e8da55bdc6f5487c65ad29d7370788aa0d09a5c7553284b44280d4808eea6ea2c351efed0f5592490db77490445d034cba88b5f87a409818aa6371d9859808a1d0a89aa2869891f767f89069776cc4b20dc5950fc3342c46cb9b194a3e5a95596958945efd0d24cc2e7af9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h2354716baf6a7a85b5bfc5da6e9689a60613cc5b4433a6ac433bc553d97f177fb2c2368527d2074f4eff89c761edab986c26b291bef5ec418033895b99062ed867e20a0032e5c9215cbbf2577cf83f964c46556680b0db1725d995f27369d7eedcac59d60df83c85187f1ce41f12782a17df7ef25f95165bdfbe3486936edd3198262e6bf6f83658a7d4b99e6e64656082a82301efcdffb8c4fc1763f2748c6513de6c4b4954b92a76d162a9a3df07f9f8cd9e1636877dc06ab6e0612970ba2427e08f2d7d07fa70d93d3b58be0458317d7d024c962f1d0c58f73fea5aa45dcd7a14dd05f026adaed32cd788d0f88273ef286da4e35a2a8a515933301828bbaf4cca1b4e5cf44c29fbc0a62a73ef973fafe9c1bb4ff5ce69ab7163809322193099996353b8c043dadb6ab4a1648152cc29a75c24a12f2ad660bae6f794f3aeddce43366b320631873f95ddbff227da29452219b6236b8c466c66802dd11a122a3cfa7346dc9eeaff6cb325f6a2ecb06bb3039ee7ee47808c4e6d4500157419c30c74cdc430571d58d9df9c36a5bf072b06b981d981cc4a2a4b68a71a7556a0130d6bb2f058dbe18c4da09c087339fada45bfff96d18548b57abb9a72a9de27dde5cbffaae27f906b13b40e0e389205562f7645fe58e9142e995845a84912af883592904593862de477400a4b4d0b38eeac16efe7a02e228b2542462136f9f9a8f81c68544f08c33766622ac0c0930d50d770aa57fa0ddd6868cb3fd99e0bbe3fbacb38ec9f7455b3b5e9ec88c308fb3b1bed758b2872eeb716017c2b08f784f6441f0166c6cc5c83d52d0186cd8d5092bd4b24b10ebd290d0b499eca8c417f07882b27065ea104937617d84ba38ad4de49ff8633d03525cef3cde384a121912cb9271577a291c95a3be312ca95c65f3b445ab7e94a922a516b2281072a82be96720bd356842c3c9384259dbed986e5d3504026dd2618742d25f5cb4b599284d076d0c20aa51a6b8cfe3a8f1047b90bc2fc33f66d8fefe4dcbd979e2d1d1fe9dea76cc1d56c45d353671d6cdaabfaa096302b06af208b36501e36fbd9adb5bad827bcc707dd2497b5d974ca31d0d38b6df4c93f664531d59e8d6b40096fcd74b4fea38f7572736bed7a724852bd1dd5ce8b00923dd8954786142afed58ede852d7d074ab7acb22b06c5e2ccdc4b2739bff941d2009e9e723f5ecab65a0d4a10b592da57df099a363b9bb6868b76c7b0b437abac6fa4f01258312edd0674011aafd4a77e1db92a4dcc5516e574c2b31f6926604a600226587987140fa9ce7fd31d9d23a2e44ad30fd4a9bf3c6c2a113a12947ff9671cbe6b44c4c0d30a72036b17232546dbb9f42a58e187f21fd68c5bd3e28dc5edd67a721184d49c60ab843812f8bac4060845c2bcd77b1249ad32881117256ef6e502d929007903d8510e3e087bbe0c3125bf896c670c3ca054a67249f1bd2dc30d9d2c585b4838d0dc4d0201d4ad04c4ea78ead6be2238795dbf309816b5a3e7e205a9089b88419400255ceb0f579310bdc962895ba48567b94c7c23311c0fc1db946a65cc74a9d15c7499d747a639034c3aa4ca74fbc8c8282171bff8e1d747d5a743aee129116ccfc86be72472cbd805a570167276178735a8611d7d8c64746b74ca542928f0ec5175694093619bd165c1c168b92cc9391e3fc2823e05e2a24f0dfb42e6f3609f6f06ecbbcc856916bedf23cb2d5b198ca848f0d81fe11a7a09d564c7110456487576d07f51453156ea6c585e812a67f05421ffec300f3b6318b6fae016909d638686bf14d8e2fce35a86d379eef5f24093ed6ce7c4f7c5b7ecc80d415f7801507932664aaaee7f0503c386e3a0b3dfc64fa05a9f86d0c80819590dcbfeb60b1ebfb66f16d46e6cc9ca27f494a46722dea83bf6ca40905ff5fd2d40c26c6e115fc1c6d46cb9494c5d227e5e16cb0f3c0a5f8a0b30b25829a68475ace5107a9334e30e8bc35ba31f2dbef68c22536fcd44c951a4d159163c9a11aa56bb9814814fb8ce02d2be6455c03651b90749b6ffb69d6443b4e3c717ee247342c98e6374ee4d01896ba27b1c6170f6a936e90d5c1e963f95be7cae11f5da1598039e5d06262c07cf9e728b7a7764f6642253d93af433d41f0470373c9021b9605c051a5e9b807e694834b7de11116879aad5b7ac42924e0db4ec1040f3369d4e5eb83404719eb79c3d43fab35c2425d87c723bc0328f734baba5859698dacb94fe6b7624d79b9810157766bf747b8037f11d15452a04dfe8cfcd15fc6ee618ffd6b0fec0cef1f4163bbfeaf107a08968166a90d2feac3de98e5e1528eede5a6f798bb5a775bb18a3e65050a0502c627753a21107ca4a3fef3329892d06cf1802f9e97ef676e7878902dba839d4b422cd3431bc7e85694ee10da7f2f1911c582c7260f29b5a7957360687489b8116208180f967e9f5a3f3b3e4dcadfdcdf4a0451d5e3cab7704c8d3ea820807fd5759526050b067fbef9fe06e0d62ada7a196685e433d3d3470dcf91021c23fb45ca7a9dc8301de404029bf94bbdc148955630e6295b6babf403583b32306aa220bafc48bba36fe06d79c74562ccb257698e64f42e58e627e7857ef5a1cb4e016dcfc8dc8d0c76583d7d19b9b9dac8cc208ed7a0fbab3b31bb95a6303ab132312f9882fab83078e3738cf0c8f19f02c6d935379107f0da219036e4a526df1850d2f888b42ca629411a7670c5f166de11b9c82223af993f12cf21a94c5e0b5325b8ce199c156cbab97cc3c1f90af929b542fe0075d677fc0ddb6ca172b00b802fd03ebb294770a60c3bb188029d5a11ba4627e3b3286bf59d90c312e1d87ab8c9a679a47538766d2cec219fa6ccb63580b0112549121ce38faba0a4c4f2988b160582920a68b9d4bceb9a00a159396b620991cf3e2a61eae31d9ebd6eefc5583d54e33e2e9ecbd046081e067621adfca49819b08f19193cc4556054363b1735db960ee7ead84703003920c19d4131be8af5d84d16131f65a54d786b6738dc9840abf021b76e95d589e475a5f1ea5e3b9ad0cf1a5fa3f66eb4e8ddb8f84a0bb30cf73325cb2d0d2ac4c27ace27187060f1a856a9f14742a50e91ee873f56771e863399e5e8c149490798e30388399ae1304ed456dee7acb273e473e398b72ecdee4eea15c9dea40596a17e1ffbd133771ac0964cfad379c66644f8e551ea0edf0a46a63daecd93ac038f0c7debc65deedff0b6aa034bfb540165ccb3dbd279277df8461694e0d0bbf0d3b82148d8f3d6c6e412ba0aeeff1a5de7ba38d12e4559c1cdfc673cccd98e6a588fd07a84a6c7b02f769ef289d5d80f467e27cf8a2b686c3010ae5d5b60b118561560f76a839a7d061d4411e414646e7d305adee811fc6313a4c0b1d5e47b4fa756f51a1e58e089e4fabdd53203b6f4aa7a409802f783496ffdaa19b69d5b9636908935437e2ede91ce13be71ab6f4a9b3df337de8b96aee69e21d51cc14afcf5d0bdb2c910671e0eac88b5b5b2f80ea1fe3339c0131651114d3a43faeffb8e0d260b722805c4c8ebd0dc7383ad1a0e11f0471875bd9f07054656abe7d31866c4c364781f64cafddf30e77b5717699013a131e0677f2be50fff18891e2c17acb97c00c799121d6fc89175004c7c3cbb62979319fc2ae59a2a2894f078309938117aced77d9f1132edeaa38ecfe1d8f951476d9193c33120a43b73ec45531ac28a8327effa4e56271c37dccf7d615f216d05861017ae1d640497a3ce4f3a2d4186627a38619816728da49eb7d02cab5dfabdda23c18d1f85a1f80b7cee06ef9f0f928236a709ed5fdd14d9b75ac5ee7205699d6c8cab21b9d7ee4d7a2bdde9933aefdaf5af64d04a357874341ebb00f81393e4dd821b5a878625d38a30bfc82bac1c625da3563b271076163d18f531c412be6519aa8076212caa01d5c153a6bd0e7b1c882a44a3246033bc484a6cfa044117468adbeaeeea394f9a46f5dbf57bc8c4613ba695421703ae58cdac1f54243a0bf9d96bee821582c3e7f32273a9ae0a36ce3ff1b7827d359e290ed85220b1c9e10089c62b790a272ce75458d07fbc622506a65e3a22426a9437d64c2616ed33a8cc50aaae77727aa7b5ae5278d8f2cd2d209220bf04af0e5f8fd7df8eadbe0275b46fd8adc2eeeed58bb030c1d50f950f8195182fe7b8923ba91815b9bf16df5f34d9a21dfc20e96e9f27c46628906c7063c843a6daa835ee447f7e9846873866e11243f53d18065cbb073a15126a962a4776ede26d5fe0d8e3a01b10ca60e79acc80d2eb2404e4c10c7d8261d3b18c43738bb0de49043a6eb10fa0a97510806d6728795ba08b2e3bfc7f827e0cdf9a8c1cc49b1ba4780138d456ccd90464e62664ce282b986706dd2db9fc5c117b2cd3e716a409beed843a956650c25eb8c0de9ddda68dfa72523d19f714811e37bc5f783b067f49f40d4501ae1ffeb07fd79e0112d8044e6c026564fe2a32e2829961d74e8bbfb9273f4ae2bf71791ff5278383003fb9b44a5cbc976fcd37780e67d9a193bbab3a40b84b6d8c669b81469b85c708896ae01ea10a8adce013d8cbc3ff301f6e5b51f0109c0fa5da6e32fcf48c1478ba6b4dd8e6d0f52e56cddeec4932f72a55a2f69d2b00dc1dd0b2a1011a708bdc40e9c268c199934a02187f32d1cf19c605c5c13e43315c378d7b786927c540b5b81337d55605102b7509ad2a82e2afe1b8e69c6c6b9eadb541184f40113ebb5bbde14c3d2941a5faf081c9a69624f50c44ed7c967b48d29401b483c1e463772d95d073fa248554f03f21eac3bdaf9d4b397a3424fbc5bf78f33d986f77a106c2cf6007bc8dd7dd23d9f7798d837e6e416ae556d3500039b0809cb8c2b0715383f0689d63b69bb34fa4ccdb7bde3e6a0dcb5fd0b5f3881cf998654bb8cd93c34f5604775697f555be11e5f5a8ae203aa7eae9ecf97d5e15135579fcee22a7d5f3c6c52d1121b07dc20d1e02f3b37a115361af8852c357e3c3bf48f98cc0e812ad2e9b8039e1d7302e743359c27d09e3d92db822947a938fb6dc25b73c2d2a462fd93325123a017ebc2f9230bd670fc5211475f02b69be234980adca08c26a8aeb9d0651db62311a9829177ebb34132d63b599bcc6d0dadd5edbfd6750cb11dd8b4e65944e2c9b8d703adddbdf5fa1d0a00494d6053e0e46cbff075892bdb1636f0218da0bc50bbea651f87162bce466600e64a08c8b7de631c38ae40f21436abcd3f9e3dde97f55649b20c355623cb24d2ef9011e2d9a6c09616fd31e804809dbe002ff4aa302cd5e09c18c8e0880ce4b5fd94bcafddd9bf850270440692cbc4a2dc04011441c8cc1469e3099519ef46f156dc31bd83af2e32587796a9e36894b803a71e11d5eac5c3fa8fc7c74736092e976974dff43c1803cfab97fb23ad5cc5280d147a127658696bb9b7e19cc77efb1a50392aad1b8fa7c6919de0741f9e826fa1deea68ca82ee9fc268a27b2b19a7dbcaf1673fc8aa981ec0d2af114e8b82efadd9166526303e602549d5be9bfcec966071bac657047b798fcea691df32f8e296eba22e16dc56a09a8728ead4358b8921d2bf2f730f9fd48a32694b91eece286e2ab1a7c4651c06e2ac2446342c7cd84457f1003f90e3a6a416c0eed1a77847a66a2d11fc9d9b126adc7164d18b4e8dd8f70337265dbabe405980a160b68df12605197e3ec77cec232ecf72662d6360c487c2cb08b96805db7650586d621101a4ba53d4123eae1938cbf154511b2e55610a7a2468d58a07a7e2b10fbed240;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcd82c9a975507b66b1667046746be3bf84e083f0b01fad97f0c403a5577fef8a7744b6c1b0db2ebcf187fafc40a85047d2165d08ecd77ca045a732d96e42c3651a402607961fb6c5644df19cfc13c77afaa81645d7826158c04a5ef4ed227694df9fcb5f44bfc8c4888bbc851f74fc6f28deea6491224fa9e11563e2229c32549ed08de1e2a043379b9581a9e420f80663a5586308914555809f5c3616ee6d13ad6a53cec34b7831e3ae059968f9115dd653148c750de79888072561ea9c02b4d30209def6623e25166daab81e4224bd6a515d4bff6ceb7d44f467c463f6bf06d5046ab6bc493a3394c130a0ff1769d4981552005778245482ce4b509712197cef47db2b72aefd0c7a4f386873d1c6584fa6fe80cef8d683a909e55587e404ac5ed080f709df613ff811e30b61626402127f99a1a897e6303795bc4600da6445104bc8b8d8ce8e1fd01ccee59cf9dfdb3d70ca9d450c817313aac89ac0df4fe6b2808270a1512a3a91039f2ddb8cf62413d3d109d2203838b0e0b1d9be46f348be29e6cdea02ba46dc308323d8c57092feedc6a783007dec320d01d2449e734e064bb5e6fac094d4558b6d1b9df09dd060b71ab47b2d24079e864e1653563916e5f2cb059cbf71ca9c1d0cf598231b707d513a3a040124d28df0666382ce0498c9e704f34ade9434478a6bad3f46e3658c04458799e1173f974ed173b32246bea58e2856598d577af78b7d6f5a6c1ae1ebf4d7afa0fdabf5269712abdff85bca11818aec808ba3ea2bc6e41ea8aa0cea5c07c87c403db5b2597c30d884be2e03f750a0f15ab6c8cb98675fa6a05fad20d215c6691e63c2691af57bf42eeeabb42df4c8344083175c6678fd8ec6af71d491943f296c0ffade2f97637f3b78a2dd47be18da2e9050c996bd349ca62be85c8b6d02009607ea067656c3effd512182cc4a42c3de502fb813e60e673a2ec796cd1f19e3898aee6ea9d05996684cc561e6e109c44a16e24e39c8073985adb3b0833e0c73f6d752bed1d81def2ccdc9b62e36750f57950c3ba0c264d8c036e7ab7984eefbdf4214348129749f7e0092b71a5d546e7762af80f68c181bd0b79974a713b787c67c8e62e9e09d7c45d03103531a04ee5e7b35d7587500d9d89c1c976504ec3e5a613ea13e84b1a2895e90c1e770e07bbd5976d79bcdac4f35d6896f5b6d587066b426a451f54dd7eae91b0c7c3efe3e90b219914d1b45fbbede6c85bead13a4edf8d79a8b79937de50241e42da591eccba55e9d254b4122f7cb792e171d88227c29601343a179d33b52e8e35a474e8aa4a16ec4a94bc2053bcfb5228a882247020582db17d478e103ec5c5855310fa7da1b079d991cf78ba5e24e43df5a39ea340cfedb0b3ecca0be14e802edb6eb818a2dc3984ed1c17fbf16adcba393271ca4c88b62f3b09c01bf0206696e52af0cfb9fd483101a02dea20c1a7201b691a1d77ab03e80fe7ec893839e21e5e85a7f720e63c4d10fc3ee361c62300f5a68e172ed40061227fccca659f774de9b6a1ac4e9a96b1e573b22dd4b4f3ea48c546a35faa9e1c9f3e469cd8e6fbb947356f6fd4091348dd014c6d63cea12fdd6a4a9c58a78287e8ef89c6f50819749c1f0ebf3c7a2b8370557b08245980717c5d599cb48232fcca3c4392827427bc154f4b6cff28a71133ab420225d0090cb3c68d6494f5da4bfc1656cae1cb9e398ac412a8da8589ec868551159499fd94873536c0a23a51dbc9a92291fe10a31ccb680077c725ff8b2bc10a987fcfaf1244e29a6952f3047828301286001a5f9651f15bb19f5b059739ccfbad42c40fa159a34189bf90b9ac1ccbbbde27d976e30379e80dd34d8038d37e63efb0835d2cb3f60738fffa6389a0236744c6c348fe9f583c6aa707438cf09730bff35cac1e24716cea7b7405871d082d6440573535443efa9ed854cbd816caf584507c8c93577f647008cde9773c34d3a57914bc04c59e543d2c0347017d64458b8f3f6f3111d71494ec8591fca4097a968379acf9436ebaa9b5f151a52a01f20fd38c7b9703ad75625034705fa8c190afc3f4dd8e21c9f97c89627de9cd1cbdab95960fb884ee8bbabc332d7644ad7711bd1f0966e21cc5f21bf8e725ab12bd2b7866f7e57d40d55cd0717793c219044a7467a221cac2dc1624f0af333176d7e345777693b77a0ea97117413b389a0f8ccc42af855dd46fa0d80f5ff228bde64154d2a3d5ed03141c711dfda1ca0601e774dcf0dcd79ab0082a34d4fb6b2f75728d97db99bc0a0cdb2dc66809a3adc487e85d0c05f7f37cdd7536cf9d489e7b2573d683dda0f0bf813787977e249c45ac727de6f0378c8e32bf5bf1a231a303a1dc571924134098e892f9498e1c58e78fc4d349e0298effdd397203a43f1ceaf4a8cbdaca4065eee3adac0d9e03e8af169f5235efc03d79b96cbd701a78b7b5d5ad4a732b99bd6479c9f2bee2048e0ab523db31ec5c553bf8f340311f920873e9628e373a99f516d006736c00c280253dfe4af6be1155f8ac9a5f3ccaecfcbb020fbbeb251dd00b3b1ead92e9217a2fa5891f55dbabd0994066e82ba24a7d1a478bc5d9ea467a8942a09a14b50cae1b32bcaa69d31afb601e95fcdfc625fdd1a73b380aa83b9443d7be851850d15d27d2d401c8f42d18643ea5fde674d397db34438e912f2004a776ea3549620987552ad529dd4bf47eb74bba9ec36339492eaaee869b8d7ded91bd002f2a4b0c05c6bd38fed1284311e7f26fcdd531bb223a5cf0fa201d32380740c0896aeec32eaebce561e52286a755709ccce066eaec22d3d479bc9fe6ca7b677e6437986d1ad2d836c38c4022246277510875d07a28139e25985e6414e762e146287956fbf14bd08c4d0211cf96f800c61ac9549df2ad30e43f48b42bdadab25752dc302f7b348914f755b8bc6d04815222444c67b50d121a04a1378963737a1c544aa5e1a18519387f0b0ed356bd739ca0f43aa7c9ff2f1bf2845465e4c901a785729acd454bdb26b3424e49ef3033670269e3b64475f664295865664195de86d147d798ee7602c3b9168272bf7f1ce7d9fce0fd2d3c68202084eb484dde6d33d66e55e8d95d235ad7d526403b0e5874580149d7d22ebf3794fe25557906e5a89a772f71b709b6b9ff8aa5afe77ecc03ad78874ec78f6eeb8aacf7b11e3846d83a77b3508f94b05a84eea69ff7ba881adce5d0d1d5e07e45b3e010246c9d909fc3ea57c8f7f98c7ba069740d40364cbbc3deff4702cfffd04b1ee74534da33b108515a21860d97a210e1ee9f92c0d7d895accb05d27e81726e87f3500ae6a584617b08e113fc75cd78a2f0b199761bd723c8d23b0c9c5dc4c4b9c857858cb7aa27158a9cc2a7d964d45c78adb63b0d3cbbee4101a781acf16967d33ac523b3b87c1f864abc740e8b70186354f37ac1f80fa750ae3d45a6c071e7fec3274bf4a87a1a305916a5084db030b4c43eccd1e9e1e70ae0c3614ea140d73ee0b95d77d64254859464237a1d0a64d6cdefc0bb6ac69a7168fb01e5eeee545ebd8e1f3b301c7a2c93a14cb2ac66a33bc28c0d4ee92f12afce7dfd8b29e6c7ac2d6f04900416d5506c7c9d01dbb43a4a2760b727cf7990193eed9588be6f73a788a2599950b4ba893618977b5c3018eb168706fce975ad9a0b1260046a778dc20ce2c5324404a85b4019dc4891ed09d05df06d1f4f2d0e57b65582b19045ac47996268dcf606774daf0ea24e16ab59dfb52a9fd808fcbae6a28bd543f7f0a2b303cc2d24b499d3180d2897c9623be7f5f1f793c2cd5c75e1cbcb64c3f2cba44d9e053f3eb52f17c2281e1b3058808a528400df9de6b373d315d448ace0ace1dccb3048f9a2967de67c69de2ccaf88e07a2836145e687b17f21c5e7c87a9f05d50368d30152b11ec36371dfbc8a82f30d8d1f6853cb1d2dce787f5ff7edc5b8265075fe83ef94891118f198050d03ff7b0b0e5066cb852c00acc63e6e2c8c3b1904a782631f58555c454e5bb1dd236498e275ead4a0accd2fea136b76123abd2699531ee5b7d6346fd57c34e067dcaf3a75df2a7db0dcf55d76c251223f8cca5e75ce407967a19b39b39727b6fa305a19a246c2ae7937819a32e47681ab9a6266cc48d4d9e4ada353023bf8e781ae1eca8ce61473ec648be133efae95607c06b574f40057c4839158bce3fb03ce7d3bcc2aad29809e7308f8361202465afa9bda0d0d7823d39878e600614b76aa5535dc061a82577314a9fe35cca42e0f2739d86f93177fe722d1af0884b5a237f7cbb0c2202a953429c97c827ba492fbc99a8efce17a9910f59a8d45a5300c55f1ec6defad42229c332538b7ae4f7fe35df037b317b93cae59490bb2be528df40856ff551b97ed9f39eadac7c45ebc07a9a608d95068ace8e3cd6fb871d101c994ba7bf42fc774d58721fe5fb09741b3066691208558575fb4ea71312e7760294865a15e821c8e47c130c06b7f67a4b8b981633b0f6c901d5deed1324065a35a6f10ef43d41711024faf1d6c27c0bf29ba29db52f49eb7e812ddb0608b029594660b133d0643fbf73ef4de48005fccab95744bc2ec22b5a2c857da1df08e12cad3a0c4f535f630599cc31764318a2e950b85af69a3e6b40a64f8cb1d093ae62cbc5fc884b484ddfc1ad276c0b619eb6ebed022f972820196d4ca9baf0247c5328e48a491292964631ec6620daf2709d78ac397824e6068147c32ff2c3cdb1b8f3ca3ef4dc83d814d8a5fea09524e0638c2bcad1558982983da79107be70b25814c796e2271a7b3cc0366be63b9f4977973bceb69ddc7189e1ec4c4d37b72a994fd8956f097681cd6d4df5dda998d98f18934071245ca8fb7e7333f7692586cf3a7487e15c5b46f47f33792f49e45553f6443b8b00439e46db3c9b4c8258c733dbce848da88f3054315fe6047785688a184be4980df9fa719269064c4bde5e58a8028c398a8bf38a2dda736a71565ac949783b1035622b216ce47e4f8cc7e0c17d96d1ea85d6d6571933d78c8e6c90ecab255850c9c040ae5510e6961d285ce70ee819da164efc9180538f0d36f8b444a689046f91ef05749e8d3f6e36490d831f2772bac127034a8fc3dd692e93c60e285893f161eca30f8c2006c9ed14b5fd509454a0bfc427334a9a0cec41adc5a7554b15a7daccece22c6ea29e54ccef85b1b45c53f04dd19c7b2e74bd3d93fc34d83a34bc7cf8c5237dd596629fbca6a8d867e1381a30e074bfabc597dd4a708b3e5bd2f4ced7d0c50d945927d04a6ac53714a7fccfe4608cf267fc9c48ea8928592c31050c073e91d20554fbebcdfe68fb03c8f224d2ce297698a0cec03fa3864b038ed7c65ee0c1ecef6d9a46d089829ab156f7c17b881a7daf4bf1fe79e5fb464da149774bf4a7a0d69e133b3aee66b49219eb44fe0a12332fa9d90dd65a4987e94d33751d0a353d1ff52f466774971b749a8ae3cf90818d1e50a4048bf58d1d58008c92bafd22e47facebb385f0b023446eb5e47e97d336bb26ee878a8190a7148b986845276d21c9e7f45992ed4437a5bde06d7ad55f40aa0327d0138fed8cd56623675d1d31d41c044b218f344b6fbee59051f5db664e66bc81fc9e39d92b9bb2941755548496584eb92e2325be90207a331c974e3fdf08b8bd9f678d16dfab33c5a12c74cc09cc221468fdaa8c72ecb52c3ce3284bed8e8955907f7556030715199f5073ed503adde46d08b4b5cf7d96b9185553bf29a5e50dcd9e709a8adc29558c2527f96642ac82956ef1c6b927fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7821ae099bcc28cb91db3a1f72cadb196d9fb8f01895893e89dfc355b57fe3e8a864f5585e8cad2a468a115286a7294acb76b301d2bf5b69fb9f5baaf713c6821e24a795bd1e35af15e309c8f4369093b7a4f46fc920b26c733b078a0b7647a37ea1c4261e8f9e7aa87a5fb2fa9bbf5f8c7eed2dfae1bf7fd26f750c34357273740c6ab35b56e6642ae4075371421688b329336fc5f4bd06ded737682838536786a979495d26161a193e5c73b596a0e6e5f7cc3f44e0584598950f97d9889eab56bbe19e1ae11acd17cb0e405adfb719bdde40811005159910ceb98ce001ba9af8e380c134ebbd8b957fc418d25fbd8987a32451f884efcd8a0a068413b7fd4d5b9afc8ce19ab6213d127e692e56b80cad1e408f7ae005af4393ec85bc956b6f6a655f12e2b463ff9d1ad49703afe24c5f3fb5f67ef6adc4fd16edf3bfc4b6854b611d27cecce423ebfcd12b668c7eb1ed406e40dafbc940ab26ac0ea5c62e21ecc4c1710d38facb6a12a0836224c8dadf432c27b736191caa5bdde50d051ef983da573689a0287e3eef1364c35e585da7ebc3bc709e9ad5bd131618ab0b6247b5f8d0aa1cfd48fa82d982bf1f1e4c243a7a496a3250e10475759de7e2bd17cdd286adb5380b8281bca9045bcab56ad778f01f645c0462bf3fad07dabf07de586caf079a55c7f45cc61e04c1a7663c0ec940f32ffb44bf77f0d3b56299cd192fcc07b7260eebfc89dfc67d1ada75129b227cd8ab2289f88887d8ed4768a2779a58326a2e9181d204f299fb9a7f61073fcc9a6a09376aa38d49f3c952f7bf91d2b767bebd374671d2627d758f0497c75405ed5ecc70a255f11c8d4aa2a49e6fcbc1c24bd498719252e327529cb592abbd829a591435125bbb2c2d2e1599036c26a81c063eec224c4d5eed952ad3488468da3373078566bcdb29e1a8214f5a8300597b742891fe3417c0d4da42351af10bb07203241af2730f62a350c0127c69e7b63b0bb297da3be6144b32a2706bb47acdc16b20998a27db537b22588075c228872052a1f9fb28f7c8d82c6c1afec9162d97e9a9045460f2b43b50a374d3f78431ef3a5aec97999a150df779090f855fffed444dea8fdc8d2f4df2703b279eebf28ceb6ee7d47eac70cbd299fb30b819041a270d3faaad2e62b01856bdb9810da140c99637c7b4de92449d60a5fb78b9f9cf2e61af2fd977fc2d5828bf822ecf75c0c9147b90330e29e4ea89d6eceea2e22df3ea13578e6f0e4e47b26f0ed4ef92c9380e1cb2347696c806b8c82ecd2b7c2914048d8069750b89dab24d0c44275ab09b83fd05dac7314dd50b7d20d7a7a4d1527ef82410cb9c1500b4e06a8483f75278e63a556f153d04d5def21b8486c2becef25b0f2597c1e2da8739cce2022e62daddc79cdd0d86968783f501fdbabf526989d25822914b0815feddbe9ddc5c9173e12bc568adb360dbca93ecef3fe8310eedfaea2b2c1d8f8251f6de41d8cdd2d4a71c5627dd235e647b2be99c6a87d53e11e4d6535bdc4f26c965b0d2771bf63c27474ee98f80b13f65bce8729c4f96e8a7bb0b0ca54a844832cf8dcd7976a5004ae9e2adefb9084c7683962e31d545eecc30c6a24f41d1faa46c37eaee29429d054a3a3fab3ed867d969ace402835cd77883a9ab584f94852d2b75066a3e07c98c56da27c80e79bcd6ff9e853754ec1e00923603ced44b9da8938a96e27ed41380d5b610605c95ac9a2eb8ba67968a5f3126cd6682759e932875d1ff5a7f9645b437b442d9075ff294c83d9919d91274fc71eabe295e30d0cf2262e818b172250bc88e3decdff3a98b87392e95a057e9a409b70a04343b5f4fcb23975f3f4aba4e43d12ded697f45b030e743e6af65ca1031719429299017eef5e0d10f96a801c45b3db87b1c5393017e8d23db7ce09f2d76308c128277c497e2f068fcb84336c5ae1accb4ee384a6aad0e89b818de1e39421eb39059c8cef7121bb7867f954c790d20d217942c2e26e44a753271403870693a06b1cb97e4727e7789f8768d2579744afcba13783ef4541f74962f6960e438f618695313f778bb57a97202e7ba8c364b5ce02ea08a0d0ae798c47ea875ed7ba04128a0d5a3315a8ec6520560c58fa07f5690f24dffd15f4a7d61943c20c4a7d288b671e321355fa8e6bc112a1868ce8fc11a588e4663ee993f9bffaaf9b4bcf19078797c1a5b2b0e06c4826b9908cba02919f9697b73f9f5dc076940b450afba097bc6f057d494b31124a7601b0da72009f7532c05ee599db8e8b27177c71dc731643bbd62fc4d0e6e660a46169893659c122ac05ba24aa8ca4f5f3cd9f9de27035d798b21e4b86d729b86ce11ccd25d657c4a40f49cfbf55afe682da9e584294966c45a053f9459ba08e28a4809fb46c6a932fbd2745aa50f8c5a1b6ea7caf02e8d832c4f4804654cb50ffe3f3161d7b3d5eec53c2a0727e516dc5bb9c400b64c574dc774d8c4a8daa861b727164fdc1e253e93e9e9f1af0c4877034b1d1f5f3192b9522d3bd60c469c7887ecdb13d2dfcb870ab0c7b2c9bdabc623f158117fe143de70330900722dc160825860eaac542c3567787e263583c39f01019cc59f1324a2eaeb1d6be4f91e93561f8802aa92c28f66e81a842dec1cdeae2b7b8de71826f1916aa7891d30a3610503f94e252369f30cb0c79ae41c43b7a6ec438dbbb3d6e167d38c2ec2a0d2a983ee0dce885d84d08fcfd88a010c3191bc9132cd9e19aeb1dfabb74d610af2e6a2f0a507987051709136b5955524359f4a69937305ba3f5105edda2a021e4eeed980b7c08c254193c01b0a46adf1544f883979849c0be74565a42f90d0d339cd8f958d82e795781ab542c2ce34fa51ab3c886bf71b74676d7a800dadb3ec785fc86283819234801a237de1c65d7ade0f09dcaeba9968152ff3e82010e0ff3d47bd49dfe2edff0966799b49120e0b286d0f04aab42e86bf8caf3b1b2133761e8d0a4f223e9893b460ee0008c14675f75e07ddf2501c0d9c72b897c5512d8898763352c17bf76fa2a359e13bf4449a0dd9ecd3fe73ea865b1dc943be34bc9ac96d7ee30a797bf68e58d688b28c3d423b354e4de3c0e1fd69721a6f053ea983734a9af8c3eb328730ea19a7adde7b9c7febbdc9a6f75def4447dab2323d9979b41d538c81133fffe690af96a177b699e55f7b4d4400bd374fe6821b0128ed8f28a4575cc87dc5ff0c2f4dd28fe7731d7002abb4d82fdb283c6fbc85f754d2dc1c0caaf9b1838c88ba1a1f83ebcc4a9ef989445c6525c35ea35be0f23b36c427f0d9a031eee89034debc432a5dc42c0a8e55c53b9ac4b115943b52e17dcabceea5970f982b9b074202e3aa63bbef7ad66bac0196d769b4dd621e02c755dbc5d77152422715c5a14994c6a43d0950877d276ab250ef73b0334ea86f183b225c00ccf48725415dd5b330acb9aadf059b4122dc57018c5f04c16b442722777890c01f393a15aef26e12d295b0abd288e1b1bdef5ac41041d6a6a39d740637a3ca173169cc221f2359bbbcc45c75e1fb81a40621ad5f9109e0ab3011fe4020d592b0b9f869fe1d7cdd12401a020a24a48c92a980ea85d2ab4c6a4991355d6de1621060dde5cf9247ac8ea2872c4e88a73631233ee32f69b7920b2a991adb648150663d1248580857faf929c2a37ca3a9d381656770b24ad0ba38b82db773347302773bc19be84712a72fc311d1f121659014f05a6069c84c05a1b9a09f61be35b0011883d74d8842e2229d867bc0ad7b76bbeea39eec28cd1e1909c9f0beee1885c78cecee254657601772554b5aa9570c3c89a8cac9c478d30177d2ca3c7c0bf0a834e1c7a5bbaeba0c5de885542f6a53a8a1850495b2cf05e194ce015b1e315dc4c395075d034b7e9f73a920b1eae6cb6fde939584d1ec093c3c54abe12edffa71da1e9b2de661e8404d45441c6b44e688cabeca78b8e21c8fe2c60c3f94fdc5719cf9dc846299b74ea7e82e52230b0956becc2153d736f7eddabdc554d6fbf0ce5054f9dac5a9e04a516ecb46008e5645e955498f4d3ec74648a0236496b778c769519ac33b9de6bc1556242b1f5fa3ba5902316fc2b7b7877411e2402dd676b998c119645e512c18b39bd46327b8977a238ebf4a53f3aa6af6a47facf1517f3687cf67db678b8d3cbc85164a3706ebd89908d350f1eb7e04ca47b3e89737793bcb6e914ae2d885cb835e0bdfa7660806fd3b5af3b10c7a3a0c4a368bee9a09358c099527c2795bc1ec9b92b1d559252879484973f2ab2b8a6a271b5de5a27b43eb626c1bbd2134a10f2f0b26743c24590adf1c7d82fb8a1149f106fff09fdcacc58f984f6ecc6de5292ea703d1b036139264386a0168da762a470ad30c4682a00f273b6bc4e18e5edf7793faccde75c65566bcd594d4c3b9ff13bf71b02e2a5b82f458a7335e8c3d882b03d9bc01761b45ab6e727a11efdf2b5cfdc7c14fe6787341f2673e9dcf5436b9a2d83154821340f085b3fe454371eddc5816ac76385c7a836b02de15882728783b65696c2aa0e05bdc8d97c0f5e526ab99efa8556dca437d51952a45c0ceed1af22ef19d6a7050d7780e6f65ba03e29299e64ca591ccb2fbf4cd5fb14b4a7f47aca51399a624ab05784ec6882f192f7bf06b2c17ec13b962517d7786791eaa59fcf541a00cdc4d731449c2aca1279c6c22d36a09b1f24d41c0068a161fe5916de57e37a1bf4fce12a7dc27ea529e762a05a6456c391080ed947e0b7ce383d364d8b8c9de3d3d73e967e94baa946d8a808035724c624ac0c7fa3f780b799c733eaaaa5278a7631d1c73a124fe1a623bb0d3c8a1bc9ec0e52ba034ce1cec099f11885a7325f711276d9948ca8870733c6362aced2f3fba85d425fc3b885042062a04f7143a188de71028bdd24f413c6f5f70263660f3f442cca74abae030cf3043c58e3d4e3c11e2eda9f5be066ec9afab3ec0de21d78f0f0fd04fe5c4c0b295cbd5c96faf4abac58d1b81f1ab6ca1c272732873b54eb0268c2794892442ac26b6951b215b574913e23612c15a8ea75276b2f6fc65806f3986f8a4a29f052641b0cc4e807756cecae19138761ea18b8d94d1215fa90e5a2e50edae4e31864a4b625f3099419343e487d31c6b1754aaae07d0fdf36d90d8cef99b13f467ea9cc317dd6c0f6e32a8d85d3b324a680ba164ba0d52c2161134c85feb3c4629e6db002de4cdaabef14f7d57ba20290429a3c88d9ca712da11d5301bfec11030940b7e6795ad330a8cedb18590199ca1e7c6d8a8f23eba435d234d78117a668bff70a9c064563fe647c92d8a3a9403e07074bbaece54bd3acb5e671c4a62ec073685001d6e266a97f4d72da177e4c4bb1cab2fb4ef87d1bf4d893a789dd2063aea0fd02e814817f033893a021487c5d14eb98759e1b1104f5f311b95b7e7b0ffdaeb0f83d64447a64c211ec08e58b69ea2dcc738670421e06fdafa6ad59f269bd8a82b328216662dbce8b1edd3637feab403948e702744370902adc973878ab9730e32da4067c44f9cee253d1fa3a6bf9376bfb875204d0f8cdedca989776553c4bbd5d524722a7e782264326880705d5481396bbd5103067e2e1ebad6b5eccb32159850d60965cafe05a3b58757f836851251ee915206828c49126045da1b683840dd7c2fde3ea263c02a168955e6e8d66336f480ffef1734df800df5ab3d46f895f8002dce1f7af4cf77c844b84a702fe282d1466b30da1192380853797ae726c6a568138ca5a6c7493794870ac0d9e2fdee5f176f2a57969590;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'haebf4f5764e059286b809bd41752a2db4e3fea5e91faa0770443e840fbe8b43f4b3cf44b37cf3d2b31755fd2aa50ca256e5fa37b212f30fc53e431a73cb578e87d4ac760002b04cb98b4ce3e3c3cfc4f1312c873f86c8ea39eb7e38465719f0680f026dd08b253742cd9ef611d9b4cdb29d6cdd4805c28d808106a6c71256c287db56a4b4e64b0f2facad4058f495d19e7f7ae9ab9bedadab6670a7bc8306c646450dd08187cf42f847c4362d778626f8d95018ee5d1d414c66f0424d61445756925247866d1592300d0e76d4d608df3d9b910cf643aa3e092f9696516f97aa894f16cb54cdac3b25314d55fd7e8ceacaea13b11589c75656482c9fd87732eeeb9084ede57ae7aa972e69725f802ceb7c6a0c9d811cd5509cf0ac684dd1e4294c74238f31b1ff10c82d5b9c61dc5a2eed670cc966e3a8395fde37d496573e544320846b56de786f90f90243cf8ad36cd5269c9aa8bbe73393d6a4ffe57a4cb2270342543bd6c34e1f44052b7c46d873482eef0df9d3d97887cebbefa021ae4c594b67710336cbba80a34c3c435d66f846b92c7794103c2f87d5b1bc99571e4e031fc49acaded70458386b796dcb4b3e62673bb9acc2a1411cb84970d3c1236b3833320641db405e0fc43fac202bef7733566cecd3fe0dfe8c1c4610ba9e7b26700327bbc5614aec7d05d615a4255fecc7e8062429ff3b90c19f91efb48abde69598c9432b1813d657fcfaa938cf46e696882b8330f79c1b68ccb1e151d8949e99a571bd6ac98c9e9ab6dc8e5064529f46546c4d4fc36d7e13023173edd6cfaab319f4abbdb5006a684208fcfd94d4bb0c787081ad228b58655ec021517e566c001c27402ee19896716cf6bb0ff0dab5a8736c0eb0cad620b879b177554d74decff43cc66466292272ea015b86b89858d989527c88d54932e56162268d811abd3f7dbb2362043c56a776e456d35e2c1135d3e447f26adab3470f2eb7c649ea37abc6a2b284afa305a6e9cc8e2898cb3f5ef0b68599f0f53002a69edf7de8a9c395c01fb631e19af2cface2128528cd6841f65149aa36ede111559b2199e6098816b2542eaa0f8e89009aa6051a447b9e2efb9553b7b4c75eb6f69feeccd25d3d5d22c4939be1dd2418cb34818f6d1dedd0a1555b8de736a4a1f7d421e44ec075f9211d83340bf7538bb133cd1851f941cc753e3f96c3c16a00e9a174777ceb8703471a27930d3a062accbac35e990edf669b9d860b8379c64d1b822aa90ffc580209f39929f54f69710124fbe58d3f3ee0dbe9190d4a9f1ab3592360b03834842ff57c90871269dfe9aa33c12070a296f582e0df9165c1862b5c9c20f83b11ca707b1fdf331616e4b6fc44c5700e1414db07aaec27c26baf5d931cf648423d2ee9393c04cc1656de5ed1ff22d07cbb1748ecff8d400f8afc673bf308aaf8527cba078ae134f263f0d48bfed287ef12b6c6c646ce62753e492012c2351f733f26b04e1a9107d4818dfb655bf82d6981587506700498b0e4431e702e2688df75f598d337e3381034e5633753e6b045da153691c324e10b18d2753cec317ad1d7d30cdeb3374816231baf5a132d1d8c6d4098b3c8c1e7897d052eedc231b3894987a84bc83846d7988974f03ff0441191395a06db8c296acb0848295c27d18868e566a195530b5d74314f931169e105ffe4fce45f5fa67f4e8d97be216e9ba2cb5171710ddf0eae7f7615c2571a173ef613ed109403425c663b0c06e6804b765a443140f5e6ed29d417c8a610539707864b5c72ea0174836098949b4bb8be87f124561fd394806e7b0e349a88a4fb2ba90ed43998bb4ceae8bc309ef3a2021af8b3f712dc4d4906ca991a7f2f87f9d7dcb565df7cd9efa0133d7ced71a3bee7fc2512f799c9c0f9f1b25a7f402711d41bbf19f0cb287c36e44fa058be34cbde673f0b788c73b5546c7eb8686779836e301edb60dec481ed4d56f18338ed79dad050e9031abd22ae52551325bf8acf1b6043e4733462b184b852a5d43b44ee8d9fc864e0ad43530bf1a59608e3a841d46eac3fb3157426de36b1a37b5708a849c294bb39487d63e3114e04405fa1f15543590e2e9ca4407e0e1be31ac3e1d9eca8aafcbe8fb1d493967fb3d7ad89c011a536dddbb9a134cacf4e1208d9a1f019b6c10ad1a1eed87330c4e9908c971302fc83551787e19ff4a669a813bdb8b4113c9770a38a6de8059d9dee9113d2f9ba71df072e1e6e535bbbc061ae839ab125f8fd4c61774a1f2637d50aa70d64848e9c2d85655427bef71dac72be51b159746518569cb5d6445eab9a22cfae51eee8b102984b339932415d5468d6f85f9e0b2821ece5f8a1b38a0acf0a0a53c1ed54acdd42751f98a87a1bd58a5eafbf5d076092dc4e0a4c53c4119703998c0eb987d17b78a5e00ad1e3bc188d26f216182a08ee1b3856d231a43f24ebdb265b1f2e1fe9687a6fbafbd2404bfa1b15a3b6d8156f52ca0dec20265afd2a4f5d61619a702d605055a6eafd5d013c738c083087ad73764e9b15d669a1d8a0df89707fb09f1bcc7b4080df429cae466ee934095ae211aab9dd6b583f19938eafe0cb89d02706fd7c2b98c2b520c7f2380ab880b7c09be2cc5182e8a16205f023e4eaf40f45ddcab0ab32abb0346d711c542ba983a2903cfe1a2a49b6fdc33310c4dddf58177f235b1bda1525eae7a033748f987c59c7f90dbb6f03e21304448343adf9d60d357b391781f5572778a0361f05fc94f13f74317881afc860db2350edb579dad36fedd99edd8dc0824727bda9d8f0a5313e8dc3344e7d29d0226285da1ce2a772732a9ad38708ac4da15b001dce37e804d08b0856fd75daade93ab79a421dc0f5e56585916408803ec6be56977c7a68d374757d83d8347bf37051a997e77cd0d1fc521e30c59d3f2ce09a226b5c3810aed5007bb762a7b72c99e86019299a15e38f2cb7e6c6a244c8fa69ab50f623d19d3928f713ba2f99da4f66335a1f56322ae01e95d94d28290d2ff9b9dea8d3275379e0b38c99667259fafbad9f448a2ae0e56b2e894052abc9204b565971fe68300a9e63035444cc171ab8d81f82d6833c37272df1a1f9e6c8a920182b8e999b4af4312f47dd479d5735c74ea5890c2acc8038b1b26afe144440ca57fafb6836275b2bc589324b2dfc61bf8e45abd64e568f97cb43f5f36b5d7accb7cd9e7796a1ab54d9db56c8d40c9de024bffe2b94b0c2e0a268509c5029e3253a412da8d87fac56d93159413e73bfc28fd59583beed696ef6bc8c1ee8565a8715dfb4ee7a4deed790307e07d2b1f1d6bccd573da907727c7054aa72830d76b6a68f9226bda5af5aed0ac3378c5ae2b3ca36bc728ff781024e51d0231edcd0d7fde11139b7d22ef2d085ea8f13cb7e5ac238b021b6db2d7bf10c7f15c0aee8a498ee4a83c695f3af3a131beeee0c6d0cd978cc0074a1f8f5518fb592f615353ad3cea4d977f32f78826c24c6e65991a18566d3f2f3d2fa40121fa27467cbedf3c3fba574b2c511dc733ff12f5c6879a79954624c47cc3ea20cd5e0962cfc96e1209df7cfab50b7ed95b291160ef9ddc787ac9077e4b35dc8982602328752e94e6509a5207d5f07b833bb575464982deeb0646907b86b1c24a4dc921a192695d107fc9edd681baef4665be66dc7be8d232c77893aa69b68cabb896f860835aea562369c561ca699e1cf25d8692a65aca2d0ee160d1d845f6c991f1ccd007fc4d3e416cef073970b4b1a4e3bab5994cea2c9ae90737f99873287bf1a19644bb426277bd02a69287dc7f43377e2ca4850c7c9246ba14dd5509a6c3bcf1fa195ce7d7f99cb3113801be759f53de707909d7170738354a3dfdc21a3a8fce9001d13bf1646a27ba9c23b8f39abb42d5f5588921a0c7b66309185eaf47bddb859ed7bbbbca15f0729501d27a33be5ea4e02a172e82b9af3f8a58ce197d4e128ed15566821ac674dda8aa0f9a5864e89c834701ea0ae270170206941bec288d81e3d2958902d9870cff82675b6003072f4a40942e6a7d084b4dd8af2b76baaf0156bb6188b5db736763bfa58ae9b86aff946ca7846c3e4f2df2ffee2329dc979918c67f177ffdb2bd3da6fb4a1e2baf600f0c43e384c0f970144314350bb4f03c1d5f5be842a5e7c20dc19115e96369c2f920d97a3cc7ea6d3edfe7ac3c179d69e2be6a3855315b5ca1faf1d769aadb1fc51b5e7bfa51fade7be8020c6d68d51a67e2d1a11ca134cdb026faa48525f65370206c23e2fd7f88f7ab68827c70a0385889b47326ec109d44b461c874868c31017079f841f5865bcab7b23e9ad399358d3445fa5ffa5838991807186f0b03a1e3d76956569b3ee63a91513ca996ef9504bbf743c502076bffeedf3b1ca9ff330b5650b5c401ba041f4ba75da4b57fd737f1fc6762ff9e68079e02e009137389dcf4c7161e6652c2035bbd5b12959267fc47271eeae9d16c512b27d6459b4d479518d8e79cc6004a5151f360388f6bd6bcb32d91a3c36910b41e1f0f24e3dd3713506bc49d4bd3fcc758bc79cf4bca7865d360e78dea868dfa27bd471283fd5eab489b1cc5aca91c4fa470f434e10063c343cd5d52089a792f7e80d4d5c7c682bdd6382416f57ce0e99d6265bda5643fc4d84e0279ae2e321fed2195cf628b82d02b42f6cbc31580fcc1c4e94f71687d7485f14283f340d7af324bfb979147becc3ff44fb2f6e7a11acca4714e0eca6976a49b5bcd68b0ba34c02abff25b1dbc88b7e0f6fa2b81b1e7c22428e234a59418e857648f533d04d7b72274b36ee9f50315e8bdce5031419cd4e94d6d526f4e593dc06be9a5222a7ed8e9c6f502b934c1c7806f722e45bd361d6b3978f90bf759c598d7175981fa12c46b222984fd926a6a79efb5ed827415572638fac77ecaecf5badf8448026b0f7cb72baa429a66879e3d588b55c7324bcbd2bc2c6ff68f574e158cedf1d8e312de41a9d0610a020f6aa098b77d029a7b32badc20c5bb437f59de3cb80fc902c229581d650ebe9a79c7d158b9081f988767eb73a2afda823030cdf96a8bb39ae8171a81a451f277319be8d72ab705bf98fb256812956cce0096baf4c50421488178856991ea1f38575f3072fb64f42a34b8f458f9d83aeea0052424963d2adcab8270cb7df58e6ad1e44477105a647ae38d3d0636cc488db4d2592f8774af4eff5d0b2662b830faaae2f68417952bfd7631a2713594f9dbbf93ef7bb598376e6bdc73e788265821ad528dcbfc19b2843c4ee5d9e60f58bbe8081b2fdfae2c3076673d63bfe2a673260bce8f00ac09ea5c59af60447e8949277db31e1f722849312b5f33b0f29a9b07078a8f6ae04e23065439f2253f8b5995ad134cc164ccadb0d883b6da3ee24c5792a93674385d361478847f539c9fd3b4f33b937d544bfa4f71169b918497b17fc645bb15fbe4f353348207f98f2bf421efdadab7085f32a0df70ad3dd828d4106f00e87b2fc1a03d90c25e32e64a6a74ccb37382fc65e3cfc7869a2c8f7ef8b8badabfdddb635d7a768b36dda087829acca68d9d6214297136b54be7bb4b6b192546cfa1662eac6a710017838bab50797765d86f8f8fa96ce3f1f63ef021c7bc0d3f03f0ddbe26f44d32251ea90c770db67b2b54837a19f0962bb15797d46fda0de37d0db4839f5d046d17d02b5e17be8bc68ddbd7513165ca27a76cd473971c91a4b1997d0dd4f424e39475de86e7de89faedd0a555aec590c729322e833cc297f40102bed14365684e10c12ace33e09e1f6e30dc1abd8472d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h76475877bcb72d551858b0e2d02403e2b2dea90ed347aefb798b0505bce17e3f5870b1f40545cc8a9ea0c0eab1801f106c03270bf5dc1acd7c1faf38b250fd4e6f68b7447c258e2535d3475e643734f507fd3b28f87c9851a341dda38a6368416a6b5371397c32c0b8853cc9f7ea4407c62d11bbb5ff989e75164ac823dab7c1b38717e75577817eff26171b9a94839d30a18986e2709ae997d2778e0afbeda0bf76bbd2060479f07fccd07c2385c07d06b94331202dc970b0ca4ffcc53e83d7ce5ab12c0de001855a26e188b99517140a9a71c72dcf3d2ad92a92db8df9e393705edb779d9dabc5b376a0a322bb63e7c2da7ee9336e8fc0014145f6c60017983781d7227dbfacaeb23706ccec6960d78ffe57aec29c779fd8255a351e62b6e32e85797a300b12aafce74cdcd0ece244c146e4db3ca5ac4920fc985fa335bcf31289bd58c0cff78d53af6cf43fff09dd1c153b11c9d595e96d9634ccaa59bd76a0908e81795000ba89fcc37671dca18607af40fede44dcc3b9ad132937fab72dab494a847564d3be5959df0090881121297cb4f8027a99323a9a3434ba0064f04d2e366e5c3ca0fc3cb9f999ebe163f4197cb75287c913ac7fe1deb781f8ffdb5c82a46b7c8a327359995da860e811b2e50b7448a1d52fd91f3f7cf10a5043cc398031f7eae850b44e9e2fa14e84efce0daba0692c365bc64a97e04a40ac3b02d437602d92967e5881b7a01d4ae96c473d27262f92af30708775e98ddab3ed2d1d5565c7c3e5fb4e0b609b8e9e93991e125dc90b932d8edb44a89c771206c78bff3ec23cfdb309963724a59be59c8aabcaf0bd6fac33aff7b03116c29e004d013177b1d93caa1dda8a2b19f39df3d0db67e5169953515b99b8c5573efeeb8277146d462926a744e644431f953ce33399022b4f3eac9ebe4f66d59854f919dfe58e64c833d73c2e95ab83805f548c6dc69b83d3c5b07876111a4d90db1a20aad8e98193e275be0736cf54a116ed804ce645d7b605df3666a5b2d948cd66ff87333b835cf189bee0913bcb256a910d4c9889a6c1171fdc5461494727244147789639c5ce76310aeeb024ba43f4e9a9dda9665f9a09b0ec713d089c8361627a4a6ccfd8a041c62645882a3042cbbaa2bccb8d3c8e3094f1a5ca739905d7385467339c9e7f645727a81628f74d85561e6b83d096ffcf0c3e8d51aa834fcf55aba8b3f266484ac26492d0cf2da14f506588a6409ab8adea7ac4057d9fa7df65c7ad373b900e6b29bca7c056f8ac81f5913158a21cc41f33e2cfb449d7bbe3df54f624ee6b5f03755accddb3c1bed237ac6da6dc4475ccbd526ab1e6ed7ee754ab3e3d3e6790c232072445287c67f74b1edcdb9be8adebad51984afd42d3feaa591487214588f6fa99b6eea5efd5f9ad3f46c0f0e37dd31e5437bb3cd92be4ab99a195e568b11762218e21d7f53aea7577c7215c48ced968173e16a9cb79269de82795ebda9c8a31df9c86016fc489d8fb57a134d1ecedd3c1507e13c563c31620798866a98a98303fdb5e54989f8498a5539f3140319bcb20a1d0707263ce6f2295eae85d93782323018621f25e585527f498e37108396ed6c4b251fe78f626dba67dae6480145d84a00a56acdcdd4cebee569e9f62b60cfaa7e199f7569492e2aa66f3ee714e3ede860fa4ed8d7eaa15a7b5d153c2ab33fa2726612417d7838595d26eaf20543ed2b145eac68de3f8efc4f3b8aab400cd513b1c5aade03e654e4a354457b1320b17265cdd3d06c4679474298b888a69c9b252ee85d9db1b5f04a6aae98e2e03654e93296dd575665ed966476eb46a9eb12a5c8766b301ecfc9e52212116d33f821cc24b24e64ada36a174b7a81ef238c13cabce205bf9ff060113c7ef266dffebe02a07ac022fbd2ba419242debe7570a23a20fa8b35bcb7a5efd18c6fd7ec080e2995206cc21b0f0aa9c02e8ce0937a22914f21cf3a134aece0a832dbd4ca46f11661957ce81e33eec94d589ed7cd08737adef0fbfb47e07051ce7b868b45ce5000ccffe529597a59a4dd7fcba03c77c0523d1b5245efb9674ba3924dbc048a35be03871d8d5cf77013fc08843d2a495eba69e78ca98be83bde674328e4ca101180dba3311c9e646a853d241ac348740201719e349ccb0aabc647d7c1bcd9212b2b73ca63809f4c45c4bd48b06f94c790ea16b2a55e36532319e0d7186b1055684344c56033058a78082030a6ba6e55496aa5edb290afa05ae3bf94238836e63d671195f6452a6b8d59bacea2ffa488ca26ef1b11937680c40c21f22879eb0522850ebb1bfe113728b99b9d7ca4f390152476cadb9baab2e069fff9f891d9a62b1d65dfffe7d03bc5e0a00541f0e944f8bd3b995191c991021029875b797f6e1e28a569ff84bcf445d4e691c211b858d3c0eda78f5db75da3dc462fd256ea58e89f78969f1046ae2e1ed4610d5070f419e47815d0611a236f98f7961e4f62579a6f2149a2c8560055088625cb4fd4b8371de61d2b98f3ac62552ed49654a9a0e65bd560ecad347385d1a47e6ad2136066a9e1355d7b28489f7ea191486c737931d1d61feca14bf52208a0566ff2de7b4195b9e9bfd255ed012236ddcacd7087807c902a7eda2f44e8eb1b790a845fafd282a6c0317bc4fed74c86add0ee6127ca85bbcd814c33f5d6af1b494aa976dd1e65d1703ab6cd32c5bd2276ee53a05e681f7da02492e298d9dff386a49b4773d875c4bc5eef867bbb7b1f72582f95ce84b3f890f79cd41665cc403fb56239bfb6500b538a7a177f7e00e4fa9f00cdeea17991308fd5a87b2d40b6b4816364e3dace0031ebd1104a24708cf99ed1b3aed53165aee1e8b877cff328219294567313ac78138617f53fd56860efebcfe88b6140862d6faff99027d19aea1cdd9f6c4a8310bb01e52319137ca43be30399ed94ed15da943347e6d6d6752177d6b37a2236401fe2433ddfefe80450550c7c52ba0d8330d2403d6d3490acfa598d1d9ec0f9f870e6809846693c4da50d8c9ce920499030c0680ce138c21310bede74aa5eaf4ce472bb8b61bb702891ac7c973bacc11f05891096777beb0d819bcf16e90f0b635a3734e6b397e2ac17237c98403bbbf806a7404c10ec2a97ceae87a51c29f11aebfaa3f31c240d0b161d88c14f5269eefc6abed68873be87d796aea9af4f45400574d27ed6c40a7c6617ff60600d7b689260457f251a8d7888c5a37204df1b775451bb3f911bec2a3753db74b0f131cd973b29d0879bb02ef1feb6ec445ba4b154a88e57dca8713aecdce3417e13fa64536e7b4c1003d703e12ca959f15638b0089feac8ee646d64c3262a662fab666930d508955ad875cb139fa75eab61275ed07526f920c847febdbb51209ba50f5b41253d678238c3a7292d1488fa741bceec3bb3ad6018b9c0f2f4b1761df7e3221746e587f24e266ccd512d60c649a59ddda1097a075f862f7b2e3a1c4e9508abfddb6b3b9516a2d971f73b432c2e1d14e8d585faee61513a3d88468f2850c72b2467fd465595cd64643ffde187408034876265951fbcaf3abbef250224e07754e1305a78ac318067f20d71876a1bf62182fd82281879e666236f1e3d5a792881e9ce9f796bea987b41bda22a544ad334ea2e39f8f022b4bd020ade1d027d08ef9600b6ace12db9130f2a18c62ab3f8887fd981cb40e28d8ec5bd106b6a11113d55170f31611a0acf9598c97716a72f79977a3e163b26f573a1640fdd3130cb053a7bbdc339d2f22667b3310cc15a614c5bac507d69887c039666655f5c61303a517ffc82bbc20759d1cd468cbf04e5fbee3df5c6541e10f09a498f13ae12b04aba93986dd2184385a7736de608480eea920c4dffe17aee0b7bc9271971f81805dcb0c448ba370b5d1ce782f848cd3683c69140a39b4dbb9618ff443404de61a827751cf978e7ad9ec31db26c936f8419cb03d61c4d129e33d0bde29dfc2e9608659b0a790d49099c0988e1255480234602363af0ee42225489da2c9b18de448fdaf123cfc2b9ef3897254b3e22abf5c5ee30b5142fa055ddcc322fc734cfe181a2837f01931158a07836d14e5eab4b3029e1e27204fb3f20a0c6c1402f17cd433bbd51ebe9832498b56e6b569f1032f20cf5efe758988827d8328b9a04b2e6e4a4c08085d97f81a666965bbec3a4cb9a9dc862e16a5284ea61de5dcffdd204db4f46c6a540a19b5e09852089542fc5f495a9ab2c7535aa1d83eb05500a00662248006b9cacc8778b25417113fd641952e9307265797488a94c062e7360a4aa80c5680e4a313f9fb1ce025f7474d60abbfc69974d3aab9e6c94a4cb71c871ba738262f40999b86fc7190e3d4ca726440fd76c56176b47049f74e2467b109c971b1774338c8d8176472e04d5aa1d6d6d819afc6400d95d22717ab15c5c047c03838f90e26f2bcf124d706fb1a3443cf586abf583f3395a30fe96b4bc598a12ec3c3389ed60c3edda358eb0fc21d0ce43fe369776382d995f6c1e37d176a9e10e0a35ead05e8d56361b53aeb79c9c1dc6a43dc7703eeab1b8e534cbeb1561af11c6e40f09b927dd392e6482348468f8d546a936ba83e8843f83093db3734791469d56739bdf649b712f0332fba70ec8035f06cb2252b1c74b41dd5626cc10b2e1beeda3433dbf8e3708eec50e033572b957f9cc99ac0578054083b01120aca2b2b25a9c2b83fa552120e5896d4a00cae609d07ef6c0df699a7edfa7e054078107f76c812d7d32f06948dc3e0475b0e22fce7daecccddbbe73f54acf210ca6af586c2c0212e1316feb447493129eb2f951b8503112dbdef10bc7e2bad92cc6c3c0b68138e2bbac4e82ad30c2ce915c6aca987ca4609333f78be40c40eb32bfb3166c260970c1af4ad8cf5a410261b075e0ab4ac5516c29d514154a8d8d5a9b34bef8b323abd63ce98bb80bb97fcd258dd6be6bbd9ade7c74be864240b5289aa8b484a52d53166629da7974f06738c127d819322808753c1302f1d113e4722897b6da3c03dec8d3e9aa2e8f5d9f2bcbbe107317a358c6f7564ff92486deeae35e56f7fe47b05b6356d44e34c73962feba9244199e91b2d4a13c9a19bd651339c4b77c42dc3b044f6f6f75314777a4e629ae0fb89cd6239035fddaf9ac8416ecfcb725cf70202677258b23af529115191120b990653d074ec7ae066d033aa2dcdb12a75a3634a91b62d5d13095a7256e53a21566c8cbb681e3d8dd9bd698a54dd77a163317d3ff39f26f9e0e8e042caff903a4be0fad37f86235be3014ec9911bb20681267b30fe00c5326e8f9f3d67da96f56b24a41e6ae3d3995a0cf9615ac096b102e8a535b615abe4a2e90fb1cbe39c3fa8bc1df021208a594e361beac8ae2b674dd5d145ef65d273c9c80e4ec5fe83332d8dc1bffbc9586fcece0823ef797f264c5bd74581b32f95af3745297e9d437267cccdb04aad332b76bdee4e513a210c1d4b17677902d923a7906170e0d121d762f67ecf24b302d054f88517f4efc42fb5c07cd8fc52f04bf49156134bf2491736405861383a5929782e4483c69c6fd7bed25ec3042bb99c86a8224fce5358cbce826b49c3c983e5bd879a5e01d762a5eae607801ea1d54a89b2c96233d39b44ad560aceedb301b9740570815312fcbc870d66d35893bf546c8084b5652fe413d2d0b691c08630585fdf0c4e7327a4c9ebaf5bff997b7e35c42a4d5da9d4637fbc029afd0cf5113d97cd2d944daa38ebc1869c7782b0d28a95724977433dae9168b06cd9598a48f470;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h90c839103eb8ccc75d028de01f282c740228c1f6e98293cd89ac8443b794974dfbcc1b814d72023571213647c0d90684d12849f710781721a140d3755bf2829dca7a86eda648365909e9c674d9d7d5d748f6108403f6ae6d9522f5d1e38bc007637e51bab474dbaecbaa31e0e0354ff8bc12665ea115d9f84d4f87761f376ff32a2c31cc49cf923d94fcc942a55c6a7065460fa8fc0bed318a17d8f3988e23ea8ffe2358e08ee3039e21f2bb97edb1a729a184b698daa51441e2a1c43144ed0b3c3d6c4398a3da507233aacd1507ddfe3186ce89fbc2a7f024bb98bff9972d47f2d612a5781c57a95db8e7cc651cdddb71f437cdf94f30e9e01d2e44b3757203f9f34509e4eca1d0efc4627a01b9b15dcfe4e394ba1b7e6aff9434ffe82fd02580fb1a2d15679031ef0b755eb07afdbbf81d80a95e6f9de22cfc7ccd22af7f21591e62b9c9de9c0ca00e5e2b1cc71ef162fba9ec647fd3acf4b6fb058e07357d7e2fce78617f6851f1f7124240718967e63bb31366e6606f1bc49418f7e4ed46cc5126e01f9448c90648b96bea9988f815e5b9cdf9f0fd562ad19c6c9c1c1083a3acfa09ad8dc6d9eb4695170489130d4561978d0df16ba94e3f22ad1c4e74c62afe3b222781d50915b6b681aafd6d47a496094998a97c0136ac84314ea49c8326b4565bb06f6fccb7ce7a95e04e9cb14de9d1808a4892923b18677651902b1fc296ad03e93f04aceefa6d3001627dd496b3948c5433d95c9c218729c977c7f659a6b960b1773160e479f9fce1ff00f7106615209a47e5c23913626b7bbf693d4e7cfcaee54d1c38fa3a277c7152ccb48442cb7c81af670b63cec03fc2558e56e5ae775a1af0130bc7c54dc69ebf51d1eb4ce2e976b7c5a0549fba2e2271012a737524e6f9bcacfe1338bca59ae33c7ea7cba7477e8202f97bc0b7999379739f99cc6af3879a232a41ccee22ef2db4f743ccd51de665d1ff12355aa8cc0d87ea0dcef150efa7c11dd29d90454fa3c5a1bd3492776f1681465836b54b50f8dd666126b3c91b4fa51b714c44d1c1b663d01163c3ad68ef07450522e87b7a36612555542e5adaab5f717abb521d11eb6ecaffc404d7413845966814e2edc4b9d0c8eb4b64a1a2be7046bf8d274adc083db0beaed704645ced1fdddfe814513a25cebc024ae787058cd88ba82db7cc0fffb53361653d3c0bdc81e1d5d3ed9b9c9e1c11d98c3a3c91302aad71c3b29c4e4ed65e689820cff33a7e8b8fe6e6379b66f7231f4179046ff2f067bfa17869a0c1c75601324d4d774e61e5bf839ed6e11e96ad776b5281dfb565df3f740a63d8b6590d942fbabdb37ac3539f80ac40008450d88af3696ff5513ef1d02332240809c05a7de77352208650e971aa9f1ed8d3fdf0d75ef8fc93396c1db8c2e3058957477e4981ca27baaac425dcd2d9dcf90cc804e4de38e8e87b731fa0aee689ab2c96c7d362c84cf95a2b3f1c5edef5044352b2ec2eddd6ee8b6d67e75a703ebfeefeff60848e817cff696ace0ed7a2f9ac91c1fe5b1136c48b055d148134e8874595bdd5d681a438b88663a9bbc8838cace4f4ca884ca81047de7a77970d72623af09f9000328796b026e7ef9564902d13ecd8500befa3caf95fb90c3d9b655a540726474c50c2adb9de12aef95f0d5135db11bd6e76674b703c49f5a68792b757dd5060a464219fb4e984aacc75e413196dde7274c94df6c96d5cbe7d23c5793375498e31e1f2ed43fe3d93e882d6e8dbcdd3b574c3d7954674d1ed318b6a89b176df3ebdd2ed0441746e94fb4d0f7b5460132138066c8552e28868cce9be29db8174b1b698246aaee8d61f4bb8b5cafda237374625d86cb4c86b0e8f4418fc82dafe386e62e88d88d1b85e0219aff82c2092d11213f4e0d3c98194bb609b70f5630f48b7cce70206c2c43de4a23079dc2a55c63a312925c4aa8a77848c4016c98158ddeb728dd7ef705ad784a5abe622175f6b1195c9654fcc6a380fbffc79fe4ffdccf65e05a60a96c9b7ab3fd07a0c6021acb96599f5752bd44e9b34cf1d8db6e99200d6a11a03692d54fbe49c0461e6aed6fb9fbf3a273dbb7533b18831a3ff5b3edf10de11daf44ae58ae0914f77ecdf48c7692d17f1b66a6d74663dc18bfb528c041e57b8474282f09bddaf2d50ffa2e71131cf482d7507d57f34822a00044da85dc601f7663969174c8879ef57e359e83750be353f59b38cb3676190bfd4a3657857fbd2494b61371e9beaab1ca0e875bd828dbae39838c9899530565a2d5c7202251e2ac6f7fd1feeb885609cf5e8c66c91f69e084cee627d74563f548d4e2c10f4c74632be1bb09a3ef6f480fe631061205e1c8be07ba64ccee203a4b3624bd6748268049503b5ffe987d2ed76038d6cc30bff4678241d327d2ebc004d388c23125342d6da9aaa0d8fd1c9b5ae5a025e81bc58b4972c633adc0626a368b8b3e2aa3130ac6b4dab7e4ef2a12fff92c100fa226521faf600b9dab2410a7cacc68015a8cd73df71e9c337ffa570f27fa3dcd7aae7de3406a089bcad82acc4f010ed993eb150e3a2c9be738e5c616518d303d09dada958b18ce902228a1f9efcf3001b25e3ffce6aca865f82a55207beff3e044c71e547674466987f66ac7d9a51b70eb0d9dd51ee1e1c613c872f83cc3a44bfc7533be0ee7d25af5a1633103db80c4edfe606fae67d906c2e9408271b494453b4d68514276515949d28dfa548d4435763e5ac3a0bbe8c8a2006edc302fdc149f092d015ab05e209cc7f347cbb19d94ce7533365bec1c4778c0c307a3cf17b3fe0f3a207850ff1fa8fc3a741baa3cf917545e3e0de3aca89d3cbbda684f9eee089b35916e93f62a61746e62586c8276b1127f22dedec252be2a62bb6e5a677e29bd5a0949b61a5fa47197db697f59d8e4d9b940ebaa72ad968c54f6781fe8ab68ae8f6896fb20c83b683e4542b898a4e1567a3aff1dc2ca1021d6dc8a0e37df77af22cdc59c4d70e10ffcecf4d64db05e9e9407000f272c35b770e63a524cbe2b0c26de1f336e0889a8dfd19a72ae24067e6807d9e71d2dc347baa9c30464daac3ccc39f013663f899c231c4888f189df97fec189a5c2e4189eb33df100b996c73ce359977b656fff2aadb07909f7733c742224f68ebf507eafe3a5be48dfc64a0e1e1084a04274bb0565a94fbb1d84681a2b1993e4d050a372836829d66440eb9a7da7226812cf2ab7d3f79ff4a89fcc53d6e323158b5430703608a63b6f0fdcda90a723371736a122fbbec98aaf4d8553e3071be150050897ac5bff2ea6c3401cd24b528eb20af7dea6035f6de2d5f835d41396a1d6a85cb43456f6e3a7552b5ddfb21012f9b3550f48f3815a33c5ab31ddf678d8ea19cbcf90d92ffb71c9914b4cc2725480485e29f198cc5f32d46e6161bd4111b3f72723a5b715ca9d251287b11531e61faad809327ba6478f9cf29309d6b97327b487784b2adeec449192f2ffe4c3dfe44b929d7e7213eff3efffdd71f6fc4898dfc78099a1812476dd9cd0447eb29a1e3f68f46c6e7432e021d007f3f782e0c734a98020b28f8eaf7d765f725af2831367f2e1ad2cea1b1f40541fef2a01987b32f4e514bf6badd51f9c5944e489ffc20bcf31b6322a9cb6b49e000a73049e96338540d089094849f76fab63dfecdced3d698ea6b62a63dafe47ce0bef32e3fb96ef1b46c1b096bd63fbd630d88a57954b067ba22bbcae820825a415cc3df96fbe4a8f11bd0b049fded5d3a82c5d15b0c26b0d72bc4b025b4107a931b26a3bd0eaa577cd42f8c03c30ba7ee2f695f579a7de9decc28116a26a6ed4a6b565034f07a8b93290765c7de1352ec37f8c1a300fc9534cee33ddea87469421c9f92f4bc30aa7666d519aaf52d023a3861aeb8f120ebaa763d655b7e2e76794b653517037fc54a4094af7a7177880bd4a794caa6470b2c1fd729d0d33fad33928882649995279dd6dfaede2a564aad8ae3db788b81bf455309e1fe57d7571824268fc80deafa090a5e0296049023acaaffef8fb8d607471816c621c02a586ae95d6fc74c7a6da8c0069b237779939e91f1993e3c1fc93a8a07d57a8548b9b08d7a2597cee2257626d297aa6c551ad20c5daa4af7d0b5fda46989b18f1ae739d5687f627d6be42fdfce7770bfb30673f2400751f4ffb404f6236c741a4a546d01fac5ffbb1ace034d64a4e4a58f28e1df7faff3978b6fa8fc50fafd9921b1d9c6ae5a2e081f4fafba97d1cd116e2e3c40ec5d6667f6a39d60da5b54b6e8defc4142457e2e47bc8d16c0b5870aed0d8cfe6bfc7c757ec1de454a30aed3d9edcd4959e4fa56c3460b6d9431d3651c1a616d9cfe55f4753af92e1881d2775055eb89174b7f882252d13bc0bda22ffd2ab72f09f2b25e81084a2d1d2a01c80b6166b2163609737ff9995d1f32a10dd2f5152a1b0622121f583652c511328f2b90476e6b6a7bca14f099dac7755b98c1b784b72edb2bcf1eb7ff0ab6b27fe9ff872e2cff7401520e382cbeafcef4c6b5b584fd5f28c9d4ccf59d4c5a42672b5e652e7e831161ab3080a6143e2a257866f898e0fc55d760abbf1c68abdb33066a28afd311ac9a7b384b876499918eb00a1cda6ecfd8f9ad5606ee2d61dea1dfca9b6db505b1e262531c6abdb9464c22a27b0da8040cb65382aedb49c2a4b2bbacafaf23bd5345374a79f8f1e05065afb5f05b18e26e2bcaaef4151972e5dafc762c189662697b218e09f29c2fbc124e4394bc26b92e908da7e4acfafbc4cafe5b304b8690a1300cd43f86ea474e7b46e07ed26b17b8d8deead4b72740f9a334cb09a5cafe24611e07637c05b91a1e80fe02a8fa5f8be1676f43a65d0b28dc921f1b0bb1f12e75442e506292c6392202e96d500584b84840db74bbf53376dd3e65cb7017a02b320629d67d80bd895e4006f3203cc7bc9f028b73569ef3d349dc05b14da35ed825216cdcf292619f41cf14c342424a09e71aca3366f8b7bddb5db0278238a3a4f91f889e45cf88f2a2f6910bd3cb1649be95438567da86320c887b7ef1d802b05d74289c66c0b43791a8ed9f75554e49b9248920ab2a79dd33baf3ca29da3a8fda03b810a5402e3ab538b80a236ef287d70a1744c4312272de8934b7ade185002d28008cebe83f0aa768069cdcdd44dc8d67f30496330bc56dad30b3c95f6f0ee6a079603655c4bc40dc062bdf457d8c1325da5eda7dc36a490991219c6e0a752aaef49c2c76523b8f01e9f40b7c1d50c1468b38792375736eae9552f288c1f63908f9c696f59e1bc1ed47d9037e299d53696f7c205f36e54da75c20b0afa5c297b0213bb8221a98a83951bb4ae7ba5353b46e2c15eea69d49a9f8ba81329875ebe8fe689f83ad2bc2896ddc812310a1b5444f1d77ce5e82e4fed31fa29487558861cbe3bbf930522cdf3de2cbbe4950298446ff87734d24ab039338b19cd2b420c656a3e3dc27bd229753281ef3cc642cc9a84c80c3acb5c197c8acd17524864697a0a05211d6499eccbaa145a05cc6fd6cb72be3fc739cef03ca6e669323430b3d865219498534ef5354a1fffe6c253005388a3a3194bf86d7863bb420a22d9fa95519da3b28ccd211b6fee92aa32cd5663e0fca45074b598e5fcec72104f356e884261859b5dd71b3ce7dae2eb266b83ec3fe2ad38f24a57506f46b55c38ceacd2bd7ce5bdfc117be283ff93eb3b71adb531879255f25d9abbd2fb86469a08b150ccac2b35fc303807a408df59e768b22ec427a4aa56b0b37be43adef81c0e65c8365caf5a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he33cf90ef6b492c5ae3cde45d234bf1578d29b2f9e810e93f98ae93060b66607e2d69d9a52ad3b8214d8385f21f6544abfd20feff96a98a05893bedc2aa7422be1812b25b922608840143dd66a97d140665e12fe6baf86247fe6c9c705d5d72c0ce61807c9270b2bcc5008182e6d592a5b4f99d3f71a0d3cfc5d105c6f42c3ab6597e53d043bda417cfaec68c6ad52e3be107dc3617df53724fb4619612b83881c54e35cdb1bf24a98b8a40d12712ea2056e2045fc96c5396258120919fa11911e9b26f84a397ab1882759a567c8c35055983ab0c75a18e8bf84d8aca6e95c09376d58fd731949da0b416834aed585d8e6331635bc701dd8eec77dcf6287124e7e0b5cfc2bb6c0e840ac41509de282d0e8f6c527b9066a504d6ea925816a0a5cce40a4d8a7f27701356d66fc0b5f252cd12becb77fe6aaa264914b41fa8661581e1ef1884e76669c0ad15892af29b21706bb2cdb06bc98bbd78c64b38e08bcf8e643cc4b3f73903bac73c5081cd12be58004b62ec3367c38fd6519b905781f0daca25674aac80c5cad3befd6bea8d7b1a2767f18b5b0f16e3e4fc208e92a8c56dcb609baf8585dee75e6aa71889654d71ec2a83bf7f02570c4fbcc1f0b29cef11b3efaa38c814e9e4ef0e9271f48f8bc6972fddb2d57f4f3ce3efefbcf83b0d59c435b91952df61df2352374ad9663c47e3b2d0b61b5ee996871a40bbb8e19603ff4c519590a9f79dc87ac336d01ee2a762a72b874c4e2b5c96ae28f4325b5121084dab19664976e9111e2902ba6407200a60b8e999a423ddd56e9fe3293fde58f841c5791e2ec8337c6fd2c259b4dd0f30dc190d2e8ecb76001dd673e85a6c832cb33e1e121d4d388fabd5b34e7c9f13a85a3e06851c1d8b526f4164fc3e522194822852d3ea825a409e6cec6b7dcbe47d2cc6e69d6e78bf4eb3d1b38c611794dbf3a60ea9c1db8a938bba378bdf2569ba4a61251f83d43333d0303a5488844719e1ee59b4a3bb09c78bbf407cf9711e3b72b2b19f2b55270fc2efc05ce49b5356fd1bdf32aa8be7ee0c4adda4c9db12d5dd6486f768ea7718a4f5753ed5d0ae372e97c6260022692b11204248bc073817b3f07eaf451d188266043b12819a389cee006f19e5f880e156cd8f63edf01db1a8032cf2ded6a2bf256a2ef979f582b95c84ca86c9bd9a097d4af98efdbbef83a157a11c0a5b622b663e5a44bd1bceb5cfa368c889207eac305fafd59dd11a24bbb4204a7f80a8135baa1bdb016a41da5301f429b4583afd09557f4754838e9bc82081e3d29550dfbf4631280fcda278ee79be37648ba45043c7a50db2e7e7765ef6604465ce00f062f5a6ec1fbf7d7d54ee5feed010a055bbdc842ba715d9dd52a1d8cf305a0403580d6ee639fd598e72ecf5d381a4c92752781964149ce6075d7aec4f9383254e244b3d6f0bd3f641a16d2c57e220b4bccc6bf651c9d07b5023161451861725fd4ca5d6e7ec00ae7f19a5050c83465e932025b986a809396e184673566bfe2c5c37fdbf078a704c35bc14a9b165f1c67097789c95473cb7d1d41648a14011b21c3031321b6a487bc97c893327f88a2eb67971e8f4e1fc7a6645e15971101c7c5dc08aa5a74daf4fb637783551ae57bbc89c49d5657507cbb2691175eb51bac1a659fbe6cc3f0d0c2091356ab410f1368ec1084fe638ded626f48378e7d6665464e01d425b4f8f74a0dddbd2d181811551d2745f4c50d9da8c5ddb2514647afedfddde19759e94c3f6d0f76342000d19224d1f39f29bac90c69a535e77231348e59cf27ba32463110a36de6076afaebceb7101194bb937a1d3e803c92ae70aa0d4e0b7b3cba4e54313f04baafcda9166d482a4de88d16b1b6f7860df01a5e838582da94eeda6945eea9bf2af08066e993d39e94ca6b676ac93dc95cac8507872b81895e0e5bde8aae431a00186623844446a589cd8464513bffbde461968e2c8b9c4d285779622fa21a7c9e84a3c7976b1e58bb0a90b7150cd3e479d81612840697b033c85c267c2928f5c9bbc6c6f35f179afb0e1784a18fae99023ee663a166db65bb86d9162aa7c42907d71d2a65c1b23315354ddd0b108e7db9f6cd13f4f88e732b4df4ff30e1019b80f060b443a2dc0dea20e2ceddad20255f216567db0731dd3a54f9faa8a5e5a2c20563076b7af74ca32e447c6a0e6fed1348e2c06b5bad4ac948f8a6ba143a674f4e222bd6bd78b29a957c1ac8a2db5604c22ea291efa2ef186d771f6e50370e734986e852a0201a78a683a857ef1668b7e17adacc94a270a057dc7c09e4f9eb478083ff9140dde74ce9b142d80b9c613e5129b04543b51e738720266d68542a6c450c1c7d7efe6207350a4a49c23134828170cf682095d0cb657a1fe072bf3e3a13efdab01e7878d3cd0a71505c9a9ec0882897ca61c7f9f186dd77c63e854963b0dc9d52daf4c0a5a6d49358e438c36d2f282c3980c93205756f6b33cd9af7d1e07ed8f70f4eb10e783d929e20fcea1975271d404c2b437ea38b918fb6e3e4bf9319fe2feda3b9248eb7ce644d871fb0eab794cf4650d2c9953c7716465f400ae28670c18c4ebc9f998c1693731d0a62e9a02b3bb488f8d0eedda5065eddc60c3d6d21ced5dd3e43d7a8d5a7929b69c732e940f16f0190ad5b841e67eda3fdea125a357fa5f516000b489d106d80e180970be7ac56f3a7b40100cad31bd8e58f690cd9195759717ae66495aca6453bce4faf5d59580f497e3841bb65aa3b4fc1624c60c68834148770bb49a5934fcfe483500c75e4020bea0ea816bf31755d4dd5d57b89a6e649551913c9277cde6c18a6a38ff3cf0bb41c22eb8a5b7044fd935d87386469c989c9dbab70ef8d3de6d04be4f11628aaa1b23c3bbc8273f5a473880ebfa669d67424272319a830c8cbe2fe178a1056c0626e67a212df8dbf24aae5b23f0324faa692a1c4b78bc6319e4a2d402d3eae984484822a3a594fbf368d130c28c0ceaecd446a90b920d718ac46b4d947daa5031622d031b375de492e7a26684d3a54a3b5b74017c73bf913fe2e8f259ac11f43c6523e31b7a6d990378e6b1398a8e8b4a8697d124c34d33af8ee21e3d1dd340c66b1c9968b3a91c3fa722fe29942f387634bb43dcba91df0708389075e76c069a9b5ff7a7bd8d7694280ec5cf28176764f389c18b8bf075345be0c36c47c4a7f3094c20268da525940cbfb2a077e0c7732308e97586de67da6a902803bad2f1d9dfe8b139cb47537447d33a34bc757c2bc3bf9f8ba58a719be627bbc0d365a7c295f1ddd072399dfc0c1d2041dc084941d3fd16655e841981aa68f9a77aa6260b7dae89725d5aedd9c1f79b2f4477106ceac61fc6949c8d9d041da40374fa9bb85d3db6572f1ab0a09ac9a53af14aab37c0fe493ea28ca0c5c9f97d9d2ee7adb5fcdab63f1b244e59128e57ec9fe476a41a3ebb62229ad61a4dd78ab851fed424d77a9e221cbcc7b462ba4e8979629473222f114d9edc15ed17d79223bf68ccdf59cd700df1bcf2df547dfb4f25fa4ddb22e88b75a7d1e62211d5b4de938331358743e8dd26d14c72c9ccdf709df057b2b15219cb3cc8765708cb0d2aab5e181c8589604726ca4456552fba780e54aedfd551b5f789f160994717f56f2bef7223551aa3aa4cfe00184a20832668df9e7619f3f5f60c2912a70160ebce091a0ca835c9e6acfaac2ceb77cfa6039ce679784a4c3cff15765ab277065b5d41f9bd3305e4cdb3524780207a68767bbfa8fd0fb5fd8ba2135942dd1994549d64c2231385668fe1bbf72970b0f1a2484ed1fc7e5f2cef66ed6bc24590a8a61d76b89ea8100548396574f8ac6c23d9192b9a5e0d50b3fff185f986fa936830d8f459a6db4ba5f7e0970926df7bf2acfa9d535031c4d7460ceec511df9de773078247f5704358b19b2afcaaeff0990d8a10dc91ae5bf89cc933c9cd1516c3310bc21f9dc9e007761b39e0f2584cdfe8597025ea949be223ba0d16e6f11685780a5f21a9fb1b414a80c9a1818bd96dd7b02a6a7e6aaab2f5b64f261278aad6d2c92fa85d352b9d57fab4f634142eae2f7000e32983c5280f515d01d89dd8c2cf98c50c9e4dcedb1b689673e13d7951f86c6e8996f3ed65efef6dd270c5ac82178cc9dc8e9661e69c7d149b7064a09bb233b333e1145b6d04b39372d7fa5338aaaf96baa950fec002e66699faf4de3e0079b61cfc9743d50278df24223bdd187f8382f9acab6cd929b681f8d948d8935d561d2b1c33e9b84b76d8cf40abe0cd45d742b94c4157aea915adf346d64b5169398bde4ccc69e74b3bd497804feda5f4b1c41577fc92ebbf91b22d679b65cdeaa738dd8649f65454b4a7d702ea210252dc820354046aafa317f61f9c810f8e57ad802fc4556ff7b6ac874ce5d03ebf3c3eaa92c418a88daf3dbf7a2b451e86d1c3bf86a22aa78b1dd87d94aa47545018be88fcdd6ddff4a9ea716abf5d3b47bfe6a1195d25de7a4588b14756cb85c676aea379b740183634c8cabc25bdfa54edbf4d48285ccf4dfeafb0b30537ea9682ed17dbd380a27369b1783c585f73bc91fb5e1d09bc75ea64245f7ede3f2ff32863bb7a369eada9d3b2199b751c3a77a7856341de21f877c672cc4bdada68ac0e0ea2990a01160c4ecb1673842309017e7a9420f5b6cd93e2fcf0016d3d672ff003d2479a1f9312df2bb753a9fdb77ce041f60fb7b53ba29a2a8d1fa1005e76991ada53ed868508121ab3aad3a0ec9e489e7369117f323afdb241e52a854e2c82f50937517eacc194ceb3e6c6858f29ff924eed3d44397fe6fd1e747954f7807f4e51470aa214728ba5c2dcaa03d2c63d76bb7269d6cd31eadb6a4137d564b44d81f2abd6c69ae7190904c26dc3e967d62cce11dee2b54c44fb35d41dfca4b2aad7a4e079a6495924b3afa9aa0487fa5efd99fb423c325efee11bbd35472ade7ea2ecac5a942b528fa4f6e8e4fc9177489d25f2d5c67bf1d5066ef24ccd8c571c92e8823982acb5dd43ba986f8b4ec05d29a990107cb06c8f9912b006e8f5ee5feea507ee87945a9dd4f9a00c2e75d0fb2e0df091cadd4e4ab42ae545aea3dfd197618c1bdfc5f412c03bf37214f9fe61e8d5691818378994ccd40f3010c5b11dd3487efde2494eff9511adb4c300936369b58559cc288a7564a1460f3ac26ce5026173b6ace4277162c8a1696f3bc211b63f7ff86355c220467fee35f02753407561b9017a8fcaba72a8e517431e0322134c6e2c6edac0c8618d5be0ca92eb3e23116cb406bda67c4c64514f1addb3614e7611640bd131264b993d031479ae4dbde1e97b1a91ead5ce4aa7054e337a4f2279c99397f82b58f1aa9ccaec73e16bcc198e72ed4ea45a31e4fd801c634e131e98ea596990c717d71b2d67c45a046797449364a5fbf30fe83ccf3d7412164d91107bdc2bb0759839973cea1da4dbf7951cac4fd585dcb039d63cad96c610ffe6e4784ff2aac8af5b078eccb5c4131e9dea99d9ac2012c6cf2f51cca7e0431848e2bc3feb60ece1207a5c111072a15f567d3fd709e3fe97c57a939686acdb959ee33fa7b6fc0af8bf8d0572712280cd50d79281b31657ee75fab053dabe57ea6b8e52908940961e0d19d52a1c46802146286bea1b07451af5e619b2f29451ddb62fc7c9ee908f7e80d134ef7df9b242882a4b97a5993cc39eef0bfb0ed12c567088e4a00c938a91638200b052e8c9a420a1e4ba978044cc57562a65e886c1f8b0d97964fcf623ad8acf642502b395dc914e5a41f3dd230d98179;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h988dace92024668f1a46b73819e2285f74bda1ec683c522e69d5a3efe661884d39c14d32671b8c2baee7d9821e43d8d7afa220cc08d291c4845c69d6c95004bbe40c4f2aef6f1a2c866ca2fa0e7080c8730edfdb2a2fe3e31474182c27567414e7f1284abcba59539bbf10955ffb599b39f0a8e553ba596b9fbfb047e6a2290ed68b41bb543c182215231b06b5f498be2b2ce60a40018230ab7f409734bdf20c5caf0faa9faca9e925d3d65ab7f79f61c1434c94e37f599a93e30d1b9beffd800dfaabe816844c91fdf6b72572f0302b0428e42180c7d57e787bd448ceab0afdb451ebd1db9ffd2918d89442cf44e5d26250ab5d11e26ca23adf4f30db61adfd1cf16626a2d3e38a400154735b2fee6b28ad4dcee0190f91d150256ca65b362fe26332e40db90189bcbd755333def2010ce5fbdb0ff716c179543d6cb9bd00e9ceaeb4c8984fa3c1448e59ca4db580a507c8edb0013537ebc3a5f5294453eb0bbda86d7d379d8ca41ec56339a5232432bc3dce0971a79f1434438a37dd0d999f3218f2d1ed9477bd81cb2de9790bc0655f37c0692ded97cf1c6846002d98777e73ce58a8192d5576e5315ac703eb3dd329c9e8494433ab44df75f1fca1f6a1d80a1c511c3247c426cb51057965c8a88a57672bd722a6572f6385e9870d5f567d490c35dfa1a0e850ae1791cec100ec0c48d3d50e82bddde7b26ea20b3abff05c328b4a9626f139b2248080db6bdeb697b9b95acad29ed3a2dd06adc05a4cfc6dec2d6d7ab265a130042f437217f249cb158effe6b0cdfbb7afd42fd9306e077617791a5ad1bc125de9a32a35407ff13b598bb0029855d613abb82114f30347bed5eaf6656801e159eb56ad3721df801fa4e5a40bcf10706a12342fc9e8f5f7abf6f4a8404deb1ce825f968faf7798f7655603b236f1abeba6850d9702275f3e7aee8cafbd292c78c17b615f9b028f0983e5ccd488a918ea4cc2873f390c25be9b337c8f0e403a04b305b8a494409c67c0c2aba0d4dd49d7652c52f94dc77feae246d6190b9fedc0f241a8e0b8e8c7253e6ff847f7cfc2e28c73e4b7ce223d8364246fedaff768741ca1c4f45ccfdbab597b4a62559a4e59dff7d3ce16116b8cb1d3138857ed54d81739b0f3c563d04c4ddda58a3289d1bae459dacfb4d401fe37c9fd0816af357c78ef5a20370dda2cc766bbd63af040f4fa8fa51d9dce72aa17fb19387f6f31581623ff718b72a466eb03af4de69137c12a9e8d26a2474ba1165ec6aaeac6423c83862e7153c9f6422e6fd91aa9725252e92c086ac54e69e94b665d4c298efe804a7a8806b633dd04d0ee0c82c0d49816207b5b4bf3587b68397ec66b759fafd81a3ebb16fb6b3cd37df2b1e5bc2455efa45a92ce719fcd57e2191ad277661851d075233531b1452e72b89225a1593dd44227887c3a770e7d750d92bcbcd4aaf180c8551850a7fb088de814f77dbe23b7c9998f2a4463108e6a332d394c4ac09cf8d37a35af7381b02a61b76e177195e5217cfb12f585bfc09b273f54a87eceb6c887ccd9ba4ab52f4275923ff030cc322201b2349214338e0bb0dbc906638e32847d2d7c7c9d91f9cf4ec884e7dbe0cdb10d6e7ee23de4c605c7f79bd0668483a35310ef317ed65a835e160efae176a8b570ace32598facf0c8e520a2818c36ae899a3dd557b3502a7b557c9a5b8ef30e63e213046de287adac1385953d210ae994c03791afc24cac8171f45daddaca01f76ba5582db49616a00016c2ea9d6453a14739b476880c8e9f9c4bc62ea8c97249142fb6bc7ad7ebbc91ca55bf7452d41488ec2964b63a1ae29cf4e7cda517b2a5ed96074527b729c80a6e30519254f54f62a9cbb7af771472b0b7d3202ca212fe56e1a86a06815733996dd194a49b81d771d7dd1c0e172f54b3889856d5485dfd07d4f3f5e271b96a39218ef3a682e7c7ca9db294b34313d8fb6ff743abb0225c728fcd7dea19a6345487a9b9c03d93cd65738c4c099dabd79ddfc6bbb580dd4d4247387325ba1cafbecf99db845ef2af4bbc3fa0f207af5e53e7b867bb8d953df98b34c6e7e615f9d6f2dfd0195c2ee02f530ca60379043d803a8989442d9c1b03f68d1edad5b0ae1e66561eb1d161aa0c83fb88310aaeb387408abef676af8a1a676edf7f3f01e2b23d362f94532eae95ba87324de7bd5509a862803c05595d17c28c1ae7309fb62ac5e3676ecc0959aa18300239b5fe399c45f49c8e78b84d7243f005e024881781c72c4681e562caf9afc6109add601a976d1a5a6a722599d0083c1912bbb666efe60dd56fceffbf4e0beb35b6b5dff7277282e1c6ff3ca6b3ae66bb9506b9f5080f9e6d0fac550b31940fd63dfe63f89ad17db6edb84b6d49355b407fc392d90ca5a2976466c47854abcea8cabd4ea42f908255c5745554361c0a84ce9304797aeca54ad22d511db756c2532125d404c14d493fb1ad03a7ee04b795b0c75800650ea6504ba846c775c5d0a34f2c22f91c6c4f1986a25e312a41ec9d0a3ea66bf1c956ee2f6a4cad6e7f15b86b4a9ff3f8f6e47e3549633376ad365a999f9b650b72d0e1520ce7f96bd85de5d91edff41fccbd9a4b797eef6ba567e17b061d74bd9da7cd105b30c7ecb3afd2a47a7e0a80c5f3c09d63a30ef13580e09b0b3351b82f3e4a13585d431d0b1a23bd820d6baa9d87d432dfde0ded8d23170214abd88a286bed18effa47e7fb8dcd0327e6295ad0a02339fced697ded059e83f062a28e14ed2d5e6a285a2bb333254120de00384b56f9bc46644ea7d5250599f6a31d7decb4864fafad2833bcfd3a3a23eeba50a0586e6bf1521493d8d82991049794db1de181bb339ec26d074bc3360a7939dd1746c956c9e3925b261924dc0fac44fcfc386005fa42abfd6e508f2a6041ca9aeb6de2073f475ef2a562eecbe89249f1fed1e74d5fa8f1104b23e997bb90a962a497fbb1d8eb7d748348981dcd24763167ec7be5b01e0d51fd4b9a8b6758fbee737f219733c880332058c5d2f097092a3a689b19df253e0dffd0325437b390fab99c65049133984a73fa2f1d70230d4a8d18efe02d6d496069ec508da9004d1d2649c6fc77c828f5edb4c3a8d0774134de3d6b280ad796659435f03271b3da6a1815cc5c36179853b8c20c2b0674edf6cba8217eaf8f7d3c5240dc139762bc69a01fbaf99513b80a6518ca1cc6cdd8c998aed3b97ed26ca53d18b6a409fe7edaece54686ad2624c570cdcde55f038601af8cfbc82cda9a9a313f18ee801c802df9570f8952f7b355c1fe4f0d23fae7ab35297e0af0adebb3e18e354b2c81c09085e967fd8bf25070cb6d33a0e08926269a83d0689d0993366448656f74744a5f7772beb251bf5f99452de9dc4dcb51531fa74649e7c29251851c6e37b291feadd9a3fed8d9ae4f4054d3cdbe15d99304d3f490641e65e0980ec64c4c9acaa56a7c2ab865b76375ccdcc30dcf6c9586772318ef94a8835954bb826fe973e58d0ef1544a6a1cefef0ff97feb2cd14627d2f4c1a81e6188d328f4af58cc12ef249d11525077b9c5b6752e26d75e8144846e646892452c94fb0c7b6860ded8a8427109e4b4d4325a71fa5b18f1cec085c96d2384a68e9aa480fc679e0ddfd9d77cb62cfa2b7fb1b7c30eec4f94695d2193a2d8e39d63a1ecd2fceddc5a9536921daa9b1b4de8e6bed20cb2873c04ea0e69500b21cf3bbd49142846894e91d373c90a8813845d4fdd6dd7b60ea6d69caeaeff68f45838f6e840345c8d094c17f6990c27760d7fb53637dc1f094baffc7b0cf13f9cf1cff1934469a5b95abac58bf7aceb5247e680988730dc969e48395e600cde752ccdc8b3c7fbe1dc3677b9a034c51ad2bb1bfe9b2b48c2f55803be81a48d4df09a43b6f83d7a197ff594d61bdd2716c3073c7fa457dc1f62ac0d6d64a1f4412d537419ec1503e55426e8725555654b03e582ec502afbb2628d6758278deed3dd93708ef3dc05080788547967c17a4217ee965e5f01b04e0a6d69653ff43585c94dbf0fcf45651a58325c4c71bca388232641d74d173bba739dbe9e3d74fae71db04b5d00d6222c3ee4f779a6a53a49d0306a040cae2f2c1c57d6883cef5989d3c88e50145eaca2903e2295523a8b435c8a4eda818c3e54478711f638306e251d71f809f4a380d674f3b4927377ff35610f4ef503a505b19535bcad294fd03205680d4f97ba3cbeb5aac628ef9ea63841e48bf04558742bc351c99c4891573b0b9ac022a75555ed45e1e96d989bc2d316f6374aa910f86d99cbdc2333e26fa103fa6f909f3b2c04a3c99da2268ccf5cfdf649868980bc8afb6ce085b9cdb64fdb106dc8a9c8839a603633e4537a965599b4d524da84aae4b43cfc8256a84b36f76715742514687d88b5caad38d350883dc249bf1ef06356639f33eaf8caa7e5cda52b117c389f42f6ce82da1ad6535dadcb6aad376a6cb3c8806639fa6744303591bab070f7af1f9732240a45f458288e65a9ca1c9520a2199547c7b4a9fe5c84b5530815a591e98920a470c3ef96e98f8f32c0ddea89eab4fadc4457c3be920b87e8e1fbc482c447602ac8219c9108a1d150ed8c007b76f72050605ab2b9a3b2df26b6be44683e0fd4f137a543a04143920764d4e8b7a294e4a03ad01159eaad9b255aa7bbbd35e5c9980830adfd9f9bd913cbb63201cdab0ea0274ef5915ef28ccfd70316a51146ce2aff10bb22cbaa7342c3243922aff0fae3b50d4c8935da90c97871a57667d85821a4605ded84830f7d0371390382c40ead1e99b2a7e23f94be5a7b519d6bbbfe5336d784fc0654febf39f1b1973e227e3f506b47446fdb00d8667ecd3624336d36c0f0b7e4900885eadaa490a4e5458dad404e483b8045ae8a4d12c953bc1aab97fcfed18746850700bfe97a8f571b0e5b1ec76cdecc6672e61e8119adc81eeff41b5bfbeb5b2828e7bfe82dd4b80adc0abab4809f764c52683987ac7b0b974e46bfa82501c346df92068dad346279de4223ae7df3239676cc96985c4f97120a8092769d90ef085cd5e363b57d1d11e04200eeb4551d31e1767ac5614776157cea8c0fbf9deb0ade491effc8185cc6d66264c49129f0642ffc71745ba0a92271a8f2246fc4b6848aeab98a39fd551c65b589ade23bf3d9c253a275a544e6582144252c46cc0ae6d0922721382b6563d3ab783668384b983b902e1ec74dd1f4622a01c068004f88fea5ee1ea9bf46e8a27c7e5a4c0e2249c9650bd3f43d980c7310d581177166f7b0e36c688a1ad0d6e2bcd36758cdc29f1415252b3f2725d3da8658aaa8c22114e46d6e4528f5cd3ec3cdb1c508a772b50c7646775a2a46e568c01a0b9f7aba9bfe98e377747b9914c04b791bb89ae81a75dbf0d131964ea53874b00c6d0f0549a20bd1ca9e5ab037b7721d6d66765346054c1a8af1addb9555203cb4a0fedd453853c7897b5958256bbcf741d2d7149dbffd2e62798d01f695da7d914d97ed7fc1a95c98b6c7ad28f4195ca27155b2aa7b7f9e4c912d025c8d7d8f6f3fdf391193c4f2ed2a6da1e630d8c5eecd7352e0f738d68fba772d59a66ed80144198df73c7def3fd88cd2e338342f9596e314312a7e3036b80d828e4ccf258abc341d71d21ca13c6bcf147d094ce1da5ed8373c230b95112b56f4165909b96abe53d05bee6f37a06d133eaa362bd68db6360d7aa1ac60dbc97cfd63467815010c877c154f2bd60698e7605a916235a754a338b14c4eb84d2cf34f36a65f73abb9d7c12991add23e2f65d1f33968f169;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8570fd0d934202ecc96c124708dfad1177ab63cae34d09f5b7e8bbffce8ef1e9231c2949a964b029599083c5dbde8bf3fbcaa7b0d0f8a2524f5826245ff25fa96e584c2651f09eaefc8adff3378eb1d5454981613b98d68fbff39ee676335c9ffdc8b5f062d0fb4ff32aeed5686307604314e9018a85bceb7f7e00c51577bfaa42fd3503b79a40705fdac6ff11e76a199df553d2d28d2440ebf6b7fcb29e991769c848ee66ae4956e1a209599fd98604e13831e8b099d884ba008e7df436953003de4ecf2df0974842f3e5c99aa153a763a09550e0034d7a8ae7691f5f49b0821b241784d3215d8deb84da03d49ae753374aae797143c6c3f5e5d9146e21980731e7c776354ea790463bce8f27afbf134e7734a13a88f55f316c24ef4888f637196e2f8b2c864f0ef20b3cf710c92530f7bcc12ab639d3dd95ba93f6e552b3a3e7b40e05f60dff76da783ee671fb70c4ead9d1b5b0fb9f639dde93417d3e70ac6c3068d00af510fe649d5e208dba58df514bd9596f2a9fcf0b844fc711544461bf11bd34c183b1ce4a13d160228dee86b7680674b25a90cd5cf46a6f1403dbcd84040876253ec6be31122708c9895399e1cde29128f1ac720a9003e4ac47bf7bb0d807c565acd629efc3d389304759eaf4bdf08ec1a307d67ede87741c37d856ea9fc2497699caa6ed3916a21fa1060fab65cd163c31a32439f247e3030741fa9706966aa854a5f639e92a749e2b374cefb217636cd6d7b0b6595166d14b6a06b1e0e6c385e2bdbb870c59e59f9747b7bcf34483a9416ab37a688cf320645fc439e670eda1996143484576e732c7cc3de49b317469630c3e73ab9bfd61e74202d90ac26aaf3c18a95541d47913808e9667fb41933b2530ba1c25a6cbfe1b6bc023e84b4d327bc39ceaf16f33b99afbc45e49f49b9f277b4d11b8ae08061e6ff28730eb941b5e3050c4064741add9ac724fd497372d1b331d0561f7b2794b4fb8e446f9a4fc019118c731c5b40d85f7e402882faa289a51e030fa3c8a56ae4165a64c6bba1208f1e0c698d9179646f7b2703ca5b67a07ee08a601134a63db67a23be9ecbdb3c12859e65f51f205cc333e9ece39608c9ca3699d1add4c14d791de8628c85eaa758dedb24354e809400cb7265a0103285927a4b3e7964b16f347747649208fc7dffaf593e34bff1f797a63527069725383ab2252f4fb658d50d17c28989402e4b2186d127f07574545527ac255630afa6ed00e4ae7cbdad71e8d1647f0faf3423bc48ed1f7d9d3719061568bb972a978803747e4e72de9d6771d443689073b5bdd68de8686eecdc209d51c3f9164bbae6cd01a0232b9afa3a1ca66b82cb98a5b8aab46f8199d56dad3d8185c926e508b48101660e567d5bb50f61679c3e1a37dce6473b4337d0c0484193cd36c0f6bc531b55ca906859febfae45583086630a40ceafa6e214e2ba66dc0d86990d379e7f83f85c8c902c6dec19ad6391fd20df136e99fbde669115cdc2c932ba912428e5d5a4cb2ec1992eef1a8b32a839ec4289b458f017c11d00f7ebceed9f7d2e24a211a66a113d86af11ffa8993949512af03f8eb8894acdea0c14d2403c7f37b0fbfe985ddaf8d383774a35ad282520d8bab1fe8fc507a31840f5c4e991d01a1bbf246896c609f7b95a604e88887ad1a93fe4164a696d0b64fe6eb35f02938c3fe906de4ae5e5613a48308b66f95405c1ecf880bd02b13967fc4922522c2a8054143567e8e05a877edb0cfda838dc32081db8b1af508d3af0341b4d626e80943386e57ed606a0b6d89b4e995462a7b1a9d648620f8a0025fd5afb2223b9529583f78cf5314368de78d68047e0d099e2a462e6d87e1a5bd2a4a6d109bb511ceb786ff9feb81d2d2ced71db555ec5493f64735f1659bbf3d38ee31b6d57b5d9b946fcd3daeb3f325e3f07733ba02c8d1f3d3967a4c295286b96d0d29df109123ea06de123f7714b27b8d92842f1fbf9c1e3cdfa2dea24f50db0f0c53d3d919a51ed5b1f488eb4a4da613eab8360114ad88549dc6b8df6ed215d0c96fbce197edf85a074dde08d0415db507f56c784ae96a50083b9f05716e13463b12af8833f2ec90d87d7cdd78fb1d6e0c9e2625ff3c46989ec70ac26fd57993f8b073718fe5267c5177bdf8b506d195b5ea0b1984b1b718c111658c3f2ace455efad8c9c149b47b2863f9f24a3a286ea8861866fffd73bef52b3e3894dd7a1b13508d778e080dcb0fd7fa85ead348fb8718f5d3ab08fbf5e65842aaec449449905f7936fc33515057d5c2d5f0b146dee5f335a2817a3c902975a10ac86476463bd5b30df4bc1915fa0b99f5c891838a6c4ad765e6cd3a1b6d47c398430dab55f0dfbadb51319bbd359538b9872cf3e024e5ab56dd07f8e3565f84d609698d6fc6466ecfe85638075e08fae4cf0400f406c1f173caf36fe23d1fd5e60c90a121905802da3ef40278f380fe7a04b52f64ddae1852c5ce5593c5d33f4edea7458433113233ffc1fae7397cc5c935ebc2e3cf52d225d842b89c21e3a784f8bda60038a61b6d88196e860c4c964681432dd0352e35d5eef709b533865b39ad705f8012f0a57ac6d255d9b1c6e78aaf833c81f08b6fe6845a825e2c4d1d51ba6767fa53cd15d739a755d641828d35c9e2aae719dc4017259ea945e07330e48390ccfce4165c99a46c75b9413de33a87d134fe8bc8fef5e84ecc97e0cb14b460a7949237f9eb052cde10c629c25320134154510943c78d651a164203b23fb26dfe26683f44a13241ef347da4ac28247d574fcf35cce4b9d217b2cf85206896d9376025194525766b7a798bb9dd2aa4a92f13e9be886ceea82d9cd4cfeeadc7040cfc458a451dca5124c599da1068b3d14d61cda711dfc2aa1e64740da66fae06e3ca916cd82d7e71fe26ca705e6edec2b5ffe363f32926a2ca010dbb6193e0ae42d23286e1daa9b558ed7e34b794a06e1088eaa85f308cf2152952a6a8c9eb044297dac397cbcba50fe44bf194f1777f87250ea65a47a41d446a9afcac2c998f8c28a030453d84fdc07339d3c1fe9c6e2ebaf82c85c502c5b68129ad3e6aaa00e77f168c1f1bf6c7b5dc64bc4233b8c355925381d7bf3612b27d9f42206d99675c38b9477c2199851e73ef464ce80ada61d75183374e4ea64434db2f58d8346090b73d140a0201b91b1cc70f0c5649595003fecf8bf366ec007e4491911fa3935ea64a5b1d88795cc39ff604c7b742caf18b7a1ea4229a8b4d174850529ed2e96712fb19ecb76a9c93736d74587d0afac2c3128afa1c0d9ff097650532cc4419e3b54581005d7c0edb9d8687455dc3509c4ee1037f3466b38a1f4defdd7d7b1d6d5ce3e186248fbcad0b722d39f0b897f9221b3660578d6133456b8bf2a0b7d8e44a01614cdf93fe2d2d62324ead3134afff18b4929c5d1a780a22938962eeac97550b765a5db01ac7ecf88f6516a33cff3cb1723c897b73d080cf2afeea8ed94d497815f380cb72b638f6bea676d05d351a22c4ca6441eb641e0a06ebf68de4c58655c7a21118764ae2f9f0a5b615e15ea6edc8c04179e23435c57bae8cfef9f76245aa2ef27d83162884e763950a375506546b7fa3cba77724bf051aeb6499449279f2fe1fc43ba7e88ed2ce127f35cd79655727ea3ab7753bb4bc0a317e1ebbd81466a0c742471960838499b55e89990a46fbf3c19fbf65f9c9a48d1f40ff5e0434129404fb0aed02a852c8336e9d2417e0f3b15f7bde5f5d97173d0246f1638b00e87ffa77f17d630ab4ef163710af32c1ed5b697057a55084a8a28e35f1a6bf0fcb840d42a790327145244b05f31ab888d570153013729a076a9c4b32bf9df0a0241ad071b95e128503781f461e554150105993bd739416e21045fea17056ebb68d7acab83805038a0970cf4fcd486d95eafc51f55c5e1a48a60743ad7810d3f61e3732f6639c4c0d3d329d2659b840a47a06750efe87be9220eaa57162f9d3b156223f91457c7e805044a0b7c446fe144e333524749669248526d0967555023f28712cd6529aadc26b33a5221e3301610369a0b96c926e811acf1561cc8eed110a97d7b414dce21cba5f1398f578325260b17620df3120502445ab41c094607b57b9a7a2821c7b76273659438e550bd5b9d23ad822238ba859965ed78b0f39aa30cf12067db761497cb7191c9812cb0867e47c9d886f6ceeba276690d3a18622196a1cd3536175068ad8dc37628cbfb94cb136fa103cf21b6c441c20531663abc4aae571b896fea4d4ff796c65f6ac1b34f6b4eab4f290db1dea26e2d7a6d0e68bcc861a0a11a78802ca7a9a08c527e6f990c7cd72224460a5b8c3d543045c3db96701f696a01bfa10c8f0f11e39663514ed0fd3a5032e94a695bb2a45e50499b0e0e8ea83086b967f5bb1fd69e4c645f61a1e2603a28decced24baffd95cfdd28f13c678d21f25f8848bac0880365ed64f1e933abc02b4d28afabeae781470262f4a6f6dd1cb156cf63111eaa3920b302fc02695eaaa8bb266e168ce39ad4f3ab6b63308f2705294853ed27e267ecef4c44e8360df89c2514f47b1e8d4b95e671ebf7ffe8bc6e095d4461665db8db73252fd89272c1d1ae22fcbb60282235b7455ab24fa4d5792543e867ef5a290d8ed0e3318d9e7710b5ca1ed82e7ebcb67a0d17c8fd4e739ff5fdee2e83811d346b583b201feb7cf7ee66fa813cda530344cbc5b0855daa0834202fa568564da1d73d737a05af99e3651ad7c0c416c75e1cfdad507a70ec39ff73afd6616499cb282de9ad4488d62907ce5896c09854585e211be4188a229ab2b873b24ddbb43ed27bb8eed93c7947843f5ed2fd335dccd5389e44cc83a064be3aba7674a53d272bcac273773b9ba384dfa33ffe744d75a911e1a0511c841cbbe9d6a127d8c1aa764902feda5f2fbc9391f391bda84b699ad757ec996208867039cf796c5573c97198d85d9f56bc10d17b02aa631fcbe18c2b86bb64e934c04cbc9faa4a55d530c2f6b6663298124afa3d7ddd12263f6145cddf71a2d2310f9941a882f08d6691c800621d188e1cb75fd6637064d363a5392d58601efd819d2b98ed075862f16cc205739141ffe00a30da7fef2443628006cd9b4add7f1e961adabf49d87b501496b42808bf0a4da149557169a5edd57fbd5b64785c9d989f293a3e61fe0cf17357c5f2e304bbd78a2a4aa207363835a2f7574f60043018a633f16fb5eef92b2d39df39f3b0921bdc1fb236dda92c2e96292723ff295e9f50c272d35659e6d283259a85100abbd5fd7154bd1a244e324ee48c9fdf99213bc4150f5a3d8249cc0e15c7aeb3da26742075d238a241c4e1b4951f0e028eb0adc5753fd060db2d2ed3c032d5aebdabde450d1efe21e6de1af4430eab6a351f97d58e8450619522a632665281cf5e9059821aa16b3fc899a43e5a319418658d9d404a95206c3d789d94e5ed5ec505f2a52c81569662e0b8ddf60fc5d2a6c9f11894f65ab0edaeb6c2f9231c1b466f89890aa3ad55287596b72d59a74c37ac2c5fa205f1a21c61db1c1a72a8f659a845e6009b811605b457d33d3f122084318216abe2f5c9635107f1acd8b166f6f3958796c60ff679e24fb25eb2713a6877573fe904f5abadf3303dfeb84267ed912f8e345efe502a1895b0c9b712062ce1a535312f6343ac1df93bdca234c7b3cd1df1b8336059b17a5b7dfc343129bcf019b1d897cf28c7bb0f0159d1af8c6b2fdde8b8fbb14e72883faf9473b86a8be305c3fae558cedcce19d9d16c59fcf4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf135c8bb679f6a0b3a826a102ec6e372388dfe52c9c9795dcddea8ae0f9dfa7e22afde6e42f6541bdca8b1d4d1a54ac394199e3ef4d7e42af76661866bf48ca432a21ecf8e128f41f4c85709cb99107451de99756c9fa427ff922b2f29627e6429dbe95f3c78c212411441c45635ecaa1648a7a67f4234c7989abc3200e099362ce5d2faca9049b492c9bcc4b0ee16d69f812f4697377c224f5b6eb71015b17d16a7254f2fb9da819ced4ff3224e45a77d539a71685265c7b12dbb03bfb81228dfa7eae1da43424a59844dc890078767f87ddad1edfab5999cc02665b9ec02c142fb8b4b92baaed89e704f0f73819ef5dde155ee04b7199c9e436c9ff9069162a52f56be350b7a06549d64c78d60360e969b60da1ffd8a4569ea84c6ba55557cc09d89108a3da3040eedaf8ee5795aa523a29ad6487372e6b2a49a1795f9c23afa6bf9e30d95eb60c5b2aabe3b8ee13cd2b6bb26001e5827edb99746093b8440255ac4fea1805111a6e39137fe542170907087d5050ec13f8d5ac10377d210ef20f0321203292d43abffda7a828c2302bb00faf2538d0e5acc899e308980b8e49ff8e67f1a6d1006d42c39101c646b50274e8aeb8621d185f176f1bfe250e33eaf1a06687b014ff685525051bb38b821c2fc8d26bf220de993e09d720e53bb544e8c4bb8699cb3a8d98b178c05b115c7bec84bf225c81d9539749d2145893b1031b8c07e4c6545f1982bc4ee30004f7fbd0b734dc6da0869fa267c6753dc2407cbe7feb6fe5ed91872f1ba1fc634def83bae878b77fe53b54f252b42abebb7997df82693d7bd04156753ee8688c52742df74096dd81a2b752cb59d88a5f52afbe85f67a5922595a2a61672d19bf71149d19e6184e9c6ad9e65ad7f8961ef54d47f26a130949ebe8fc0faaa6b015a317711461c34f293d008a7bc2dc5e161df0728f7b562b23946a865b5e48cc2fc674e92f09d3edc581d07ab8c043b5affe061d0055bd02f082632d071220188002320b5687883664addf2215dc074649f55e9e71e01d7a6c26ae4014e8f95433624b9172428e5c5f0c537040653b6f87e9a642897bcf3db9ef662844728ef27a387942dfe867fb590dd8147d44317e0db870cc731a16d6c81471c016d10009af713cd3a55a85644d0ea60c94327729668af47eb3580c3c9e91ced3ba73c19df501e175dbcda19d88830d9f118d94b6be40f57b841d14f3b9d345630bf4bb60ab65c4d1eb4fc20026a8263d508ce85473314449758b515173da989f68da46ee4f12567cbe8fe3539ef654f099961a5c4c4e9fa1ac2639d5fda51db71a3ee7145ce41291e45901ff016934a8737a0200f876e042a2e07bb10e8de5a1840de1d5751f63a286f06d31c18ffe67d5711b9cbab4e8f78e14a5b0648fc7acd6def3050656598ff5132e421879f9001c52782f9dcaff106cc51af06bbad338bf9c4d0816936874775532143751bab22c46a4e60662f6d4433b2ad50ab1a616ac68039dd940db1e98ba663330a49a0bd1da1d827ac38020d8d587ab7cc3bae461ea7d01ab50ecdd64b22b6691f9089fc60ed3a935af0a974d85a89ff206d997385b5185f8d2ba0480365c8f2f6e06c6b684f6944e4b6d57eebfd1ecdd73c4955dabf559ef4a73d55a698c6e6c5a6a05b67bca09ce5854cf46b48ecff081a172cf7a169c863dcc3f7221c4f68eac7ad5797e3585c456cb56ee079fed34f9d25ec5e7b6bc0c3ce1a9e547639b6582daf10cb3bdd2145a6aac036024dadac125dabe7fd3178f9aedd0342ab1551d9539eb99173d8719818b52dccd9fd8a303f0b236233da173d31bc9214fdb76650a514a44b227ad08b5c3a4dd0cd406f937ba54320976ec75d0036886deba09e967deae73b765a03bc8caea6933588dcca67a11b10a1bf68c48c4ef9160373f86264e6e18bb10ed02ee8f90104f7a3704159d508b4af576afdfc50354516604669bc4a45529d52cdd9c369a7fc948c2d2c2a7074f8007dd05df0ee99e61b0c679e3822438307fdd1ef6d802a9ed67b18490dfc805876519def71e3eb11dbecd8c44333d955fc7a3dd49330259f8ee2637958c2b0435958dc76cc01d6fd3b768fb95db8fe348c81e5a9f0ab5b4ea8b09efb537777d7ddd72e04b402d975656a59d51a6e0365e9d4c4f742cd3552897b1c22c97502bdc5720f01f8072f3155e527eeef8d56946a16de667fab6864f168c16b3f3bbcec9e335afbb8737c5b8f038075a70a4973acdf4c0bc734469022357b749a64f943c6c46704157697ca6fda1d62c2d61a19f63e3763368a1f7559bdf9e38e52b307df2f4cc471dc19383dc0c62692f2e0fc64f189359fc5826b1f34ec06cd5d50d51ec7a76527ecbe705338c80a2a1a7d07a573d4761cd10c7b58d82b48c555983ac9e55398139c18eef37773908aaee06a550558d8d482f318795287748890942114e231cd2c5ec295c8f3f84ba50f503e226a2780ebf3d894e099b12e060edb6d64285fb41f2e0dfcf11759070a7e813b618dbd75a408f70a4ee71b2de3b6abe25ad38c765966dc5ff62f9e6ad01a3de7d13a97c17afa653077a07467f163fe43ea0e45d96ab2a8183a0f5e80dc065128cf0e37742e31227960744cc4bbb4f1e0ad629737f1492b21d825e14f8f36f949ef938db908ee957d9b675c04c5ed4054845fb7658325652322a05c8fcd1b5c55040bcdb81880ccd3cfe8823c8932262bf835aa146049183904c658eae9de87d620c53514cb7e56871bff385c03d4b1830e7332c826f9c8c7f68cb4d6132c1b510a62689cf7aa083aa348f93582e9e9cbdfb53046da45ec1fa60c7c5dabc713644dc8b38e5cebbc05939b12c453615715b4f0ac9e9b5174f8a5bcfacf43fe11474f5d94de544b95db1f810e89cf668694c3a7fd2a3dbc8a4d1c690eb741171932a68da87b61af42d5a3253fb4670f66eb8904d27290f8cc7578ecbe7de4f905ed5914cdbd5c9429d15fe4f82caca8af95fa70a354d6eadd566bd8da0c5fa1985fa470711da768801f8937ea3d7ec3f33f34daaee2ef117a38388a391a20c674d8f3ea9898aabc7116fc3a41f57396e816cb31282a8044c95dc3cb3e8f7c6cbc1766089e90dfc93093e00fb534bbe16c28aed880c66ec72025f68fac44b9082386e6f323ceb36d40e458613f36a07050356589e1d66793c8b3c6450b9ee4f13ae63654036e956eb5e4e4dc248c24dd44e3ffccc69b4e6b70a2b863aa0da952130df3b3e63fc301f81636f1dc7d7684c8c1c6e7786d35dc00dca5960cecf738fea6c58b06040d7132117f4d8d423fe616ffd18be0c50f652cf33d191d0e62e30f2a3389c8ae7dc9340cf939bf649cbf191f43e97eb81d7161b6b0e132300d1f6d2ab89185b21502212b795190aeb2181af02284280173d62c437780bdbcbbcea112e0e4247d413cefb2240b5a060ce3a9d7dcbee395227798f426937db56460c66cabfa2214bcd6d971283b4e29945d65a906c5cb4be280a8d5dc35d19cca9938b49a402165f003aa49f7554dce8cfa45af076bb4ecc64f0ac73f27de0d7cea3e3c988f6c190db920dce5f5d93b37be72244295a942bd784d9e73aba830fee04f8bbcd8fafcb73f29f0a0f4e02f463c6e515a7bc0ee5267cb4f079496a037fda0fdab10afc6c5338d4f9baac084afd2fb02307b80ad96dd0a551c112f1d0c478356fe95f803babdc0b6ab741d9e42f53b06ace5a71fe7f11d27b9d50ececf669835eafe22936d52a3c9bb3db5a4dc3d9edee8f26260da132f73ebda460382aa519d12c492da85f4d32e09b613522609c749f0494319233616beac8d5f27d2d2fc05f6065fcbea1fe9be1881c48c783541727e0334e69e5f061964ac685942e25f5b7e4428b46655d9a5a83ec0159ce77e02a94c5a055112ef018358798ee223bf7ed6374753359edf537f4db23c6dcbfa3c3510b74607f6a47a94665cde612674276bf828e2ab9e10c83df2f2bc036ae39ba807ccd60154846095d8962115b432ea6d36cf5b61d29d85320919347890e0a10408c81c05a18ac6f5d4f3047276db2fa0ea2c42ce2b1c36b668f06d460266124197eb8a0ba59323a453230422f52af171eb26ccea6091e0db27a797b6df7b1200ffaf6ccc2985763b0ca90a8232ce349b2f1d5d21f58dfd986cdf8e1b1509475d4464bd536b438bf8e5b9e91d65538485951520eb32413aeca11a8f245e36ec76f2364e9dbf6619daae5b43b1df99e19a8840b10beda6eae78012ab236977a7b43e3d2b97303fc825664539e05d28fef4511bd3605a24ff46e3c30cd5921ef8178bdc70bcd7020dd89cc9bdb3d3f0482457cdcdc7105776d8bb7f226e52bdfedb92a00f3760203e3d3c40a1bcf0cc0514c8e7074ca3167abab5074c644d051ae6a640d3ac806568fe5bd3e17e4769f77a996eb3c8c370db96b5bfce7434ee6d572d4f6503e53ac13b988d879de4458c6e4c190ab7e7c18014949cf220d03d6daf3ef0c257584327c05b6541ac924cc5263746c7d6efb15b58f5aa02fd34555f6ee68aacf43cc12f04caebd043e699f21bae418fbf8a0a3d4a28828f234baa4d22754d84f1bb8840b7485b4c57165eaf433822f079e8b169f599c6c8f0ff88c5633f13dee6fd178293b5891a9a9f4af5810cbb7e39fbcbff109e287f97bc8fa478b60bac39841112dad7ce62c355d89690d9e823ad4eaa3dc68ca7827029456def85be9c90ecfd5c3fcaaa75fc0d0ada550c1a24122343a8bbca2e857d7fefcca6b514095f209a0a7e29c6a7d5cec944fa17f6d633d61bfea603306619021471992ca1742d457ee6cc88d3827100b63d853601ee54a9d577da064af85ac002646fb66205124523ecc523388a34f26c7599e32d230820f2f9473653c1c1b20d79af134dc415e15fc242c17754c6c65df60f308ce7cd07c5d3bdf5c802ed2733ced24c254ffdfcb04453ca0b4e37dd705265660df0e65dd306da787038e59a90e66262e605730f09bc20be3b08e83b5d1cde0803b9f9bb796c1a2596621e281b0b6b94f5f535f7dc45dfd87b49a23600958279b64ffe88994201ef74041b0f7a726d7e44a2f7f138b75117b2b8b6d83c43cc1604d2c434b8f4cb094ad10b5d46d9573b56eea8d3607df6d23ff6ad00cfea52a72556f86374f1df221767cd6a63dbfae6df06c26fe673020ce9dec752e10575451e965592cddecfbe2e26fb6ccdce8d08fc66db60c6b5a2a37dabae45a1a6ae9963e1d90ac67e437a699a125b61674ad05221c20f2773d2ce4cb9a47b6ddfbcabe3f6dfbdb4c942c43487b730642f7de7d4e9c316e56965f52189c45e06bb896051cc6572ce31703b12a1bfa0cb7eb223fc11c5a99758af80d3abcfe3a5ea3b7ccfd8b3e00ebb7d2063a56b055f21db2e86a664626d26ac675df77eae1a10df1d6823340eea7eea78cd90583fcb63fd7d7ba42f7d4e248d2cc469ea3e9fa841e6e556e118434e3adcc32f250f406e2825875bd92971db763e3120ed6148dfb035ced0cdcf900cd424d859a41769fb5f5a2f3469461ce5c83213eb5b3e2b4c395e73db4367d479661a25f96ea303d7f5d10d4594c5d36a6d383b39564f5f19cf103ae23d9e66af588b1cfbd69bfbddafeb949b107b91fcf3641c9ef6d851ecd51bc1fced06030baae284e7e8ad61da55b1ec101d2c932598a3c89e5cea992cf42ebeb048c5808c8d960a35af2ddcb856e39882eb460428033b2a4b9a5ac216863e3e0bb9d7a1dd3b3417110b3b1d09b19051256cc40ecf058187e30aff9ebcf2d05e69c750;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5f9ec71c3790cbe47baee04dd8da4fe615178d84997efcf83dfb16e6f3e04cbbcef9ca8edb97b4e62f1d9f4b6b037e41d2f8a28eefdeffe69781414e099f12b1c5ec65abb75c2244c258e9a25e7874092c2919da1b757463a6f544a4356d42f157859a2b7ef94ed13454c5c3d46ffb1db4e650e6a34b509308840a76c5e43b9acc7e849a947a0b2f2504168ad0e69590c6ec59f42f2914d452433380855b9fb712541b1745a6fff976b714a27505e8e838a5284c354b862fa728076342a4fed911e0301bcb0b051d117e8a220442bfb59fd2b366e28216557011ef20df3af9b953b6764a2b7d15bc24b934448c61804f0e98a0edf5e512cfcb3e6c4270184ea8e7a98ca9cf726172f1c36ebcb82f45b9545136be2968a2bbe807c3b9a70fd345d488f6e5e0f4b12caefc98174c52dbfb14d8edbfc5fad32e30da32a99581bb95213588b84c39875c42b7465fd05bec60ba73ebc1b7057183cc5e9133c28588136a4d1ef3e8cee14030ecd76997f69039e3c10e233cf76a3d078c73aec6e5dc9b65ae35593477e58ad4cf648b964afa240410c9bd463ad9a711a85f1608fa5f9c0fa7bb96c692c136a9b58f95e89041c9a097f7e86eeae1a6822c4012901c90a3dcd0c73ed08fe73e60c16d0cd662b274740b92c8033b04061d79304c757ab2a41d21af53e72d8381efe6335a449aa3ff75f8e60df9dde16b853139647b16a27acade4c675d3fd7fd7df60d376b2d9b4e6397bf8b1a491963a5d32314499050d64d100cf5ddb494846568f57bd18834359a28bef5fc96d3ed83ad26f8da672c3263dd37deacdb61500f3d13d61a56ab892a997bbd574e90884e9bf761b0190cbeb39c12f3e17389c74e8c69fbc0c619efed30e4e5572d7eaf41a3b7e20960e31d1379d4b3397bf15fbda09d65d1a588982af09a54b69b30e8a936545a8256042ea134096e8222d525d3b6a474b047746da313c2bd736acdd653cf0e39bb08e2563038eb263eeb9fdbfdb07716cc4742ae7561861b599347ab52672f434cf5619e0cb1de046d83deb8c905ffeebadab4b060c1133918f1b0e37cbd3f373a920f2efb84d9205e46716579377a8ff9b42746cd77e7c55b5626dd71d3f3731ca281185bb77e34a9a1d670b3669e7bf16aa6364c3b5320a3fc3f91f13f9bcceb78f2e2b0498827aa2e7e6819336051662c7917ad20707dfb684a7e7281de538424a7a0d15f957c86f38a8d874acb910b9b694297c763caf316f21d56506f1f2185dfa7589cd4ba64d36986feeffea680e81012b7a5b10173147f04d4b72f0a2b25b0181ed3eabec8e08b65e13a9422894359aa0aef75237189f67281692d0e07b24faaa69cfa9718b5aa798c06a3f2369bb2924004ff4497e947245b4f9631391c37111b435532bdb3c6943da0e8e00934edcef12f861ae16f703ef621a47ae7b054ecc6bb2e28f3fe042c07a552e9724e5b47febb378822c15b2632791d916f5f3227b446be7c90367ad8200462f21d888bb306100da6e7aeb835b0866ed637894dbb142e1c5fd25cd259fade948a1c308c30b791c09eb14eccbe6c804202b44c00ac1719ceefccb3b988cd3dba6bb17ffd5997c77d3c472abf514add0cc4b132dff09c2d67470042c5675973c4a4f7f8c18a983b5cda3077f98826d8715a30085876b0fed22185d2e4fd3af0349ff08ffde53c1a4d30a6505b1836d0bd8fb5896b9b5f0394fa71c001e0f7c3e4015089237a5bffe1eca7209d80983b7c3ed00155d7592b87a08d9f516810197e9746d776d4ed5a12ed3e52359345bd25c58c564c85e3551a8961eb01840dede1ee1ead5a6aa16abe6cb7c38d23ea5c7560d4b6bc02fd549d6dbed7d8fba0c9ed697bbd403ae117d66be0d2f3e21b88cc0a7b18b2128700ecbbdbe33254a5bd9eb728114a725056a90b5d0627b25eb1e24e83df49e2115ccad99579084e0a76898d9000e974823520ad1b2878960f684aa0e3c010e0b9c0518ed6969056b8029314804dca0f76c868a58bd255b8819b7ba1de3a6ad0f783ee426a2ecf026ad0876fc3f432d8cd84fb36feb57efe2bc57fa9e237b657e986097527d5a5ad2b50a74e3c689f25c16a429fed8d08b825ce575bc3fe7e238803dbcbc44d450d6f7508cd1aa907bb19d37d7a48bf72c5afa52f9dfc4082f46d0d06b2f323a19bd6a0ca908e16d7e75c430630cd1d1755eaf02bf061c49e1b03577068fc65688b28a5244116e74de447aa44c9e5850b71a273ebb96df1fb5642f03602ad487dce305f3a0e294ab3e51058b42c6e604685bc0a7b25f42e718306e6e33c99a2e878b68a0246f1ec4d44a16c98e9271535eb9dcf2a975a74f84ed99e6c4a91eea9f6194af9925912fccd646ff9ce506af2a7b58bcb7b86ead8ec853b9c94d1c15f3806976bc8156c82c2bf8ad6951ed285f0e4cf8e404c8619587e819d3854354492e3aa8385cb199f3020985d0103065e07479da0ef3ae80f4a8c249ea842eea231c21be07ee143ace44f343c5aeca8441b6e140ae6e97a176b2041b5304e43e2883cbe65202b103f28ddba98b2a968b9ce4c20b92a4436c0fec9ab98efcf142ca921f842a6661815c75bc8d26a77efcef4802823fc755e091911d66bddf811265db0cea394067e497ea7dd7273722f465b232a04194de91631af4a5bd9c5d33782196e8136a0c23d55f329334081cea53366554b211a0d2e4535ea735374daaffab38ea6d9c06b64da4a16a7c31647f71daad9e0024262c75a49bea63047627e16d4a93ebbcb3e14b0dffb02737d0b01dcbeb6961359e635dfa4a6e36f7117f9779fa5dbda8144443c6324032f2259cd5d892a7d6b5c6ca2c0f3a8cc532d48ad159dfb4b638f8a04d9cd7869e20662d2c9deca6a588bf200d58c9a58fd67919c4be7e8bb97055d2909fa7c3e6fb59a07809519a7f9a463963a16e00d868a687215fc6afd321fa4e6dda2c91bc9702d3bf117d1b0ff5f4098e35cbfe2a70a2eab8f136d58722df7ba7392f0b5cf019ce95d925ead57f2466dda9a87b8f394840ef5164854a065d205797867e06484471b879e042705aa8be0912e772376bbefb9b6ea8fc06b749e027018f97cda12a7528358caca08ff776dd85bc2383f3520884e2afc7c9b38014094abed470d18e2f164bba0d1632f2340509f4e94a1597955e72e6cabbec0d2e217b2cbc37504ce37175e2126763211e694a5895fc05f3c68908d86c77d5596ab328c6a963fb80068992e0e640e75e40224c0bb51e2909d081949d1f8da04c899c15ad35d6eca9b98d51a8e95a005e35411eabd5ad0020f165c3ed994ccf32306cfa5cda62303509c9a5b9b6052428154ecebe8fb1dd302416ca0e4cb3318fcb7cf42faec28f7ba391031b33c54e89120f484281b6dec2ca9cabf2a72c021f66dac4fb4cbf04cfbf5d585dd28ecd548ff16665f2bb00664a01def95d6b429cca1e4691bf321ca590a13b932c5399ccc584a4666aa8b38909300c46b48d4e32852506d7c2aae2746f154a4048d973bf8ff4bdb910827eca3e26794cff2ce66146d249205014961607bc1782f0d556e9cb7a11b0bf6f4cf0056f8d2c3d5093fc7cd9c62e7f4e857377e39f8b3bfe78fcf14ba2f647b6675bae328e5786d264018c50aac0031b898094e413b1e1f90d6395f0f9c64a87608b530ca322f30f199953f4942b1ffb08684c0a91040d4578e6671a995d39949e6e51b10111dc78ad14fefbfd419de619dedf6e274e9a71e426be5bd4ab806580d5420e41b6d3267ba97b9ce15e0ebb8216b7b15bacb0cba66fcdf934f12e41c0c444e315ad4b9a80576b914a0f858952f34784c403f2e3b7e843af0182e23d6fce769db9f5d7d9fc6d6e35b16fa204a6d10b522d2c5669c662038e62abc20dacd66c7f8ab07356e106f52b4ac419e7c8a5eebf53498ce7f2d29eddad80f03cc15aec43029742bf54f973f84bd9c8732cbcaffecee77d686f7361805e3db5c67afe6371f93c362fd3d38af493e053c50534d1f0460ab3f6c3b9449e7570538d071dd0f5c8c994b7baf5b39431dfbb2d5ec8bbc5719c62a9ec653c2e0b3cef0b199004c04244a8b02cea94114b42c68a8dcd95d52c51c1aa6031f6793b402a8f9b013b94b36268d11ca452e310885ec7d5e6a6e71e80e44fbf818456c6fe3276c7f44dfce0b6f8fd44043862f8cddf5bb8d02154499c5e63770e83d65df1f2992dc66a166a2a09ffd75e3583fe6eef9ed174246f48be60a2e46d893bcca5b78dc4b6eda5664d88ca14a2bd6ea36b42599ae73fd4e3a595944cfcc985aef5e56ab3d2a443c88972028e5fa35b55ece13180d1f9c501f6cbb2ba55d457bc79063238442a494efa68e13623824004d5919e4ab3152ffc0439cd2a379b446f536da74d893d2533a1b9cc142ab7e234ef4ef16f9bc125ce958ff2d5c93b7298ec55ef3b516f968dfb43684c37e9f5aca3e9a69871673cf537452fac92ff9a4c2c898bd6d6c345a560299a0f8f19a8992e41a4f7508d7ee0753fdcea72e8ff59788bed5fe9195792f15bb671ef280b808324d8b494650d6ac385280384dc53d8d53c0934e36921d988a88f593f656db60b933cafdf416c57adba8a3ef74694dbdd782b61c25f8f720fea7c9f7f7cff3dc8dfe060348a0de5fc316cbb834d39e467b935306fde160cb1790e8414f346f44bdc842508a8388c246053751c527e473cbbc698623682d3a945e1f3150f85f2c19180c1f321e3ed10d2af2dd252464fd6ef704cc836bc4794bcb4e55e3aaf6f33540af34126a31077850de33ad1388c67e865018d2aa2684df1fa221bc0959547fc797576bb75fe2e032383b2907dd3a13d79cf7bb43ba27eaf1631d501279a7b79a1ca8388914ca69d058d5e230480c125fb78a36565991d1203bb9f5f0e060c66c1ab1da53cc3f0fc8b5d763d8c53603b36494074b82aad2804865204cf4b66209000b6f0db40707f5b50ae2d6b55ff27ec5c95e9add909c3d7586a77ee0d947b0c35592a9e6394cab91ed70206bb411c0a7eff63a271bc6872f57d8ca7f4a5c1d2682204d9063d469b3f69b1d465e89c5f2738f529d72ad2d91cc8dc07219dc765ed79249bcbf8b6d34bde6864e327cd7bcef7e7e353ed49d7ec1fd4625a735c3cc8222ac231df3d64c9792e7c0fb4cd54fed5ab2f8d96880cc19101c3a5f85c7369e75f74880dd540ec9be263b9c01386526d50814fa449e8a00d678ad5a6c7b80207281e3d5d85157f398680f4ba7682ff8a7772dd687d010724b08a379705068e6e959e09dd544ac7f256707eeb75149e78959ff92b5e974ec681798ddb199267d573b9b7e5c0e34792cefdc7beda1dc8d88120f8a015a767a5a4662d70b31fa1cde80c681983663e9934b3c76def3550203849d84a25a06735fe53a8508700aeac49a00a09b23d73b4b0b71bfbf1239a91cb22d3c5c64077094b8b81e9a5a8588c70eca738cec63b99ff5c64fa79202e625ab9bf81661653addaadf42c5dc82b09ea62e966d1a6698b96134f3842aa03d03a19dc16859e546382b721c589af1a730ab7dca64fd432d169a1caaada58bd980244a0dcd98c37426fdadcf1ce13d3cdefe5eca8239818042a6cb16106e189f42768a5305d74e1606442a9af1ee5637fa9e3f2eeafe97610659e779e2a6ec78f78e4af7f6a66801be4b69ef1cd7dc3810d6f79a8dd55b9112491a0e54db7c308cd94ab779e362c2e6350b2b5457c6a27e3bdd926b7bd21a8bf2ffea9415e2ace88cf369daebf339d3d55855ae5f4c2a0937c4c53d6ef23e4630af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h73f1eabe3062f470849f23a2b0264572df31aa6bb5ed7d841b817a66938ceebadffe17ef1faa67d7b499e7997bc93d79e54de96fff2b1a0e4fdc3972ca386174a82ef5be0f1a6879ae927005674685227470ad3d70a49208b0cf21e8b5663b956d03f3c2d3e5e830f8203c170726f8222242bbfc00450ffb0437654336a12eaecfa5424a04e46ff01bec3f56ad9d1a1448feb2e5d52931fbc62048912cb83129daa09d28d453cdfcc58c9866e8c6d0df8fdbf8aeb1e4887b4f0eb57ba24f51a1244df210eaceff4fc60c1680c171f0b6288bcc64e5a0e85f1ffbdae42da110d1df19804ca7503a37c1f399579b9b372768636844756085cfe155bc9c22daaf63544eb02e8e156fa55cc111e577bdf77793cf5d1857ae8e861241078d871f91196298961c1013719d36e8e5417b67471312ef6502b1260f1cc0611d999358c7a07d3083f60cb40220d8ee1ad53ade80edd832a443a5421d669d23d2eb850e21a8d8b21bf951b3de42d10c56148fcfa7912c6f13c61641620738b96dabb55b4d8fdc0895ac8903d8a14920f2ae654d2fbc9c6f0647f0e63f6132682db8a89afb183ddb6acbb32a7248c91c40eb9d9efbfdd809f95eb17867b67ecdda2b008e53c2651b6eab2298890da32caef9c9daae6392011e041fe7a145ffa693497aa20a113c88ff28646d49c498085c6564e48c3aff4ea9742a08612efee747340f1d148f45e342fb7e8d17c5e82c936df17620029fb17397fda47d1ab6134dfc979415b6a72e00a9bc264af9c4feaf8cd95bdd5311d7576e4e16d9607f295a6decdb258d083684cf6afaba1f29543bf4a7a9e2cc48be088c878e640a0efe6be302189c23732a027a5dbc7cd25493cf71fe877be2bf3442527c6d25f5cab655ab27616220c8ced6100301cafec2871691da538ac93395e12de36a6a575aa085435021921fbf6579ef995a565bff67aa3d66a7de164b1461391bb7ec269712a1322bb670c176b6ace76a5c3fb4047cee840fd3d945631d3060e7eab9c20da929b3cc11cf25441511d250f09b25c83b68b8b59b9c29e64b326c2886ab331950f3b15a128062725d47aae7ca09768370afe0f528b7359d703b6fa742bbe44e6019a8ca10125ee5947aa4edbd95c4f45724ddedede788c7c04c2427886d8b251da767f1bb80caa6c66e4a095884301f0f0fa5af262339c072a9e330757995786505d0c6d50702d38a7bd140962f0bb968bcceb82807a00c0f0404f5ea56c429f1132de7f8a47d31a48eac1675b1fefffc40d4ff792fd15cc4f41ae59dff3f195563e292228e8165c9d88e0720917f4eb6c8ee49160fc1425db4bf45069f9626f35ad2fe2e672116f4745f5613dd0bd59c225e1661ebf1a567cb296e62c74b1eb068e8a104085cf1694c783cca2f2cff0ca541e4feb90605fab7c5f9620e1af9ef45c584e6897710e1abd2e4252a26a060fe6f6b81857e5f8130c8e3844afc65461764f9228034e627894638c38d10877acb52ebadf55a0e340d5a273cd8f4b42a187bc751347b69e505a9e57c750da0d79397d10b6d7d4fa6ad3b780a3b30c02391e077084bf5a4fab8642fb1eeae72e8dbad9fa65bd8757e38b40a946c09a5cd8390ad44061f5a70ce118f60eafb7b779a6b105f083c52a3904920d721964241289fe618cf20ce5df0cbdd4d452223ec2e194719058213fe38d476cb2d2e4968f7de0639e1dbdd4201bd495127b90a2c13d7707c028d5fab15d59dde0af65dd9a773a3c169de6bfa3e64098c97620763a5c550079af5d61956181fdf09a8939d11449b48bf74b50965515ee9227df5a02682fa7d546a862797db6108c835bdaedc728927c5dd1ac37fa04c0e4b6a9e9c5622e92155004a0f7e19ba4bafe742130c8aac721259a489ddc9513ea3c353b963b9d12004510ce99409e0910c00c84a2159b2e18d3ed1fd16185d57909cc017bb478fbbccdb3ca448de858b283f6b247841321b32bdbbe34a5c0d2323c8d39a53619567b3b95fade72e389708ae6d3a5df59ff85bb59c24521ff430cc424b31cb7e7ac361468c0400ab85052f5be15a889529d6efc091e72a794889d3fefe9b015587afe591bce56ed2cf4b7422514192e09390bff00145824e4f600da7be512242c7a0129f3b91bd8c02fbe82d0f2ee0600b71de8e0f99ea49748bf39bd5284a8dad488c238d5401ed832c16430054577af71f7fa6f86cb8a1b11c26100cab7a35c4a88ccc566023a205f3a4677e642ffb229ee36fa12dac10d222ab7dadd9f83159c65495c0472f711009ece59e73ecf7a8c1d0c95bbb2477ca63993ce4e408472cf93c07e7e84891e7325fa0895c442d40a98a016c91d88b325ea75d999b27c319bec431be720371c7263ead519e03e6762ace28a59aa86b6f816a5cae1f056abdbf64994f6a44c94dadb6ee50dc974bdfd72fac4cdb1580548ca4dfefa524f669084208bae688c9f5d4a7de3e417d479a783319d6a6f4859d3488256c2b6ad7ae40d648f2172715e9ce21d9b8da0040a9c1e8c6b64634806cdd580337e1827a38e7fa9b36b83c898a7bcda090359cd1c4b74199cf98cd2696516e4bf448a1c2acc9b03426541e17af57284f3ece40fca038b5925c09399f6308847e0780ae0bbea2902df9129c2dd9e1deb501a381621b4dff712df25b036b4b70110574dcdcb0aa1192c379c9f59c9cfc776c01eee54e1acc75ef37c493a155988f62cc132a9fcdf1e77973026c0127bece400c41214439d21893fc382a834b1bc018d5b3231ac5700648d2f440fe40f459ba6cd0ec7066baab0c2c4cf001fcd8d488b34959f2031f40b39c4bca93144b4dfda6c7766d4d5afc6b5eda3b651f5fd3feba7e3ed219347557d2406d1022388f95aeb78f3364a1009496f9bc83d6f2979de8ed24e4859181075032cefc07190f53938d152613e1a9d0db5bc2c9ffbc963c631fc2af7b73efd55b8b848852f4a47055ef3451101853ffa8fb59b5a78f3928d25a05f4966d4b5b48b87cae7399ee5df5a7f1273eeef2bb57485192ca448d604b72b5cb4fe08533ddb24c9502f49fbd215a600cce019df3cbf6c1eac9d21cc0323060ae35a48c6bcb5066f54e8daae41dc6cc46478030a092d95368d181465577e47ab5f4fb63fa540cc2243cef3725b5e3f343d19d310c461107abbae4f50c04cec8ed40abf87fc5b645653501e15f9948f1406411c231174988bb3ded6965d11068f4007468fa4c15300b79712c725e0b411c9aff00b67275b31598b00f13612d6df9f7d6a64dea3e1c368ee5034c18c4a895682152abcbec2e2e1c87a46ffea88c627c5884e96514079cdb12aceeea8076903c8a6f855fe0cf17db2068868a1e70d7e9f4c240850096d7bf2839972ac343c664f8155b00c38471ec977a5f344f3f9b79d4bc18e7a1974a3713a39a5532fcd972fbfbb5c9a21ae0cca8749484a874a96fe5505811d4a204f688654023460b65117f794a928f9bafee72f224f43eea59e1c09eba30b4c6d245dc477c41bf9cd95e50deaadedf31c86a8132bd599ddd48abb4e4773cdfdaf65037e58bdd79d0dbf4dd54566b0cb0ec76db4c2063ebc17a859d8ded4fd20cb5f1e36898298f1e81a29bd0d4920ea900a77ccdce0fe7ed1e527cff7b7d615899095f5a91df766a31f385980e5ca5f2f22881303653d8bf7c0a0bc72d394bcf98374a5d7427066a880624e9175af7141c8020c10f375cd318ee997779d06f9baa7b67ece6fcf0ba87fe581c62922c48f25ef66a2a13aeba86248c74c6c6f787313c5088478667d2c4562efffdfee3a2982bf0fa8186e0e4ee7089ece08f326b7c0f5421622e68c40156cfb1b0832ba29a59aa19479f45a39aefe90d75c9e4551ed715f37d5fd982ae116ba81bedd67973bd53917e9cca9aa8c09e38cc2632ea2a93e36f7a18696c950deabfe79818035e7227c076c24c3f6db1f0b404809250068b3a690560ac9e1ec52b60282c3e6f69bef3303c43cb3c2c774c5ec76cb802ed8b3bb4480aca7cfe2cbbdaeb92ba979039978c20e249a98091d95308e4dd31df11ba5355a3339c8e920b011579ccaa48a0628bf9914788c2c975224f81cce285857be4c9442bb525646d32ef7647edd1038af2701b0d2e39b818ce5df289e8e431ae374248eb7fa385341a05bab45e190970ef2ecc2c1cfe24681f3fef5d4d8aa9feea6f463cb532bc89d1288a0c72a978f62a862bc51d59d7df4d8e29560837f357740db0a9f2c6383bda7504ac14866874d2c06f06c0a7152ab6b303c0193ea27c56b8fb9cfc46694fa1c35ee663bacc45f20ce715a6208eaced9427cd42847cb1faacbc233ed66e086a80a6cbae1b9a3bc582d62999939f1408672607b7fe6d134fa051f9737e05449df7cbdd5877f2ba702a7bad4efd90766c3b6969d9d4427e7d14aff5c74ef9a488f43e0d10d2edce59b62dc96e251a1c07696c62a78fd2cb1eaf2ddd5a344c69a0f545612c6a8600de087fb4244db2701711e72acbd7a280ee4496cb6107782f91aad49db22d451e3b5a1eefb208a7fc954ba435b84f19e83c937165e386f2a460d9a0db9faa7889abac5b34fddfe226c085d2dd0e8f8634bfd785d8672bf2b829455fa396a406122332c0ae5ff061b23af7cbc19314fe7a2728d8a5587633ddf1b47405ffa74d9849ee1fec8a3f31ae44fcafc286bc7ac82793c3580785582fb5620e4a2eee9c34af722c4b4410fa07dd1cc3ce7871f037acf851b9d3e28c55e7258f998d88530a68e35b8c7d67eec08aba41835c526f22c35b15d05540877c7dee8f71aa9e8f96085dcc76c68ade7d9a0fd189d794c772f27e7c2bac65b9350806cadd4a7cb8940ef63ed319b51d8d3cbe8646a74da15ecc85a90ee8b92b51051ad7526ae13854b56a9544f109f184cb6139a997436018d69699461f473b73e9800040f8acc51986e4d60a0c910bdd400d14e6ef97c2b02b65f70d526f81710f5991f0c809fe239f1413207c9c0bd57e0e6f7599904b8e4f4b070d06517a83bdc316aa6db863ce815b47d4cf1045b55a8a25df09aa70483bfa595ab0af5f20e46a2eb7f45f3af608d69c3475387f0964e9c32bccc44187e82045674cde4b3dc0ca390838bba549c9b2a5a00381806117ecb5eec6d396c4664fdaae44a8e10071c4dd7c45ec6aa5f8d864a43f0def717105293d7648acfe75bf68f8313281d3fb315cd50242f8c109229a44fe19f05e04c89a12ea1e2d3bb166407aca5e5ed99178f1eb3b66761653f5397b72f7ea96ed80255410a469b36e29e854e9b653088d30cce147d4b41ca9a886668ab839bffc5661f5c120313b1641abe97f336f907e97156b70e22ffdad0d3c70a1293636ab2ba32bfbc80009d6a16636bede05631ce9dad40a4d2e66a35e3fce235cb46d01326eaacf2a245c311632070653341fcae0195fe4ce55f4f13b18dada4c53d6459707cc005b33de97c34ffb6609545f4bc05d02c3ce1a1174e1dec9a272993204d7e0e51c430abd9293ae81f74544913d4f94ea29a1ef95351417ae0b20d4cb3d4bdc224aeee6559ac0a2f5caa618ca1d0948cf610b0a9181a8199872dd7be6cac7f32c79b47cbd37a56b7e94ae158d746d875236b61fa9deadf81d9833d1ffbb5330e2366a6953eb54ec13654a940b5f3e484e230ac4e341a5905dd9dbcbe37f6dceaf85ad0f4788c12811c5a9d8c7bf949ee698b4b0b88040f580d9f5e9d663982821f6509509fafd57052a5416edbdc0d5898e2311625665d849238b09d3b741c6a8cac9b41d6bc54c40d57d0b287b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h23f32b96fa54362b60b3fb68562339afd0c1d31ca2416923b8875989a13446f215a800fa62c0d57df4c770a8d782adb6412958da34da12faf6366c8adb9ac9529d5c3be97483c5576a505462ce7da6c7db665777da1e1d40e31e7788f37281114ec1fb72bfb19ca8fcb8f92788a4351965c1e672636193f3907dea560733dd3aeac891cb68ea1e77c80741d5e01b2f24a9950f8f36b9b47364ed4deb2ff046e15ecedfe7008b03851aaac0c34f16c00e680e85b217f29fb86b2210450ae62d642958d7a4026dbd50603b53455263623752033e1819a584964c884aa292261d37eb4bcb9d4f2b3956ae9f7508d9a961586eb4e3a8df21b8f339ac1adf438872ebec90e9f6fc2945a72db215d99ddaa312a7fcf2dcc8e87da1e2e8b819ca784a4f107a19125a450d17956c95fdd230275184257d25139f5fcca155fe62942fea74087245bf499f1bdf9bcc8fe23c39fb08b6b4c3cbd724d535d2c3b31bf1955c36e41ff4802a25d1dcc5c38278f707374a5d8b9a3f40cb964cd9ce9ed0527e82377d92a3bc49209c6e3c2f9dfb7e2861efd398d662789587160a8021dc7ed4c2f772430485a6a031f13f26e037205c8947abf204f31b826ddf0b68d7a1d380a7ec27b3637f7ae28af412cb2e99da7c00891a3ebf0db0e091b0cb6b5acf07538a13af008ea87bbc80bb76545d03835d389ded1adb7e22116808d972f1329df3d73a2a21819264dedb5df6887c7f309479af6c77ad1d1806a3cc3fcd6b1968c17b5a52f9c02c2e51d525aa7b26be4f1e7a38468e4e4df21e961d6bb58058ebfdd891e2197887874e14dec8afd5e7d26cacc72dee7d7c247eff1868ace99ae94e2647eba96be36bca3d2b83b0e09214ca57d8500c73c7a9055a9299d816a1a30aed8776378012a5882deb2c22dd474e7eefbd8e5f397a3235982ddb9744b3939bebecb72ec0b679d87c5c8773eec5e6fefa027856d2a34c63ff1e9179358eefe306108cd0549c362551651d28be52d75493abb4642408c0f14f2ae49c9d923609b52ab52a16f575158d158313155e4cbe411d6abb048e474a462058083ac66f9ca1175e5cfae6b7923638a7273b7cf5362f808adb729b07adc98bc86f81a159a56a3b61aebee134a12d6040b176a4ba4cf1d5eab8abf8fb83744c6f57dc3737e0a75cd2556629f2d7cf7e27e8c2ec8d190b120ba56897cc34b2eee82c2cfefb3c937be8a1d376c761fedcf25fb74e867172180774ef9cfafcf96360f802bbb5b643b52db7dd4eac4a3ff5804c62a145755d1f757053493a7fd99258a1a62a1785623d6427b54a8c48c0fb10374f31a339cc563f935bdc2f52155279bcd52db68af901a2993925a66ef489016b382bab7cee0f7329db5b3f83c2ccaedafa5cfbcfee39fa0c8cd15cdba49147d4b4a9bdaf0c57e4a5a06b8032834f0daba7aa65ecb0c9a98c9d571857f9dc3de69b70477f3286dfff595ddafeddaf244ddbfb6f7be79d1ecfc56840a665f434dc609422a84ccf9df6c55c5e74a2acf7152258b41d513465ff61d7a346329760ca90ccc7314e20056d1ee7068250a86863c4accee4f5a47ab32835d90217de916b647b66c5756e3b88161c57361d2e24478574af1991ced709d4ecaffb86ebb3fe1f54135d0b47f951fe43d5f62e5c1ce8cd20354ad35af2eea5215cedb51df615606f2a29890d34e9287e5d74fa863bc0343bed95a7a48d315bc0ca028534c303c4f2a617c4f00eb791505324a7198f253842e768bd7d747f957d018663793eb2827d21dfda5ce796698c1d44db25182a3c022238b071a9b4a9732c2e1b867654b2cfa6ed60e96d945639eb08b48a53598b2cfd0df622db587032286158ec620f5351ea3f0c9c25b3f41c56455504af609353a06f454a23b1f8ca6e17287777ce1ee6cd80b442000fd00882c2b2c480dc7c93728187372aa7b914fdc0a4b0eeaca02d4aa4bb2cf836ea032f5a1d9d53d2ace6d4fd78953693e4f8195e8c2c1582b647bf4c20ab5b8738061e93c3b66cfb58dbbe01c0ff7d663ab1c99588aa6450f7ee90befaf798e51d27eac07f088124226f4c6c6ca6107e2dcdea85d88496a89d49787715c1f553a5996ee0d9315194c2feebc24780142e3e94e0243dc043ba893397dd8cf0d744169d53a4219a09b837442c57b0159271c16f87cbd8b53ab2784b1467862e5cdfd481b68db229c34186898cf83aadd32787542c5ea4fa36e0604b3e45b286ff5749947b713640adc271db4f64f28e548a2463837f2000f30ceba9947b09adb1b9667c22aa023dcf1f3f313420dbd6b76a39fe321be9e6cc261871fce039243f2c8b53de11ee85ada5c68a54f318f35bbe00a4aa5a88886a439f8048619fed6d50a5622ac86d1432c19fe681a8bb48c4cffe7ebd85952ad57f029ecdd427af35f5cc3ad2e5180804e4254eb23847260d933a105830511089677a41ce26ef505e3b88e8b98c5ede5323ce95c0b174984d030e88b6975f2c57f329b9737c83365a087d7cfe63725a50b35a0602ea4c449fe75567a85db35076b9bf9a1939929dd12f5a70aa23972b404165389acaf09ccb7af6da4c8d4adc71e3432552f99103cdbec1e48aa235fd95f7c732d226f8ed248baf1961b6e60d47206a1cf510d478ba4838f47041114a10e5a3f6965932dec3983c73576b49b371b9d42797a6076ddfcbd8e3c6a8ac1f40044dd725006e78ca427013bd31fe90c804c9a944b5fca6268b64c5bae2536d43ae782f32e4cfff21b610aa8bcd50865f29b8669974fd7427d9b9c10608911ce896227b353095a2ae108edf2e24f5511b93a379fbc0d0ba6d37bae8e7d70d595848b323dfee9fa806d7505188eccb847ac0f0752626bf7a694c56bcb20d2dc03ab6a1e7688c966877f44e1bb40292c92dcb5f6ec46ad88dd19d68b649c762c630e744402ffa8e82fa07ea67430fb6ed6de068d781094cf4b36d21ff36a694603a14d9c15d4bcc5a5755823e6b87600f1e54450571e5dba3c86ab47551601aa000714898052e24db965c791e7484aa1193d2dc2dc04617ba36b1800e3639b496051d4780b7395ababa80434ede22b7250e2d31525cb4bb744e650fcee3573a375eb3a46ef9482875c5fc0a4be8d2c13c1f0427b9b3da27760df92dd6ee31495a1eac7367d9c54b2a519a1a99153a8d13f8318739c8cc50044447445cd262aafb442959e433b8d10c18802dd73be744f57bbac422b83603dd1b45fb06c3fc499d3fd3f2dc4fda9d19f02f01b5d3db314cbd75f553cf21be39930a4f087baa7d71eecdb1de4df2c719637b00e4ce565f369c3f16825c437e554ae0d3ea135cd9ac262d5d9b1ac60a8e72e0944e43e4730a43f267088fcdfd05d5fd68d351a42509c715eba69232f23c14090367b4efe3ae1d638d855bdf22c1323dd869d9903487092fc0be5435c43195d6db2af7e359fcaff952610ebabda5d220c10f3b6be645b1fa49e5b4230502f1d39f2f48361ac9a5f5c4b31aef972e5de50ed32dc05a9d5a952d9e4724e7181935c308c970934fe9c1a33a4ac9e3d366b9324e361be40448f05abbe45ff3078f776137eb536478483ca42731c18797e2fb8cb244c2fb099627eb8259a8af24f202e1cde1a9e5dea74812b672731ed5dcb5150724547bd65b8c3640a53427a297ad10f450c9f7347fc8eb80f54e20336d879b4c6a34f98dff34d533702f2cca4e33ce415af3e734e7f778699f51bd076b298dd503cda8fa5966eda438eec4cb74895cafb78093507c01d5acd21571812990442e87b1286933488206d6fd6b836754cda939e0f9fe39efc54d986bfe91d1ac5d35b66ac7a616d38e9963eed0c8d1d35122cafdb534a0e82e0666717795d6e478939da8163b17ae042eed2aa0ddffcff0061ecc9c9b2dd98e9962b6b9fbaac90731d3ba70e41e9795c0609a4d238699fdb06ef8584456353633f9add63038ae6ae452abb73ef613e18c16e982167a668a008d505757e491efbf035894d5287f22b120ca91475c694e1e75988abf3e6b21e29ad1e3de401f119307f7ab2b55aa7faa7e4826dd1dc1e587608579b4669086c2f506bc317afaa5125c7d42c65faa985716590d95c044ee22317931416d8f78319c6d92cda78601571934daf1ad5ce7f76507dd53be5196a6797497adbb0c654dd41afdabf28538573c9eda0d5ffdd986fcf78997246ee899c3672391000aceb626d4fd8e2c9470071b4eac65edf29b4e6adc119dd3d530a52c2a02ddf3ac8f63f8ed7ea564649ec7f79517080001a14a30c272e8fc77b03da68077b54a93f2faee7a30ae982fcb2bdcc1c785448d5fb35e1076254166ac431400cb3b8fa8db79a93aa1c4a036f602656d9fa6aca9281aa979be2fdbd617f5c970abd27f6f6463569176be5237781e07141bdfc04a5941f3273fe9c8a4947e3a1ff845b62518f714ded7bdda173a6009107eb8083b96e6d1bed78b63ac470aa888e0775163b41c78e1d0322d2b2be7c89008e6ef15424b59c2bf6ef91a0ad04d6f5d7ed072e361c6eb5d25fd4c815019e49175e104dca4a0cefa18835fd7772c6253df6fdd99743dbfcdd8d73478fdcf1e7f983574b7ae2158ac70789a81e66b1a5b4fd6ff94ea4568687ca161306ef0ce423eccabf763e5445b323491ea9060624f2ae54770cee46414eaa9a16d8be63f36f2bc0c10320291fbd90ad43c5f5d33ea077330ec962577550bec6e351af5e5c97f50a5877fbef9fc55ece80acbabfb9783704eccf4ff044b655239e640a6c3574f5aa65dbf7ffeb9686df009b7874c543309a62fd105dc0d46b9a155af8a4cca779fc688e32812c36c548b06b28c928ad81cfe477a4cf242ee4aad2f97403778b5aaf8015681d50ba32414c779bb4a87bf92faa14511bec5391f7b3972f23dc4bcd95cef365d526c41273e3b48a8f0ba83d3d15c0a321414570fdb77b09371a22874c11e31f3bbad444879cfb8c65bdc7a8af7ade14e927b8e24c9e41bb5b4f5b64d63a777f74a067af38d932e7174ddb9825222d21da62700efb6381a6822a496f721140fd9d3357f8643384d4a39ddcb2ae67ded14aa4c1c8b98adcea74a4e1f47b6f8351fb4e27a2283e28297822ca6aa2801e9e1ded8b331279a63b8cd36d89fa373f1f7e6f2a101d1cc5c0bfd499e08fd2136f76ea362674b9c13ed6b391e7925c24616faed573cf37772d2a7f6f170d023a2e94672049e1bae92477da5472922ce28e7b97bb7920749a268285534bd2e17fddaa9093ee239026c64db9e6d64fe7d1ff10e3da7fc4ebdef476c64db24156ef00afe222d11ddc52eccb6e41712f7fd89b816195c589e43780da69ee78adce182e53fdabe882a24395036597a616669333530362929ff41cc5d00ed887d58bf6f02bb1134630fa56e3763a60f8de4d52c8771f1e2a4b9e1e68b2b97e85f1ae13952b83f51deec03b1665108d40b2772cf2799efa5520f2e267afbcbe523ec575492666242ff26bf93ddff80ae17fd4087d53be69fa3f2c4a7db8cd6b912ae955ba4fa53554270e8a5f4894aa76d3ee80c673c0543972b6a2e4335c38437e18050d2b852acaa2bf71a7ff2d03f1f5bd74aaf60b9f355a0ccfa8653ef5dea094c11878b31e46f5b8329815a452dbedb4eeffc4f661c56bbd3f4b89d7be7745a77da014b0c2e5071526a97d3b11480e99ee3c4e8b9660064fdb5ce8a7cd34e35a99f344c2af026b40fe699622a331c182f250f17677e8754737cb94b01d03126c055293a68f34bb936b63900fc73e471bb2f97496aa21c410d3997878520;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf8bbc8822d581ad1ecc78f2c5e8ba5ccce5d3ee53ede9c59d887e3af211c7c08a8d4198b0d3f1280038ccb20e015b8ab167f806a4d1e7b0c5455a1d6af367d678bc3b7d04f810e40c44950903c4ebe891539d1b94be66687f0c0ac860cd29588068fb1987f1dd1e0996e8d0d954a17a4cec8ac161163573e21b1fa2099205178710a6ca6e68162c07348be933cbf4e6bfddb675486bea6bc6105407996770341edf49a3cca2076b3f60de7228f4221baf6da90bb7b114888754416c7cd9be6df4b8ccdd6d11e70cadc899001eaf7cd104b690aa821ba5f2eebb19e79ab120c650afb7516b4486d0fadd15c4cf64a1fca9b971f10f4fc7e713dda2f4a030194266798f8e632bc9561506ed1549774c962529cb79c541f5e0445954e051da23563d1879216ad679d6e415f0e8c593fc02980264139e04c982f62d2f5ef1c730a74863a68ac9add7f65a3719f6bafb61ea7459d8d76792be3434e1416abc60547a2ca17c275b0a80e0159a6149097960b030a571a842ff50eb3d41a9d23a523b8931c3e9da5aacf4026dd5e7396a48b723be0a8e2cb2ce3e92e8cad9d61982d1db9ada8e384aeaa45517c2f3fe640038e63e922367537af01081381af2e9e52fe267bdf57cb791aacc803ad0659fc262b6d48050543a02e6e380b8659159241a11988da29919cccc7f8698d4cb6819b3889950f7ea55354541273686cfc0061198f89ea40b99a833b2d18fdf19e0f7c4c839276232b6b48df4c383c316238f9cf54a061cb3a237c1a9987a9813f567ae01214aa899b7588e8c6bd71b6e7cce169b236ff8ca637e618a46e4881874ff67b645c86e4b230c8d7b9d63936c57f048f97b0da908dac413590964cfced36e0cf5c9aca958f7b32163db8a2081ffe5366c70fc66247b3378caaae6cb0212835a0c9e663044bb0080294780a86e99111affc9f5c2b0593807fa67a3bfc1dbddcc64674f3c668f2c889862d1658d97cf4981708d0f351f51d2e45d60cbc3a7092020463005f0c135a27a64e0a3657019a82185675d2b6f2e137b80580e5f02768a9a61dbca230e5d44ff91487a1d8225ad4bd1288c87ab5b2e929a9a9f513034784319642f32e38a433f1f94a9283dd7f617f1fce5ce8c90075be21506b0a6f3759fc68bdf551c5515e7994df2cf3dc3201b23195e010ea0750cafa32b616bd9a614b53253596a3cb0e10ca4854d1a60d91da109f5ca3b282ab268e9f32bf5112f41d03de668fc49eec9f192bb2607b6445bfc869ada0a6ccb6a4894fadbbea93455d961552a91d4718fea76c77fb8553e2121d56d6bcfa3dd82821b03e1456173136b156203593ad467275355f3ccd1e20aeed3cb128cc651cb1c018026d5f532aaa6de9e89fa2a9fd0d0d28685a14dbe137a9f3a4cfd9e1961e37c56a11bbca1fd8a082daf6aa63c115372b5992d39e157f60d9ac96ed68b22db1f2d3fc88870406029d48fe906615669cf978b1fafeb17c992b158d443dd43dd7d0689d91c712ef73976d66f3f9e0b894c7553afd12dd16aa5254c06386722161b8017f43a5d5291ec1c1f1750c54fc87fbd72eeccd719a9762684d7b5490e16c2545db853be11a02dadbbb2196601673b282619729ae2ebde7e8e4a31f8846827e98b653a945aeb01646e4d3e35978e2a954719d93f29aeeaff945555c4a6fcf5302ad7b84e2128109cb772de5de38b4a0b44283e9e4aab3ed4bf79a92eb41715cef0d09ed163180fbbf2a26564ecec64594722a69cdf0560ffb8d793e7180d7bd5cec9da063fd22c6a9bd713018545ef3b49245f1e4caae16991f7b61502019eacbc5bf4080df67b6c89f060eddfecb8ee901226895248aa1ba35f8a59b9c86d6c4e8933eda78092581c38faa77caee54aae07cbbdeefd81f390c0675766a324d029af6d1a76da201e322a8d4ba98c6e6a47c7200d51e32ead9ec0eb4fc2fcee01758c2d5de892c41d75f41f0269af09824865df88b4426f0b3fd2dd5ed3066401820bbd9316965ad45ce8cd061cbce91d0a7104af313a1c789450084f88043a08516c14c626b5130004655ddb235d4f6a92650389ac9f30bfd48c0845b7b39f05bdc6987a7d05c27bed509137b77b80944b2a57e12828d161507d0c54995ff86dbcf51aa05c144db84e35b52a810d36188a4c8feff9ad64a2b6d959cb40ae7cd45f23ae62132700efeb30a2bbc8d762856c71a3316ede7cc4030944b9b536c207b798e46e5373d01fb263129c6082fb532d632f0362588e3d25cf6d78cd6af7ef8702840c1698a5146beac7de700bdf348171a4ce1fc014051674f1310cbc1d85ea011cbbbd7e3c2d041f694accd18782c8e1f3df067ee0c5776b7d583b5be3c68b922ad63e84b642ddb8717624371de9f9623c3fe4784d1332b55391764af46149d4cfb596e34677592d3aaec00e06ef87580b44db480ab8f5706f608fd0851ad27dbf5a0e257dc786b1ec317d11ea43548bb9114d21fb7bf284e92cd922b26ebce491c8896271fa08253e0e0454492e1de84de86efef9c778c3f0b4ad53df0df9c5ca09a6aab3e68d337d52f1835f3492767358ecba4e390da4cfa5b5524bcdba09fd9e6b479604d8fc873985baccc6c6e05aaa9ecd4ce6baa37e6b32e4aa2a12aa1ef5e527c589e5e69ae4f86f978e372a22cdd1f81bff4e51efaf264cf58872c99afd184c90991c0239178d5580a0e9658c9b82619f98d537ac542d36a057308c005c69d31c460bb6b7244114c1ec4be2c7423a94072d59c43bafe673d1ce9b7c1041370b5862be636182a168428788fb78a5c6348c8780ef672c3cdb5d10b671419480232d899b424a42438c9a8177a887bedf9ec36144b649bab450fb71d0e79fbb2e53e36a0aa3a78763471232beb80175a18a93c3a99f31f90190f143efa66575fbaf19d844c303d5dd6e37a146b2665298a8ced53125cee97863d1dcab41bfe1ad293b6e08de20b6de5b1ef034923dfcf468e541e854f0c2f6e3a981dfb6759ef90c4043c9b427ddb0b16d574c13a20cd812d57945fd89349049bcc0febe21eefcbc0900c77d480f1d58896f38c0e1cbc8a8f5a8f8bd0eaf8c40bd9c121c45adaa17284012eafe4b5fc2620663fedec04886be529c303922d739da36dc39ed4ad75968a1ef53bd2aabcdc96d2f4a69e2c0f436f424eca10e817a24cf2133273908b95124e831b056d82104890868258bd1a971260e6d6a29dc533a2dafb14fb41e86ccc210f99dd19710487b6ff4b41bfd6b30cd17ed2ad438b5bafb1197484fb0782c0f57a8cef4eafe8fb9c4ffbad5a2bf42cd76d4e222a2e949d8c821bef7568ea434523d3cc24e400af100d5bb7ce96937ea9bc79dc63814dd2eab2c478f3a9d28a59af0718968bd36972e477e9882eb23aff1d67e6b6b9793d5ad8420baabc1a51decc6a7d78934a144558cd268e06a5d76d574fbc462800ed661d5583e222e6fb2f0c92886ec67feeebd5696f633f2f323eb62e5640e964e25537a0b01b232a8025ef9536dc180a6928aa4066b0a0fa30d85b24848fd7f952cfdbbe4983fa0e25679437d8c225ee8a0c4d8eb9e726ccbf40e3043d09bb018fde5c8f3c7465e869d6c3c5afec3cd8b8be2dae1f21baaa2537033dc2a5a8137458dad841c6eff797817f0b72b37c4303aa781dbcf7df249a0145e284e21706b866738a9566dd0a030f0ce7fb171a3502cfb2678cf76534f4924f79f46112f9e12bfdb928831a4aa8c811759c4ee13019a97fe8ed4e040c06d07106890c7f685d7cc6f2ed1a1605fa49cf8cf6b3103db85dac0d7524255ab3db34ba84088a1484fedbf031a12859d711cc2a8d1d737cdc1c5065e98e03f9827b534244e586b7a26651e78dccc1ba1617b1b0f077d420f37930d34314d954fb586085b53b724e4c104823baa46473bd66358a3919acaf573ca303b156f7417dcbc9b67b20aa72268a108a1c6bd5acf0f6ce33eef7876869d4ff0ce6d16873ac3074f59457ae62cc73f20e364e7b8b3de4d2e253ef4517741b9d7a8b97e9691fbf097fa873a9f9748ede344c96cfd2a38b81575f816dec3180d7d2587edca6e65ee5425afafdf29546d2eced0d9659dd8b72df8e7b9c897df4810bc4b7c28cbb084d50f2b427d64f5a2dcc7b50e6358b812059967485e6b5ad5a046aa442a9ed9330869ef58a75113f0685e427d2f9fe9a27a9a47396fa18f6c61ab5d61a38d9942d96bf355b2a98c138de4003bab28c383d49bddd28129097eafbf9ff557ae7d77b1cd6541bc161b3e6b38bfe8cf9933e2333794bc72751536ed6754da94ac0562881d95f4b86aae10522d11d4b353c4f13e4fcdeeee6280dde402fa248ea67421ac432b6d22ac5c4715618ac885bf2e7fc1642934ebb6cbeaa4ec559919df5e056fd164a31363a68be76a71b0be1ba1ef3e7e06edeb40a35278e2f6563ae579e286d266933b36085d9377187ab5bab0ad2120f8045f79fa3f4a675cdf4f2c0216298c4269334cda7a62f0ce24ad702efe11f9ada0b9fd08ffe774c716ae2a0fe7916f42cf1e48b63a7d58c3436ff717b41e0efcc1de6bd48ff5ce50f3689b7d40f3a401d60b28ab2699d679225cb3cff3d48783eed6841b5abeca16f9f244f3c9d4ce7514684f6ae3fa8498013da0c2a0dfe4d19e4630ea29a52b4fdba232a87a11185c309569aa90b7ad1787a21f5d8ddeda5d9721d5b3d4c49be8c3adb206ae7552d5fbd36443c8829b4d53ea1c8d4ae7fe2fd80a4afa205d07002a5ab9c34e095fcaca730356d58460132c0edd74bd31c5a3f7f663b8c037a29a069e42f089cb36694c0c11586124b6ff80e3df18ae600f6e72adc125d9619676f9d99385f3c2daaeb86b72f6385ae8f80ee13451fc2736624074297bbf22f7adad023a8d6b814ed2b2444d2e083521ee965a057e05cf258a8902d88d194d823ffa343c0f7381e8b1a928a59a8f90c371b1b87a323bbb8d2044034a60c0b6553c63f97a1d792d7adbe7179fa04d0de2e9fd09fc3b58f8402221fc291325046eba14562b7aec77d9bf087e9247ffe0428030e4e4905e7c571776972035583e7e60f59fb3c60d9bceb24a8597b07fe6a81c8ff38ccbac14746ab367f599e51ddfa9c71e936eb6ba1c21c805130ebb1a0ab7a0aa7139a9d575fc1620e6656bd7623acec50edec7c214048a35ca5fed862f47fd8a4843b735cb9ade2b767e7d0fe35c10b193e0bec519ac6db2747ef530f7fb9c4a8644829d2185f1b839c646fbe90242350b36f53ba8bf6ac950ad53ea82e0b31e3c35952ae7fdd98eb3d94aa74402d9485f77d56ceaaf9d41c9276ce2770b4de32c2fe295ba17adace13ddd48ce35bf0c558643939e5709fd2cd0dc398e69928bd9651f8442a6f72ae53143f55918b4c24aeb57d3e3f7fb68af515e377d650a2165e397c23ca7d3e466ee619686247331dca0f12794dfd5582eaf5a1701ff9c948b0d1a078b0cdfd3f8c39783784cd732d0c59add468e0d67be64f3d940b6d02242744bf854e7e537525c1caf58905bfea733510fc7ac7d7718ce62d4ae083f3795556679600d2d9da4d48496534fc1053d90853a6e628f90bc89c4ffe9b56c56ab6efefdaa99cf16bc716e02dcdd79be32d8476571df99c4463ed876db46b7d9b33d38c789b65c686ec95ae3d736fa4fb518dad8b466f86123afae37163b4fe2f691c16b955c623be957ba3807fca6568e22d14153e88853e36fa5545c3f6d885afce91749bcf576be8c8a746032f0b6dc933efea3d28c7c8697936c654c32bb9d666dea1db1e6d98a0c117f90c8e5b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc354502056163fd3aed35712397e96f7ec8722341c2fbab7541513bae45ade6203eac69b7a3890f19ab6fef429f1be022b5b77b24caee1c4ef922bb420e08a82a343822262d0b39b635b51d32977bb23909dc19a9611a956739f4ccb22eb8fc0d04f9d20dfd1a4cc75898dbb6fb60e3dc4cd655ca9ec40614e921381b5f94b0f5b21f541fdb7e114b335bb8f646359c729b6fc4e02e11bb06908978b6240aa7f9f3ee0c3837af0baae8608aa66a792889ea5715b45ab4d53519488f522fa86f0c83558d10d2acfdec93d9139cb4d3bb2f8d876f871e852f6c680e0cbbe2a9b2e6622c93fb7bd8bdcf67b04b972e3a18ea617e02a79c138a53d0f62dc452eb9d76b0a44c5d7397cd388546e2cb7d9a0202565a5cb2d0bdda4f84342ca6d6aef68ffb96228aa5c99024ffc4492b21e6f88243ebd875a8a9354a9bbcb55d12ff9df79f627fd0191062d1dae16f59fc2d65acdb918349edb51f6726f6ca9dcb08808ce058937ed69b483da8ba4381fb3558635b4a386a94986a03616a4e40203e7b7c070e9f2147536b77c3f47c5574e9ce002146e63d6ca145d723d2d526396bd7d69c17c9ab35bc3d1a17573ef2565cb279677e601b4c5e6060da58e92ea90416991faad8b76798628e55c8b0f9c2643fbb76f0628e10dc9395becf78ba4104774551479620fbc07800d82581fdb19f0b2da56f07d40538c4f39332c5f356326290940829f6988915c9e811941c8aa2ce99a8c4136476e3b0f63965237e127285002790cc436139f4252919426a14df5cbe7579c8829681fd02db25b9e0a6a9b473291e86b6b8f7da60820a3a69d4e532f701d85292ff159c330ba103c6d91b1f481fd65e430a9388cb9ebd0b5a8b83200c80de1ae209e0746701ad883e1f0500a9322e603a93e98c78ccf674cb90ed8656d9e652b331391946c7d2ec2e691fe5e874d644655d15795ac843763e56ca7ddb4d48bbc4b943e99733d5ab9943b9a7e8c2ed1b20b171438ca54d2f190edaf17edcc1631ff9bf77136f19cb7ebad20747d45b2de2b1caf0666c53d9a65962dd4e30deb2185d2be6b3ea1515cfb1f7cb98cc96f7673dec6511559a9c8f3de26e87e09859dc40f4657757d01d59418a42e144b64bce18d1357daa8f31ee311af4c9d08a9bcfd2bfef7b080bf7923d39d09137ae17d1be847e254c50bde0f8f9b60218e7b5a6a8c9f9bcd9a4b210d85d66ee482f3c91b7a8253aab74d7f32ce012584c47842decf12b9699190ef37e7c30dae61bc43a380fb72de302a4926858af0d7df018ad441e914d849675dd4b40623da85e5328be707d63ca70132895ec292394d7b14ac0e64bbd6e962746891a278e4099d08916d7e9743fbd5ab7dc647de97e03b12659fc14515e4b3d18b97021b3ae5f7b5dea1d3743b5478a08cdef85a6c847c18d382a4036cfa0d0dd2428c1709226d0b298ccfd621ffbcb69215fac1cda0279215e0dc40c83ce86ae1ebf06e144f5459acf44b021b454c7b8151b10f6c6b7bb58addab2f53289f1fba89ba015f087326174a7c298f89f1292a143bf7cf42b1bd705981f5728b25e3318c7c4ef30e54f2ccfb5efa784c1f2fc12cc47548a3a3424289565d876b25f6f45997439ddb3c57c34298029479bb59fb907f2f5e99107b7e862df4b3c69b2be89f5d8c3d1fdb9cecd32498f44e56ce1509905993ae488d8156996c7c2aa29e9e655766ba85f17be9f246e324cd67cca464d3bf39783340263c8a0413dbbd72d8a198f12c813fb9eb0680df206ef773643f9d951c426d8b6ed6aa4a0fd2dda6fc4eb8379f2e88e3f0e39b5c944b7a243f0cceb8fa4dec812a1a747542398999231b3709b243ef359d32c1c9f62c3be15b8da5c217c6d797e3072a4d7d76c2fd3518e1704bf0adf0b736481f1d82ec0e9a1ce97b6b8fbb83c5151ef58cb20668c79238bb40861fce5bf815fdad5fc6d942e0ffdbe1286a783c0651ded17607b87be7fec5f407aea2c73517de4428bafd4988fe10a035f56b85169851d8b9398f5c57e35f5ee4ac49a9b98cc6f8e8786dd17f366c912240a59ab5a55ea05807d28009ee132a53f6c217e7dadda395ba746bbe3257851655b74080fb0f98a767e326cd95c8ec921c1b63dd8a40e324444a9025e1051ead1ea756e98045e60bf8c1c85b5a5a4aa8a34214ad67b7a10748ea15aa093e8c844316c88690d262876aed2340d6a4b5218aabd166e1253f56f252b027721635d81a2e8ea57b659cfa1195a66c93e8299125b7c634f12adccfe70c99f8e0f9973554595ddc7a226272ef74a1100c409d98cb99d46544ef22fd71d8b22572e2fbace3b88aee57bce689918d487dcb564e7e4570c32ed76a0968aff13533828295ef28956d132d994226bed47afb888e9c4a731902b0b5c1b1551660db0386f1d63f64ac8642f0fff9b74890341ea7094db53425f4c29c2cea83a4641f8175808f9c3d2925ecb1ddd985b7c5766a1ef3db7575b8c793dc23033a62eb4b0612cdbdd702700ab62aa31b25886ced8aa2176910bd800675d3fa975316c21493d5129ea86ab31b89960ea981fefbfa2a2d9f0c67e966718eef88e729ca9725d2599fbe17fa49c98ddc95942fa5a19feafe0d4a9ef5822db290accba6b6040dd66a4d3563d6049861f2f3a0844c1c3d5e2c20f47e6489047312dbec6e9be1617543d13fc1538352b120a2ba2ae7b9285f5b0fc0488ca21c24661cff30595eba90880f896e35d0d12af66a2bba47ed0b03dfe677514e5d40fae8805e669b235d05694dbee8713e0fd23564a680a1d3c69237033cdb1aa4826832231635f57a658f1c8d3ec308ce504d461d403b188a8a6fe664dfa8bb41904fe5aec2fb7789d03cabae510dfbf58b257294637283c051370dca7dfa35d3189b3f1c1d14ba2ecbfd019e4b6b4d501edd022c8eb130dede3717be21c5a6b13647bd2d17de4165ec240d683674305f8ad396faf468f411d4389120f6e4c64fc0e59869f4580819ac06b4c0253d9ac5b428187350168dbcb9f6958a119dfc0924806fe4f4c5ffd628c29942a9508490191c09ef787b765edd014b25dd7d0ffbbb7f9cd2aa3fd11ac43412d672b7b3802967cb801bb3dd04a23a3d42208e3acd78623720fc9bdb9a250858e20e7dd70cd78af36f59c404a44356dc639365d4a9714934860b99bf7e6edfaaf7b3920676ff3c2a4d3cc7c685f81d9685802262003cede92bbad895357a4ea2e6e5e8fd9c9e1cae56981b35ce4fd4e82fbcfc8527f1f3c2f047cca8fb47fd849c826efa07f9e1ec976f6c16ad312c541466710373d0610bc6010a4b2f6fce334beab8b4bb85d23c80777318fd72542c575ee96ad831d36145ee8c3a12659870778b126a1578ad83f43c0d58f8b09975a14394883e9221ee3ba47d730347b156bbc8fc8ccc29995cc8d4faacc9ed0dc2002704fad929b7dfd3271d0aaee56b9b79b61eb901e639ec49d202431e40000e97d254d6eab7910a144160c4c229b787b0bcaf057dc621963ab1e0064c22240cd2f718aa11bca0affee84aa9cf947f89bbc0be47f0d584e241d1a26ea579eb90a0b57080be7f12321514a6115aad8d99926e3db4d79ce22a00cc5bb45aeaa70792d2227d1178acfcf7b930f3e05d835e67aec21a8d06befbdd67c170ee89abffc599e82cea44ef48dda34a4c146677284d8744f2e200791bbf74e663dbaa677b91c81ac792c757b4b3aae1a5ccca5cfdf9064ed7176a3850712b4c584a600867ac442a580e64b23c192e5efafe067e37af8a1d692e40f052f9c5c5eae9ba5c33cba848cee0e06c54314f1b30950b5a1010012474b202ba3162faa5cd99e2031b81a8f4dd0e157b417cd66f5d2ee3b20599bea7c75219f426f4bef37a19fd7cc8465db329ffd1dca02eb15250cdf56912284ef4aec70252b4f929d35e2bf3bdf4d44e84bcd59921aa61a593cf5294315e637be5e1b2ffc7a4b9a83b87591080c3fea5d7efc807a5b4423ccbd67da95041c06c9fa4863768d210f707964ac80c66da603190098f4a84990f3c402db61a351880279e2fc67eac14f296ae354e9f501f16ea1dd949a2e71a97be25261f656f19693d94dbcbf0a7dee8578ff1f143dc47b08eb7e181ea88876c7cfe22a603bfc7a02718ed186c1cdbff005e957bb3786ce2de9f1b977c959d6c9d495804618fd2dee3db92c76c652e54368be2a35e0dcda9473cf805fbc92d237bf27d8aa1dc92a0f0cf4d725814170a85812c0d8f808b2e62ff28900c397b1a7446593f9e10cb21b269379cc2e6d72d738e526cc4ee621e8940757cd8e8d43d17b3fd6e90853ceb1b317e341aa3b9daa26830fa89554c4fa007869f37d0dc7353a62ae58381d935f2e7fd85fc7e26e35a64e3a83338221522f49dd824d0e8ca0c0a4a1a5d10554e856732ac309d2d0a852908282cefa7d2fbaa41e91c1c4c9dfe26b8b97635bf993103b8f197dca64a229f72bb6df05d7b3def2fae18281bb966b410d87af5ea40735fd043974cc6f242298f94211467504b5052cbd59997340a340b304d3f8cc77e110fe385801b583b4a6ce4f13e757eb51f1b495a988ff492fd8a71d94133df4954b30858c22ee7bcd4d798eb2b2e7fdc9a74a747ded65a973c21442ea2555c83e98defce682e1977e96727e8d2d7b2964b0a20e9191e59fd25143ebfd55c4599ad8c72c3daa8f4cbf15381962ff0f11932f9294cecd25b31e410b94ffde022cc3e9b6ff0d3ef81a207aeddd9c33d2c77d08c275a4e6e91159123f538dcd023a1c7740d845ab9bab85479dd6cd181c79b0771cc0ce34261e51efef465785bed41cfb596bfc0668bf97158531409a7f8e4dfec62b9b0f5d2ab7c67a4dca3c5ebdd724c580ae78c5dca5f10f9e9961e2e0d9822ce7aaae26f4593e64f231260e0838b4847d5b0aa6e14781f7701d8415fd82ebb1db31b897aa6601558f5b86c40229baef67d92c0267124b6ab8e3220d8cba8cfdef5d0fd07cde47d481b59be68b33ecf14957801b9000d1c9fa23be51f3522a8b304ee345aee0c6a7e2db888f7070fd5162a3cc0d71cadee7360d4ccc4e6cd3393fe07660edbe1496ceb670d4c191a851fa50e907a33092a16e6198ab4ff5b5abde50f29c56dae0c3985363a7227f5bfaa6121a74e3764e204db722403dcd554e5a2b5427979e1becc7696c1a353007fa3a327b6bf6ed0a9eaee26dc1397492a4dfdbf59dd71fcee8531f9dcc6baffb1a49ac2ae1b891e116fd800417acc320b5398216ba95a77682d720c9df0f2aaf671b3e2ec71159d2a88da65f35141847600d5213471e31fccdacce1ce0999cb518157407993e18f0811b36e0bce938925e1c36e2ff10b79f67ce54a045517776c26fea1f2c06416ecd717904e92bc5283e478b8c3efe38891ff83b1538a1e7c6c87bcd895a75c200ac1e10772a3bb95fc3555180ceefe7f2feac1a8e643b1100e6748ace80ab9bf162e4895b5740290d9a67c3a2189aa932f1f22df8a1ab4cfb1aa643a58e7b1d89785b0ec6d9e0dd51cec59b235690ebb58411cc0a76a96454060a9e0c7685dc759f2ae31282349033ae701ce95494e0ef63b360d12185dea35aac6deda9c5f18d6cf01da4eae3f7565317a5843d9900be28aba894452ff6044d781da124c001fdddd2a9f1b712604c1fed6c26e1374c6aa0608690fed3c95008b4711b9b48b397b6fbf14eb770debf738f26f76f88960a5696c479a7df816e7fe342cf5a31ed79a184268ed450ea685033e0524f7831da57a2abb8c110662e53afaf8d67d72e6819cf8b1c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h26167b6564dbb4072d64484b124bfc31f97b048ee8dd3a343ccefcd86ca0e1f737a11fc0c229089e050218f80b64f48ae807f488686217e4d95a7740ef285e00fba597f87eb9580a45cd4d6523ca5587bf6c239bc600dae153f2421a24378b3fdae2e7589f0a2e2d2148e7d7ba4050a6d4c86083ad321eaef4334e80989f9d71b1d84c98d52d128a7c5176201ed4360e30e961cdb18068ae1f2111ad91aa991f276ecd0150248a3864fe9693d0ffa67bdb8dcf4af6099be79304c7905710132d01f57d583ce3e82c3180d207b851e299e2179d9ae36c389db04e86a216fe2d212e9deab992276576e3a3e8af2248260958e2f5132316c72eb84d96d5d2daba032ef81d455202ba86ad844b95ab58af46719f076797ce1a59b9cb38d3a159a1497bade76a3f3b587c279365690a56fd2baf47209ac48ef3f2fc309fee33343c6372b13c78d8cb8cd34ebc0d7f4a97a10999fe7dce832a35e11eeed930288ced83aa5f3a454cca6328d846e3d8b6c81401dc58e6e025800cf21b9fa31813a1df81e7a11aa9229dd250216f848013b882c9c570ecdee88689ae7d4c2bf90fbd165d83e940a128d82db94f6c24e4557cfa15fb96167cceb01eb6ab272b585b2dbcf6789a42ba75d33f97dc93ffc3405564e52a7283f33070560b2301c8e06fe4067fede85f9a9aafe73086174d4dd095d7dd0c789fc9371fcb0d5c29cf2ad36f6e69becc9a419aab418cbff4dcc36aad1ce1a474b0d8f51355fe9e7cf68d59f7ee586c3995ad81810891f7f389f031a2b22af70022a394dbdf74acde6a8689246956270ab6f437c87b01551a3641634ecc9107a21f8ef2de690719441891d7fd31ee0669ccd88df945b24435575331c2c93c45fe24da7a607d12022d9457eae707f678f9b9b8fb75980a7a3330b15b0c8e3b16c1ebbc87dae738192e2525002cd34205522ecb141b044b684025c86d0ca796585a50d8afbb40d587de4e86a0d120b59f9155dd48ae9d9c53a8028ef80353996d4b59c0d2782eb97d77e6f16443f2dda7f1838d08958e60fc1a9444b5ff76c10c25732596ee780db81bb328afe3121fe020104b732ab81ecfffcc327ab8fbebea7dad23c036106e19b5c719b7edbc2305d47bf9206e92416b25a4cf6f20ca5b4853425f6852aac4165958201c2723d8344947b754416fd59fe2ee4009712844670d63fb4a0316f9c09ef19748ab236d16f236b1dac854344cf00f986f1c3f5194ef223f6eeeeb1353fd314947c6fc06db2065e4422f5d9d226ef31709f1e64e16d81fe15a4162b8c306c6a51e6c167450679150358028cb01354d0a6e30afc3a6c65be3fffc0d8ed22649fed63d6cac107df54d7231261c1332bd8d93089f64d785ed429c69cd694936f95560c6622bd487df36bab3c8a1962a59ed99fd97103ba4fdec961086f7fb7e4fbcc0f48b429627050bfcae7f84883326bd96c0164332c306ae33a01c17c395045c6dab6c2a072416addac74aa62084373a9bfccce495d7d767f8f6826249513c3a9882c6e5de213dbcd1d5aa5f39ac2a93e4886783db7806430b559588d70a756bbd0c1a0c2063a998eec34ec847f8eea560ce661a4eb77ba392cf895fb57e66101903feedd8906db96fcb30dc3d0fe89c15276c1ce3a24e78486cfcd651308651d4aa137345a65086b65711e0f43670c9bf4b0f1db0b1cef19d376ca5d726c9eba892fe828e6fbadfaf42376e05878f9b1f1a927fcf25c9ad276b01fdd91c7fbc40e2ad655999ce0cccb22bc432d59dc55b34789319e3492d9279aa83c7b88704ae60e04b6357c32953f1827e7d4e6cac9314ea85be996bb30476c23c01bcd1c1c36f8098c395be9319469f55b5fdd08b8b0c540ccb64fbdd5946b3364f0adb34c3e876a963b86cd4cdc81ed25c09bb5de6b39b620f688270ca30448038cdb661dc5ff8fba307b202e32dd2e62fc9ede28588bac97d4c0858b932021de6abe6b597d70726887dee3796c0bda5ad51f244d325a635eb994fd9ce0fdb2540dbd8713985ba4fa9b535772e58010f9f1fe084e1494c2dddf3d3749431ac84ac46f45743aa7ee92a903e95131fda2ab96751642721abd4b45d10050c30c67fd7b9bfcd567096932361728772ed663c77473e883cf6fcb76f1067048b11bb97f3039b1542a18b655bb343cca25c43998dc66583f2695f59304441f37bc1176b772bdb94dff01e8c8a127e218a6d4e102e5c50fc8365a012df332f3abc224bf28acb2ad94b34baca44c3352252b255a04ce80efbe546b3c5539ebb34bb847c53149a21e36a6778f267450f80346f1c13fb9c663b601339fa61f30d4ee6960c262ef93f19512985011b62b2095f972ca3fb2c1ed6980a0f36ae22e2a5be61ffed1958cd4f803889a9f0f51387561245dbbddbc4ddd79d64466f3fcb6cc0dc55479f7ba18bba4737992fd19a61bf47a2ff58e26c5dd0b5ca993ea1c681332b78c2d4fa44f2e43055822062c09871622949d671bba5273304c09d78a0092b5fbee06cb806ebae273340969a3000a1ebf5ad52953c1de20eacbd5a2216b85b729a5c3e598ac44854bb3219aabad921550d0640158bbf4b0b85dafc8e2f4f616105a8c2dd0d322068a1d184f95ba4847e70d1d6e4bc383914785706c5694e12d05f7828d7725d5b38eae764d6e8c1b6d17c4a33207d38a859aee1309e9f15038bd08e07591f47a715981d8347bbb6a0e8c058d0bf89d6955bc9f04700ce194d2781581b5204c7531122acccffbfd5c6ce785cd7c63ea2b5b22a9fe328b89d5cbb1eda22bd4aadd01e146b1b681dd044446fcc4345a946621116ac3fe94b76fa8ba75774177f601be504e6f42ff261623b1ebe6f3cf5b5db927e3fd0a9593d98b2ae97ce307341cedf9253c2a40ebaf96d0ab5133ee66dba973c35fad7fbfc261434a0e372d46ad81870079755960eb8bf8a92e1af770fd1ae3c8f4cc4d5308e3a889dbada2c8b0e75a71cceae415fd2e6794f00b058483a2038a1b0825da804c027636ee89f6c0804b6d2cb2b61a352480e23cbc0981a90a631d1d63b3a9136d09395443bc4b2a041fdc38f8a3466ebcd775dc0dc5ae3c748b45302c369fd69b983ed9eee4c16c2e045b3235babd695c4eff05a3e2c33a3179b70428e9cddba9ac0985a601846a18f3baebdaa5ea96c99b4cf3ddaca011b498ebee7889581be2445d65eaf4e47c83a90a0a6477c154b2558fa85a90d66e7984d3b6d22a15f5994e3293f305790277d39c442e275794ab5219dbbd7f9c1c2eff515f46d43b99dcc9bc9cb0368a9fd66a203ce2009cce2b2b4bb8e98940734ffc8b177de0829f6333a0e6154e91cb2d32b7386b9ef68149a220b8b9f5d7e55506dabba70d58d17c0d656fd1565d03a9cd97acf5c59687fe3eaed2341f7e0704aecc7027270954072460cc3d82f5c64cc22ab03702c39ccb4eaff183d5d3a525b8095dc6b33f3ab6510767a0bd50039a625106586bda545a48aee624547e7cfe6893d5c20daaf984ca9913d1678dba199d743fc31334170872bc70aab3fb606d0ecca727f5c8a8e3eac1c84b4b58f5195bbabe1cceeff5da76ae834325857272f8c9f82b210e382a45524cfaf817c6d3f6eb381ef9df4edbdb6240351850eac7e9dab0bfb1101489a7b62b79f00cc82d0eaaa308470e6030108bee2a8f7814b5305c94b3e588e4598d4a19aaf3a65964b793a6e661ba68b1c9ad0b073478aa7062faf9056294188ee84dfedb436a2fd274059c5404a1629e21e9ea29019623712579d1cb58e0e53ff761abb2f98faa72d8dd0fe08fa02d743feb7dbe30e310fd01047e8cad82cacc3dd233699e32c60619576b7776c2cd98585244a18092e5d80a26cc21b6aebf901f190fd33e48b053337039eb4671305aec70a44af54a39175e4fcd0836ab9f7ffdbc50ee2b21d32249787e6efb8e4311bc01ef8fca1861c63d14300a5c510987a653458033aa802ef836121abeb736d8f261ffbe519577c513acc78142694c12f5f0c6d8626403fbe7a767ce8aaa44d6e74728679e62c3aa09be295f5f3204e97efcd371aadf92278308fe11fe783a4cf2fd41a27c309af9ab1644379713f0d2ff296dbf3a4f1cc79eda4ec248e0cbe195336da33a2e713d613e0ee10a945ae7ac27d830e4e072282c596b43cc10f994a5316bc7714d8ea7bd70ae1580a6c6843a498588e109dafcc7df7be6471aa73c684425d9a0da82e7b779691c6d3b57ca54dd1b33f898b51a850f7324fd233bcea808bbe92592c1dff543b6778569ef1d780e2300173df649d349f94daa6d79157bc4e1f0fa6d87b749c1d9a1149e3ca6c3730daf07c79b61c3d5206faf7fdba2192e1ba2a7348f56dee080bd436aabf03475d61fb7d7c0cf1d53efade02afe4810ebb0ec9bc930dc737a1199cc1b2be32613b71eed280f7a574e25b34123562d2f5792848155eb3ccb918460fce552b02f40af1a30ead2fbc66542bde0281b531da1b1102b4ae26d2fe35b89f7ae7e0609de2492678c966e4a2f01450255d170e5e6f5c89be89200353e1602c72e7f4014c4862a88c1aa8ec5536a1f88a83872a3eda54b4521f7deb3eb45a4c444e49c655b27b80d71419c6f79f16e8a7c923b38c0ee35f5ffd8c30c4bb4ce9369b4376fa196fce1c94eb7ec58519898983e3469f2e9a17289b8f5d1142eee6b8b286d67b17d87958e437ea974a87adaeb28ce7e859c64656395adbea4873ec9f1a5f4ddf1020df0ccbb4d1b3250d32fa7ccf0a1276d44df7a6434866485783d5fcb6cd3c71427d510177ece24d1a5cbedb66a79c236dc7daa22bce7f0083eec95fb6b21bd159c4b0c84a48e7308fba0be1759dec9b3995d7709d76eafdf694c773800840705b06769659203bdb3e264057a369e44113b149f17500de54c30b675ea7fdbe33c635afcb3b8833a3c81700e9cd0e8346fcc4f9de1abeda94139e64cfc5bd82ec40d09f388cfd9bf6e4ac16d4fccad161e3f3d8ae5c257e7785cceb4ab680850c2c6c603d72094dbfe20ce391ccd4356ab5d88757998df89f212ef4f226a89b4d25cce956da382637258c7dbdfd00af49d00a8d8a57af917d83362322ebbaaedcd01650fd11ba6ecb091ad919e4a0366905889c2bc7282b0db00970fc0d65be084443cd9c07657951698f252c48395d7bc02d584ced844bc2a87482b08ecd8de08351283c6769635ec2f0d7c6dbbfa84169e7ce0f7977a9779ae92f1071f1af553703d6c503d0d4bcb8e6c65523d41335189dac6b0a63cf64c529aec58111afc3257576207879173a85231e34c18effc1446d845e2ca0df378ecc6a92416cc5c0b83c8c12bb41083937dfb9692883a659b1fa6d3662cc608f83ba412d75c9e3be1e9a0aca5c054c15046d32fc6080f53572387d2d60ac872b3fdd06bfa53b1f635c3531c46f95b1c87d535fd2c3f8df6c690bce87a4330c17b57581df9f61229b5f6a53880115c6f8a8e7d35e5101096ad454a2e83d465171bba02dc8b3303c816110f399f026ad84694a87ae8fb721aab09dac0d46f843e6dcea136ce586e1406243771c64225f33e29ac528f47e9e8e8cca78cc5f08f8ce265acd8ba2b050e84c74aaa818ca55ae9d41f7bbd50214e48672ba1c333d9251cce1a4a0cdd2ff18b62f0d67684985878960bd4413c227e356de8e651bf0d0cde84280eead7f374259256f3870a45efd7c98a369b2596ebede75a61fba899b87d6c2d79cf6d6df8647eb9c646f1d36058150299e7e4ebcd30fa45f507ea3838f8e33a270cc97262cff02ed648b8cbb28;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd08ec8168976a53dcab21f96a956bfc8e9675f0cdbdf1a9ad31cc70d7a5024a982058bebe778e71265dbb9fc97324695afa303d0e27ed5d648f3ba191bce51b883264c35b294215bf8b58cf3e3203ca4b5829956dc1f72399788c8256a0b2f5340c8917b82768368073d6d3fb34cb322df008c237e8d8da36e4d4f1456d5ac2fbd201aca1348a4a8114bb40e98be5920664200c89ba84337ab5fa17a79bbc4b267eddcee8fdf13c3114c52a4384f14c470b7b6cf66e561874ce9872eaa18cc7bd2f8602ce4b63ba034f15ac2875617a76550d43204163d97acf61b8c174769462f30f2fd1b8d89f01a5f297aad2e8a9c1c01491196caa07e0415a1b4573fc27f41e11f56af027d70b8ccef6e750637fcce8a40339eab35de46b34bef316a59e4f0bb51935ec56c9c200cb6dbf05bdfaa59261d9ea49860667979804176ea7ad1f35ffc67c651c7fed23eb4eb8759978698cc88603a87a1844c9f26cc95b6b8b08dc241bbde30618dc20cf09b806b33014ac0302d51acbf4b7c7bb3a337d51848cdffa965d0e946a8ce1f2095b1eaeddf6e92b101d9ebdc2b9df1587072d1569885ec2b82b9f57c80ec805d0825908794639583ef834cab5ea3f20fffdf3ca8e20bba73b5d0f11ddf734d564c361326194b22c2754eed7f7ccbd87dee49ddd3157e2f314e514ffbf0e1b1f18342329e3c81db7fca0f802eabcd634fa3f9dff5ee73e178299f46c0ccc56b830cedcf29a689110c5dccbc38e5b915d18bbbdf25ab7cda1e4def20ffb7d2aac5200a4965371b3f940c882515528db9eeec97a0f6174f8056694771f5826097dcfc6f72754b8592c0ceed69083602c3f35d15784f70b8bf92532c2ef2901e8f4a37dab55ecac3a9a6615c095dfe254a2f779928f36feae9f411a6bf5c4f4db0f31349f941fd2a807323d2fc053b298702a08f7575864d094fa5409eb7b58c2d15ecfbb99d77040373196092e33f9f70cb955dbf389da9a8dd715200a7aa46a3cf8a92b5dd6d84a09e90e519b5a62ed82d2dc0352e4a225ef68567ed6b4e28ee217bffcb1fcb35c4e03959c1fe4d02b0f34c5c58ff03bd4f6a8c3fdc38291d91a6a3f272566cbed5466fce8c961c590e4c61cd585a527ea63097971b715caa5b4623295f331ffec696d72f8373fe9113e334aea25501c46f58e8e7f40b3c6c374a0e0e198a75d2e3196489afd446b8e19dd7f9adaeb1d2f0f9548ba9e892897e518142db7051dc7ad03a20aaa2087a48b65f47ffbaf18d7436534d8cae6305a32d1a2daeb865751720609849817e20ed36db26e1e9f8227a1319e2424f0e3b7d8ab9f8b49052cf949b5e3d340f2421ecb7464038496ab650f292ba643c7148d7d1535468fc59d48b7f822dc7fa06c0475c456b50409a35999ba90a3948d73f822b5a0c76db8b461bb4bd575cf5265a38a1b596c1b38b50ef7748ea052d757ab421c215c6b36919cc91f09dd0df9e942611bebc24e6adead498d5678b126f6ec0d8c7957e87d6ce023916f4631b29fbc1d257600ae67f2d0f29fb50f31b482b6af0fdf01280a891617b60a04ec71de3257e519e905a6fb4ba508fce7436dc3d5efe2d500189fb37fc6e6d8023539f1122e5c62506b5d5a36b38c1c9593ca02caa36ead1041a767158b82e2d70db0dad182a0b973992aa521b394c69433a6c407859847659e8011c6ad3ed18be18c69ddd01572340efdfe44f5e1da0db84dad8ba963b8364629bbc9da8c54049cbe4c92edc9e22a7a32a97dcac6a057ade9e942222abb97bd785c9792db27a73251e460231aac127e3b63d564e8bf7bc76cdc7bd4c5dc3c022b081f053de53e5dc9c3a5d00b5bfa5884582408bca3f46f9b56c60ee9508615afe5870ffbb6f726ae040de2ac6ae28cb17e0dd1d0cc80fe64c6daed670ad43df482e7bb8d22b1252e6b61a9186fc961a826f0a6f2655aab5bde3833636a7e013e8ceb75c1cd508795d2e3a014b289c480eff10a8f484f689b15603ce88ed8f87cfa0d7010870fbdd0411fc0827db7a4529ef402966c1ddc9c92bce770627c4877a1516e6203399661d08ec7445f2daea7e6ce54291b206a46f90fc05695985289afcc1910cc77ff38c4818fd3a1435575aa176295ac0e6a67d7911c80847fb9beb3a622f79ecd976166524fd05846b004e5703cb0770bb61b79cd15dc80f76bb1eba40649100b4832fa86a8c3387df85cd749695c44c681bf40a5d681867889b7692081e5096c69ce11e9b4d5ebf3c69face504ef4d06941f446cae045f053532b93b8fddd22404bef77b9317c152fdabad638e4db1e4ba18ed4147b3febd81b28ab2f714c8d074a8f54e0a5e3755f1f15a86528d836a711a796f3e6c6f50c20b66c1a13d2e184ddb30b653aa22cb1bc34b79c9d08cd895dba595e0b394f1638196abdd18dda12fcada4e75e42fc25b86898c8ab10b2ee000012201ba7e003017f6197b04cd9e10d299739aa39b1b0c37f417d66376c6fd5d195e06c55e5aa34d22b20462388093442e77156d0fae6b254d0ad04cd36b5aee7ea1f81ef0d7d2d15c2cb53bf978ebaf08ef24df5a4bea8eb50417756b669534f7d70cdb1fd3425344a40754e90e46b46b625ff2ac3d7b5878995ef660e5cebf4f56cc626c32cc47439b5080bf71f94b8dccb04752f8d1df62cb3763722a70173d0917afc8ccdda9cd29a351e10f13aca55e59bbd01753dd75eb8be44af8713dae0b6da7b66b0b02066c2f9fc7e8351f8744a391c7f09373c0084afc1ea6a3b0492209139b6d6701466582dd0b11e5afa4da86e0da5e58a25513b66c9f960e275be7e8da432bfb67330d8d1c1cc02b10d4146ff6c5d4f2a585b1eb7aa37467b5e3c8c9c722c4ee92f254fe3587df580d0ff0e1c650ac71bff0b883cb73547bcf14070d451ed047851dedc048ec3fdf3221a16c8c6bbd4fe4e9f9667a27d1bd3500e8ad3788e27b8350bff7e5ab1e96423ce728fdef09a44e1225c01f1707eee3d01b9b95cd3797567e62e523887ec19d57363f63c6cdb3badff0fd4fab5f872c0228c44cb53acaa1127ebfe9715a9905cfb8ca6e49dfd0b6746116e60e68f5e5ed6b9eabaa39f6c4a8263933624ef9fda175a6495420fadc2366c15949499e5eca5456be23969f88ccaeb2218d1ab20eae131974c0c604967efcdac69009bbc38818704085d2aa89e2a4a3ce5e8239013106dcb273940c4f955e7a2db43912aa387d0357739f400e7e69956da94b315bc4e784e45df8609d917942f1b774f6a94d9245e3931565e420262f6ac8c5eb86a9d16cdbd0c5b1ebf6cac27e6aaf14b9c3cf662023ab63716e4ce6d57c5f7c5d5d9aea18a71e60f2d4e7975d94be46252a551026b91680043f1a68222e4f20a084feec5cd162e7da2593d9d23a5805263eca0b1f776cecb3a153af77ba73b372df9df0fed9b6fc3cd5e2234e52c4743a794743a0e1d65076b879c8f8035ed06c508a4ebdddefb6184dfc6ffed30c1652b9ff3dad0347b8a2dab4a0e9e6baa32e14afcc3cd2b57dd90bc88dba017c5b068f1246b919041fe31e3afb72ab3840d67216b15cf661af29e8ff1ff128f4f7325c8d4eaf88b4a6146422ccd2596e690334e65e2f37635eefc5b02b9534f037c90b9ec4e1117832114aaa13d4442adcf85db33740005b9a2c0c81cbf8e808e382daa110a3cbe07642c45abcb9b32bcf257c56cc4ae7843893a6da4cc90919205003be518aae960a3ad6061de5772ffc5dc63283abf509e32276e2337e3e6ea290e5440f0d972c3dcbe5b2b92f75919c89433549c55bfb78f8aa40baa70cde9c3ae6774613ea66168dcf0023f56d29a566f30dd5fe528a283a0061a61aa55aeacb6511384efd9fdaa5489fba8e2d2a651081f49eb2766f632b18b370f5c597d3c47da9f9950b988978bb7c1a29656825148a04bb057909ac55521eebef69e0c57e538b1ec29527ba417d99713c9419f3ca31cfdc8e3c6ee756b186b942e9c2b08388655a1aeb91c3df0f92bf21a4fd25e96ab0ba6355634fbbab248ae65264c9f8775ba0316c2eaf27ebe67735eb775cbd8c79de1e8ed4982dc2e5ab9fef596339648d33c0257668fd01515874e2d7308a45dcf483d3a634b8102781f1990dae3304f9d73fec88dec23a3b734bd86ba8f31ab0f7ea4b6801e0628b89f665265b0caa0ad26387f175cc8ded19ed36c6f849fb12e7a029c139ea0688c3b3608ef08e3e73ac9355d097470890166a21676ac4bec057b1e4dcb2abafb4c0a80cf41fd0c49afaf6f594e74b1a0ad5bf249ff2e9e4ef0efc15e9c78488b22fcede672c65e20b082acd8fa8f07f42690e73d5be59e4f595e86d76f7b23b34bd81e69121740d642a7e478e549d0106879f91c9d1d55cdfe63a90ca80fea3c8936e5827768dc3a4cbec14d7b1dc9210ae9094507de3b12360335866c1478bc5470d34e121c4bacf09145171c46b099fb74bcffba9faaa8e27ab6eb6336393915c5f08e7204e49a6b5c48f86acf7b089e47e9989d75672c92ce0f13d8dca7fc363336038022540d6108c22a68f33fb797dfaa1bd5b6c95b1f7f0e5bb5104244e37b4cc024043185b5e0a57b0bb1f0129b586e8bc1552a453a6f9ec2afa8f80cf244120c55aa00e0ac153ae7428c48896a98f53997aea7dd2cb79e8eb4bb5c69d8a427ec1cae345b66839c4afbf7919ccb0c603b01606a7b85dde7432cc8e9da6c635995eca1dcd306b0d25855aabfcf954a47be30b5ce0a4cb857fe88562948dccf1f525636991df870ac5786f3596eb6d70ee970ad5ba290d959486a1db3d8c24a33d90881bb9a856d1cf2bce5672d47d22db667ddfa9cb65355e946709a754035c224063e1ce3e2d15dd33a9e74be6b1d4a295a0dd998d60321af6bbd853912d675dfa082f8b04a10026eae92c7acb0e2dba007230b51395442d2c4426f8dda658f8fab5f7f221d451f5e4b6fdcbd8fad40770732f4eccc73fbe969ee8e0427de6fa140ba3ae262bd8070eedac2439f0fdf418f23041248e4af74fd9b9ddf5c3174e54863e49045b3c193433f4b68297253a5820861a8a5d2a896788c7121d16d75138b25953a2279a6a63555fd91c9d0a3acfb2a2e708d68200e6824ac003bd698a4a655b19829b38c23f06d5055da0ef1beaeefef542c34aa55eb0a5521b082dfa99b3f657f48a72b349ea4a5cac44a8d2670720af1f872239f208a1250ce0435bc97d58594e3dfbe33816c913a73d0a75637ccb7c0e64d6884c1544353a14a46f08dbc49de94bfc2f1977ba99f4a8e4f32feb75614f6eaf9498594b9a9fb2a0c61ec147a1f26546e3ad6e8630594d8912f925447a3a5601d6ccc50edd602bdadbaa0201cd04163252b64c622bd75278f6e20ee5e9fcbfdd9929ed7bdeedd3e2b50e4a706b1406b8a94e9729964dd3c61b6294858ec803beb1036e0f2b69668f80c1b45192642a6fa6f9a4031a05786212121fde1a4efa361c9aa07be2bfd0c91905ba1bd24b106a094a58e388ba8f6028764dad43c34c3becea899eeeef887ef5b97ee19b309e15bbaa12eacd24aff7620095bc9ac915eb334d422191a96b42542745a2144cafadecffc52a3ae14f3df80a944acba84d47b63ff139cf2a4f1e9770ce83dae1cb21994a6602e24e12b50515a8c3c0d928b4059b0b96f42d7204a0afcb3fcb2b5628b54c0dde599cd83d766158151d73109480e690e7fb2e1f344027b6a0f4388c28fa21068faeb9185ec8b3284b835699e48642f2f8d55991d1f581cea229d0f20862a7e41b0156f3fce1ee7e847fcd37cf5a11697f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h2bc4e35b5da54e20aabb0b285e99219a5451aabbab57161ab84935e970842e1fec2c4735a2fa8ae5b06191ba792d05bf4cbd8fd82c36966d5cdb443a61705c18c7cd77553a8c3f026c2c5f551f5c6af0b6f9f997f1f7e408c605bc862188a9c069e9614cf6dd41810cb15b35ead689f7572257d9ab87b605f93b18c13f95d0943a2304d32d7000f067875686468c157824cd67f4fb7e67c03ba3d4a0e1645873c04c78d0c4c2fab6ddb2c1a5282cfa884e072d37c62e844a2be9db6e72870137faf7a37793ec9ee5e91badbbde0f1a032a22cf97aff03a25a0ba2c096099272bc935590b59dc088e18b6dafdb056db765980b0c11b6f102a06c6814bcc591c8a196fa3906fc2dafc03f8cf35c780d9661e3ae3765f72158f22fa7908ce16590eee16e4a290c6adbe67cd5470c6a332eb12e84097f62d945b10e314036dfd765fb96a293d8e74f38280bbce3ffbc35e481f84de879c99fd6fa6a54db97f01ebabba80ea5922fe578728e75f90e852f7babce43aae4dcf1822580da6bd1f60ad97793b1bd74e6afa572c0d6ca2ea4c00217e5102fa85c013ff81349ace565723143d044bfc88ab2b5b1a2fc0254adc35dadb0a567e38535bc2f9ccb614260e8c0f261f27069a10d54d71028111971fa64517ea4db93fc547856468238c51549bc925925d35bc7f7e49825494c1e48f7575dcfe5437aefe4a02cc17138b3774aa45d967ef9a6b885267125059e1df0b367fecd9befa8a2b280db7d007605ef12bbfd1822e7acc570ad098e12f7b1be0c695cf950376697ba12c6054123926e391c3553d47cd34c34b7962e9b8425ab9b947b4373b105ea52169b280b0417628430b4e6e8b9f07c5773cbd0d07840850b3424e2bf8fa06f4be06599f543798db630aa11628caec315dd527994ca9e4c98e4efa4891c4a52deef4f18e28209e455639b2c4c060628a7173cc9bab0310aa26e5c75effae664f3bf7ccb683403e7292ee1d37b4bbe013bee2dc7939164850ea1b9b0eaea0024f51e05ac0361632cbee457b232cc43303cdc904e437bb2e08715a4a1c1bf9ef7216bb9453cd115049a3a5e8d595c56a86c31cfa6228297b71bbd2f8679ae447e90b4a5214d42fae2f62355934917ed288596a8571192ab12619be15ba9d5bb7c2e8d4f8b74726c142f9e4c61690a77ce1ed544718ddedfcf5e662cdb0f55b12acf6256ad53413b915a54f3abbb237e35fb6075057f54c97f1fc9ac803acda4afc76a07647904457e14a3c8de9f0b07b9be3fd7fe112fa85dcebf0e97d749c0df1fa538ff15b40f9c757afc88013b7847d0ac3312f88813f538483aba607f5bae00315295fbcb00c15a503bbfdff4b54d8cea3574ef3b5683a78ec814568739b599df268e46a1909dcc8458d1804abc0a38715bfb2aa88df3aa69ef03dadacdcb9f4f50d85fc6c2cce442c36c6994685092c9ac89b6803336b75539162d0311fd56b25f22caabca84b459011c6d273ba45df5c41ac160d1696a38a0751e45fbe8f8c56efb50718a0c5e60c93df0198af973e9f233fc197999e34a78dd6ddf2ffcdc0630087861168c84f5dac11156a8b3df5d3dea678bb357fbd1c9382e808598db3583ca6edc096668906cc84ab847689529502afc0e0165ea82ec628a744fbad68db85011fe5d1ed0d020767020282453949502444e4f86930292d08b5fb2fc59feb420f9725112c4a1b8f16888ec875285ec49042a69993ee247732dd70def6a1a7a1d7ab89aebbdb77142ae54de5268b932ad3ac3b6e84baa083667f3a3a9387fed15586d478aa1d3315c184297c3ea8398c0c889727dc8a5ff43fe1afd4ffb1b250023456dce1237327c8cc7c608de040a6d0a0cdb74a829a4e17cef538dc80d55fe78dcbeea44cd6af63b2a599810c527d5ad9e9f37847ed0b80c313be5acdb2468d51b8592c736a678ba3dbdb92554dd8896ea81aa0b097a9c051a76fdb580409174681a3a4726ed5991796a3e0dd354fc3a1e0ccd8891a4edbe36b58084b6ecee6a84ff8515632c989c63c95003dbee288827641404f132436d77114b0bcef5ec90397b434996757c99a9fed9258c7daa22b4034a22a1bb16e8f69bb27bd537261bf0b6a337c162e74f614bab2d4af094be485530a5240102f4a36eea0f3f6c8ded803e1e25e3616f1eeb38a8fc871d4d71a185036e1f1ee307ef72e1d296744dd653280bbf41c866292dc0dea1eca2b6c99ed8d2952ca7af464e8ab447df60b144004e5ecc118943c8924a130c260126c56aeb71a7607eb59c13fec419c28438c70de1eeca8a550facdd0d287cd8a90ac3e4392adeb98cdbc54b91bbb33202fc349cc316277bdf9a8fdd49bf31fe45f826b33154c52e255a9c7ab419f7b35973268e1a3d20fd9a6a68c1366550a866c42baa7bc482eada69523ef9f46be64202c7329d6e16c2bab23b6744686140404fc7f0b0e3b410e8f7c3ac5d3dd7294450d60ebb2c2757b81fac1fcd7165e9d97db7bd054f8262b4fc77900f7d8f741427eb513b0ecbedb90bd25bd07ca5a2238f4b72e32fa02dd157fc52a48745d1664605fb76e0f3c205e4f50f0ac9e81e24a55decec55e02092a78794d964e0c59107a93100c544ffc95130e83eb098df565e189dcf6f398cd62e18ac9e78f2388fb85b30f5e0c9d53a2aa9cd8449d377c67ced13c1ec30c65da46993348d843f7ea32de5fdaf59eb7283499d06d229fb5e5a58238ac1063b68eaf9acb4fa5eb2c2ae0b0ed40b127980818d4fd6053fd2be76912860665959fc9deb0c77748df42a500398447979775280cb7a5f4925d83b29fed7662df635b542937b9e7b4fe3812111c5bd40615e47ce3241c4dd2d6ba4fb5490bd52ec77af17bebc29dae973a4c3ed4bc49700f7b1b1319e3aeb3e3ddbf9094502ba7a650350c0a433a8d027541fa39f68adcf17476a7c01dd68eeea1f3ee7c182e7f223b7cd57bb61ac5c726623e1f80326e65bc59e37b8b8c80109d2e3d40af0046928e2d53a17df0c3a087547ebce7c0b307e23f34a740a3c0ed9d6b6cf4477270fc910b44a62c67681c03639ea7b59aa1ddef7c5303f76acae3b71760323060ca433477e21fc82ca0ccb5bd00a7371b7da9924fd26d975625fcb1fd82958f6a7ddc6bbec88d31bd0e4e452fb08c945593fec94d8ed01aeefed6f2a6e59771fe9d7aee60b34bcce775a813810614c08953fd1f0379792da3204fb7cbdfc648892edf2ba919c5c4c8ead96bddbcfd1702b17d0a7a91622f4d40209c25b8928c2d307fa31e6234979ec5591a1dc66946451aa8a1db368b54f16aa6d21fd7877f9fafbbe4ddac25a088a6954aa120d77698b1feb1ee998a4312faccb9ff053d9448b4cfc19e523882faa33af395994626912fc41fb40db844c71f9caca0bc31580b549cf9e38ced90b2b3711862bb2967c0aa24d60cb7ae67fec2114f3102b769b4b4822bcefd97e7bac024a6190abdb01e44ee3d8c8e4dc94b6e65dcebbfa68bbf842b95ec533319a22283413644aaa89c6bab5318aaa3bf7afee5fe4c636d0ba5a9740976411c330d2da316d084ca5bdbe052b8d3988a7be7dd92e94de4b9cd3f5768a5c0351a3797db2d456b0f7c06f82d5590e997a9f176c1994430f6b5b2ae808c9628100ea696626becf7a5d5f7cb72e782a9d283ccfd53ca51a8cb1abfd49225b954a7f59d3761eb65ca0968abcbe2075c4481afaad3a1239511baaa245f6bb7c2110ee06a899b17fe694ffd5969cd2fabca9ee73cd385c58a8935c8a14e7bf988f35ad4184f40139ef87b5d03e82e4d8dbc0bdc23ed10021ff121dba99562162a09746e3381d13d83a8d0510a2c053c0b409a4617163ffecb4a1dd08034754072aa8366086157ce4e940ba92d127066f900826da448255a7e55c51ab6ac7b911c57c1fdf34910a8190946141cb308fdf9445d2ee92ccda101079d692dcfb3bd0550e80a0c91872b038accbd7625c2572d6fb97abb46d309309a59a09f607713700fef1ef4755d7ac3d3f47135eec76b5262ae429c953fef288003164d7596baf83a4112010199e465ab167273f8ece0cb09f5e235d1d9daaf24dcdc7e03b0b3a63cf560be026265d9127783ec347dab747b4a54c36a1da18d7eddbe097e2d101ea3ab9abcaddcdd4ff32a09ac54c80c5698e91bdcc8043d6a01f99e4c9c1d7c51e68677a9027a09e02f4ad4ed7f1bb19b208e5ca0af796613be22ac2dc1fd2bf3b9b502e48b9e28722e26a8992d27c405573c5eedfc7ca62d59b28a686c6b2ace1b5ac1775e397ac8fa256027c35c6365f38ca982c183d1e1335bec467edb6fc5849ed2191a62de86704504b6de7d8eeeed566931a4fe2dfb74fa7fca23aaea650c3f5c1c73123300c2f512904b784ec179e49f990af7da0e90f993685189341ef75e243ee303eb45f21f1ab693b73d0bc430d4c99e05a04d24a5765ae0c6aef97ad3efd073fd1f8baaca169d060feaa0e60bfd99edf9a77a18e5afb7de1e41320adab63b2b7b1c4f330c32df941e25fbe1892a6f64117be5040c607441dbc49f0ee70b832943b04a7c71f5a322a749d7db6243f41105294bf6f6acf4cbe5af5d835da4e465dd224d9070b1462c6459887db51286edabc03e34821d7550dca084fa122983595f88254d674a4b8cb1a634844c6c9692cd24b42c37a4b4cc12715bce697bb9a0bf18e1fd49d0d3de9e317147fed6818a201d8a56f454c18afde5473847439b996b34b5e185bab8b19fbbfebb622408a7309410f1642f8d5b843414bd9d8eefbcdf02bcf08da28d41bf82bc64556a5ba8414490632128190263d14b174531c8910379b247c15b7baf8724e184637994c9400b43abdacb444754a33fddfc512ac2fce39e26cec676241fc29e23727b95949c372e0617d79d5ed16050f51712fa00785769f61f22ef009e60578f5409ebfe51b75f71519741617c428c5dafd6f530d96844804ae19dc79e2bffe925eb39484db7d3d0ac0801223bd634fdd283311bd2e865d5e90554aca1cc33bc3d5367282812f5f0c73ae7ee62662f7b80f14686afa89d6a5b8edcd571e849c1c416628629568377c092ce26a7d76de25901fe74b46050ed954ee5baf56d82902bc698dbb70bea29017632869caaabb7f62257e7f197df8e91c5e1d59926ccc72f71b67c8d9f19617ac2aefd875fe974a2e9b22bf9e2b0ba78472bb739e123a27d6a3a8f2a182dbdf205854b87275c7c06e641c912a2e0d7364fac6a67daa3779474220d436cbb5c510f775725892df4c5308d294df562d22ac900650d30458d42ac9fb1f25b42cf15bf707eebf6f21d191534363e1a87cd202b2b942e2927a8df42ba8317124594810a0c6c8ff6eace824f6f26a692e7bd54918f1d831887477d270c74b4554137946d0423475f78cd3eb3f8ba7f58723e11af6bb14ec7a90ff141ca638a470087fa0c9a72be995e6ec57f9e6699547d7df9a6c31a7532bd8b9d9130989e798257394dd2b726d0aa5ecbf3d21d3182ceeae959700b88355d980369058b30e32877104de13bdca68382dd905dd8164e782f717205c44b53225b88b3887dca371c022db9f0de9a5be5d0a765f706719b59ec89ec5ca19def76f174f437de2754fc08a079ce4867954716dc518c00e4e5c9a651dcdcea17bfdc1aaf4b58a8e4dcec117f425b327d9b8f494ac87a69f3d86b7e17464b0102015267be0e7a1294f5521b85f3ee431f1a69699bebe03d240bcc555ad77be75e04a4f8ba2cd583222ab7e303acb252a0830230af5bce1db5f46dfeac20d95617bf15;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h984361d2252422d380d79d7be54c0ecf3cf69898138eee3a84660cf416cf39236ed83ceae0256d2185a0038ca923f5d211eb0f409f6aa6534de94ccd9050ac933727713d09464fa2f40bc73fc2c46fe1d1c4c745fb70421d667f1cba64674e3a5a25d2734a23b42cebb1615b261b099bfa84b00fd652ab1fbbc271f4d99ed209d9b3518e4bcbb9abfde57323d153c93a19a1767a53bea0284c943e724529856ceffb2dfcfa86a127878d8376a41d974445075ddbfbc34b2f390168183b7d0a65716115b060265a3fb6635ae48cc29f6ddc645647fc071519e21b615e9cfd73889747f79eb78443b4b9fd234f7b84d7718be9904110db32681c9152e7bf62013cc62cc8c29db8f819adc8269ddcc862da278512c631b3dde6d35d382c9645d7d3355e8742465d80159559f7af3a118beebc0034fc5b02a155b8e182ce8b7dbc3ad6d5cfe27ccb022afae042289871e1896ab9f4b87e74ff4c30f0b9c78ffeba2a455b12812e1e09ff3c9d480e0c8cbcdabb3ea19a7154b092c91b37ec4f39b5fa5c405d517c96664e88f812dfb4beb6441da6b7a17bb1ad199487f0d5aa5685f4a90000ca0f9a86e952a05eeeb0e89603816d4d730f5f85acbabcfa0c051e9816428182e08070b79a7839e1e94a608173d10afb5555f9e9347439f007e66d1bc6b67fa643f070bc96fa0f49e9763268f3fd7dd8392fd27fafd348ba5aaeec4a5556e3f24e3b7ed8f38ed71f364519fed455b024c0a9bb4b4e72545219de92737b2189c13ece633a84adeeb180654743babc6f52af3695d7d1d0c56322aa1e0034a6e09ba68b22afbc1933132e41674fc47a2c7b748f86a9c8069f0e6b1cf6df11911794cfa6fa3f953899c0acb754275664d91eed23e5dc39eaf76f5bdd390ddac683982eb280b754fea302285e3751c1b472fbb13454cfc9eb81881289f0bbee35e038396bf1640d9fc4de2f22af895b3868880b13cdc1e2acad721269598ec342c81e8863be75b1cc768105b40f945163ecda6514fbbb9fc991fc95d8a7a91d73ba29f872c22236b52f267e181da9ffb7da467c8969fdf1e9b08800b2cc03eea04ab5767cfb951acbabc75746ace1ec6939f57d3a2187904c4db87fef1b9b469246128d23fd2a71b6a8ebb996529aa9ba5c837a64938e61556eaff1134d5ce2bdcc323e91bd0001825a534e59944052c320ae854f0b4f28badb478dc7e6c5e254adbe2514ff64368254eaa876ac61be34fa8245cba86a7aa61f281518bff8d2cb7207c46b325d4930243451078a9681e21220f774e0703079ecbb8f7f6ea206ece5499ac5222b6a34b7a894f10d21314b95b202d8c30168b37f5efdaa60e1eda8ebe175a2bad14351fc098211d9f9c905532e7391fac6b0d76c021f25f16e62ed76b315aaf4fcf7339b4d5109b4595ddf01f27b5a963f1943e1267b333ea85ce3b3d10c8dd6673097d5528dc34bf602a8dfc0f6602a91e656eac7f4c72c0b2f3d25aa4ed2411240c1c342325c50fb53db405f9816f14f6c2a1680a02827904d7c136909a00b5950fff3d1797c5091366fe40eb8df78853c1dfded4668584dcd7bb91469e61b3e6775f354a5f7ccce62ad5b9cde062b738bb3f3f69d6616695754bda06cd873938242d170a674d347ffe17657b61013f5ca6f1062e528409f72562cd3c93654f78c1f964326facee7c39df12760befb91e6e631029596699e31bdb295083d4824588fae933ebf3a43c1670321d00864d8d67d1930834b3a584f07911ad7f33c263b8f5609e3ec077c9360b608e86b9a59c5e924bbf223580beb984aa62ddb781abceabbef4e4322486dda9d63049d6a813a1ce913af49d34d5216c50640bd2ffecb4e06e3bd2798756f83421f7d84e6fe53d167b76989d717cf52ebd636d1d56ef423f84ccfa4602935f04694dabe675ad21c8de458e1d4dc776dbb5fdd3bce4da0af70176c235ff30f2ffbca9f155be16433b736f05c73b62bdfb3593f18f2d081a55b16c30ec5ceac273fd8f5b15b96d25a1e8ca45fe0004fe9e4f177c3a8bc2c20cc14ce9017ce7bde9047dd4184f1bacf73b25111e287d07c83ea2a4e89a896270be4a7c1545598f3fda876082efebe759d05c1ba65b932ca8ff58fe33a2a28c631e4a65424c64e6a51a83e5a4715286dd755ac9660bc23730f0960cc8e7b4fc3d91f797bbde2ffa489da0352932f23b970687e3f199e68fe598be1306e32629eaa3757c80b6101fdf103cb94050584c0801a1a506d8d20cdb8f4646203fe9b47e29f69c5ad765cda582f52e43d6c9c65ed1c14eac156e66964e368b75f6ec4cfaca09a9ada132e2369c1c6954ca3121ff64368ad06a9116d4a2448ba244b6219b1a2f3952dab61db95974c342fb93ca613e7d57255ef9a760e3428cfccb8afabec4ef0b3b4ab5aa2cdd01ab270eb457afc9440cf0ebaf17c24ea62af8a5b1ba0ff8ddc0fad163ddbefdd83e9dd0b468efbf705e4cfaf78b21810c5482049e29f5237618dd69d80d58ff8c0f35c193963c1bb17c1adf682d38ab6318b6693acf20931cff9df3624ae8f47b2772162a1553b88ab833dff49349ffd7cd6a137c6d5d05eb75ae06a6847408ebc943adf47b68b2f7111c456925fa0b69f6ceadbacc2cd689ace3bc8d19246547e806baf77c7f6520bd4c28fbe7ff9d90b9f6dcee6ad1cb9ff89dd28820d5391646c111e2f0829fd700df92336bc54d1671fa28f2e605fb7fb350b27d96f68e28acf81b3c6ab9dab9aa6f7a94e7a9bd8ffe284ed7f7fe6fad42d2a3c6d9498d733d9bc1e737ad6cb6732a4ae6602b276746dc5ca5690359a69a1710953bfc8fbe5034c3386f949882ea1537d9b48c6da4f86b2958aaedd59fe92e56513015ed292a30496be7c466a5ed6c1f86971b1106ef787a00e8eef67c787f25c824fa8aa19b758b108dabaea24de46117ca75c9976465b38939f6eed11ce895cb77532b9f9e06c2147a00860d2f0102da257d8c5dc91676d48127115bb43d6727bd4a6d7de46d1ac72716e1aee41b5f678e0dc5a9e195c2a3009ffa5743a1afd1af11ae1498c4c530df8c041854b6da6151ccabf0db8697336a4de0679a629a263f9ea5c1dfb9d4f0b24cd38c0fb1ef1c8c8458ebba849d20fa58bb6674b56dc8cf1545d0209205a017f6d8fb6c00b2a5103acdbd69778bacdd96725495ca82acbe115d37dd033c2e52f4660cdbae21db20398fb1acdd11f04c7a06c97024281f8c8b0cc6439b51e6c820409308b0cbec24716306a54a518b17bfdf51a3bddf8c72f57645f61e9e541ca494798c877baad5b86260794378f8eac507c0fe85fba1e353d390191ed101ec280b5432d0abc477d9d1f956c532aa10e6e6e59276e7f1add59ad514bed437a828ff3401a67db8d3824e238edb01cee0f3abef915d2092715ab8ee75822be0cd3e0b970e40c4a412c05c5c99a7b125f16ad2999316a39ebd7822b424209aff0839d37d34bbab197212262f6e4a81e619faa49f38a0c305075d04b1d84363005f1b69b7004a4e2f9388000f2546df797211d44970b0c2eb2688950d617d54278907dbfcc8f631e16467cd212638e8b9bfc81dcd11d2e2f47015057d85e7a62399e5377e12894a02155ed63c0df7075bb6d205ae1dc2135dd38128d84eb3e1483734bc268f1deaa71695d247abe472394ba9ed99bf57fb3b719cf6037364f99830485350db4935dc10a641928fd7e65a182565ed5df58503a8e66c098b73839c001b1ac2592e711b296f70221caee40a384202b450bec16d5cc558523a10e0c5760e377c7f8ce98b4ee1266eb1a3d17b3173ac987f47b320782d27a8ade3f51eeeb466a0d238ff24ca694a00c8d586cb5877e77bc1e840960cef6cf15fb8e644abf204024039dc5e3adf1d244044358d36b480a40541fc88d9866c10812250bcca2f4272dede07cb2eae0e016f1f0c4bfe5a7b60e9661b6364b031b31eafcae54a47526ef4cc767009d0f06408054d439c6f1b11c63f14253814e5605c433e49332546bc1369b27beafcc378922b369abf49160b332d57ce432f3cede6bba81ff99c372cb4ec4d679a1c9da70bb566145124282fe48764453cc9953afd9044ea934df099e44f63eba4483c6e53a226fc39245bc90ec817b969caedd44f062614f7d2ea619b61fe0dc3273d81564f1a464720d0e312bbbae566c8e7043bdd5294029e25ea21a9785be3598e5b06012052689bbbdb9a4887401b779f35c6bb41b0645f4560a1ba2383eb06353a69a78ca83a34d91a2d7bd814ba0c156edc4109c02cfbea12acc1e5743def147e46c13ae576ddcaca84a94950f97e162175f6f6c147e9a21987aafe28cca951bcd026ee3a78a3e1778bbe39ad14f716b4471b76fabb5c835ff0b8a8cf918542d0404dc4bc33debbe5c7290237768f01868121fd680641aa8308726107403f280d79151c8c8e8373343f6f753a8821785419d0535d6e98ca0aef307d1d72de5ae67e30d51f48e21be9dc81026507ad3e2108cdc1c60e8260e80ed46204b26011926d09a93a2d73df4b5db63a348b47a32bfbc2cb5dc6b92c36e9369cc54713d69facf343a36e09c64ee7c971610e110ab351a48c98f3ee9da3efc37308244c72c3832560500d3ff39c0848021d996ad574c24851a520f2581dfd85b7e4075a30aa7c0aef9bf063aa88b69f96bd31d40e98d3c4b48351ab44c1ac05c3a21b354c3ead882daf263c39569ef9c296a71caf4205e4623b274b41de3a06c786c6f8be8b64fb79f4bf03a12f920ac090f67d76ef2e2e659e589aa1698bf57fd50e2bd9c94c9696eaae997ce7a6d2c86337a29f7ad1aa1d31dc8278435263b857b876802d43ab922dc9f6f5a0ba534aed7d61db2d962acae5144b00c87fd804f4040bb00ab5e98c114dfc7c263381c6f46941bb5e205dbc505455a3b09e8db064ce154caa175bb6f4587512340aea0f0dcbcdf4aabcd338ec6c00cdd7c6cbf66d9377e85670fd3b7c9f793f82c33858996b041e1e82c6ff7a965ea8c7abda848399637cd0708a0ec1575bc7f45d00ba00c1fbe77ff31a4b8ecda405e51a1c284f55e239c02a08c2090140c2f3ef1703740f5e733526e043cbf497ccb7b10643bc2f1dfb63f737e3280dcf88310a3736e6d927538096fa21e75a92f8a04ede4719170c9ae7a3c6b3e823fb0a1fc71328c4000b70a616396982c9c1430d4794efceef6842878e22e98b5c12ad0980bdc9b025687d8d77267939ac4ea8f31af20130ffb01d4bbd068bdbdf5d65280374e53caee4329dda4888ce7e7060bc677f9e7a0abd7de0332dff3f4739bac3a97ba856a727a91b512facd836e0dd37690c4e19d0b577c4d24822aaac7fcb1533cfcf174d800c915279e3b659b8466b476884de12af25b804c4ad1eb529f2d6f6e4fc9fdcf02e86e76e886fccaadb6ecc96f2581596d4ca81e0cd920dcbc50cc0f6e16cb5b7938b061946e6094a2cd407f69cf6c97b0a7c9847e49fc339c22a7780da7510b13907ff6c0533ba6f90d09db5f6490170ea7bee06b174652abf70583de1962774e08046522d8088fcb69b965136fd83c57f60585d98bd42496cf9eedcaae189b682e1a5e6d4feb9e6391cdb1b203e96e12ea6309a99b23bd2a0a0577e897c09814878ca37e769723d2c5ccde9239c8b9adf7bda80cfade9c52d10b71b7773c00b6085d55c39ad234236f1a021f313143e51476bb8a158a5496807e6d2ae37b9eee3cc971bb542ef7769221ad78a505a90cea63194f17aacfa6a2c6028a3efeb3aca345c12e70b551ccb7b6e49714d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h65cceb6c923db940e156d95f704c4f5e0922f00b2a352896a3548c286ea1ae9b39bfd0c39628135831fddba3d3fb53f903257ba5ef4803d59ba28ba7a067b5a98de5c46c78b09996337fa17f3caa19ab7e3b600f491252f10b83279fe94b0bddb6e1c6e7a3bd5d19cea81d7dc3678d7cb1042b0ab4616ba90bbc6648f77ed666d2f46509375f404de9806ab988980ba0f1626a9cec3ba6920d44653dbbbeee308b512e2b55b1d14945a9157cd07249a14668ae5c7bcedcd136b51a8de74ef9bc37f9c2a83c72c3ff5d01efb4c61708b6c8dcf93758b4e8fa08f6bea70d2c47673762223a41c68de8fcc9670f9e0fbfc1ee0c6749d4b48010a54f46faa41e9de96d1b0af82aab2db7b1f3b17cb1260f59f3855b323eadce4d820d4c7a3df261ae6a6636110883b94ee21076d2fac1ea80a3fb79778690e592529309db81bd18e50d7ead06c261bd63dcda658d66957751da3b1bcd61fc877b72cddcd759b9f648fc52a170c333e18c263e1dcbdb5830f3802b40280fe016309c5d5701fe852d965a7b01b3b277914f787736b6f87b60b9f0a29c18862c7135c588200b66545a388d90dc0bfd99164ef66218dd3e521be7df5f965fd5436d76606dd9a424f345c75039ecf09ea4f7d4b156b18f2372a0d60d8bfb61f2e0993d29036f5946cefbd2bbfda4c41d59cf81a0f07532fd78acce05a553573c1a65582d1ef32d658522faa1b34dd3bb5fcc655b7b64b14012a2f4b954cacd8b03a647acdb029ae1b7ac39eaa10ed95c2c26f738a908c1b9660a3034bc2f9aa549c567109cdf7704185625871c9e792851584a5c42fa5c4076a7cb577e79689c8711495ef806e0e8abe4de3f4b3277d66c9909f43ba21326801f189b3d7ee1e47c1a2e30d322d7da1290616e1566e1770b497811b3784763469e28dbb6daf93969cafbc51fb75c95c9e7c127bd272cd38de9ead4006efbf91d47dfdb2bd638cf20782812025551977e86c014926e8b3a543f2aed6db1efbcd3cf50b5a71ff13e496865f13e54870511cc2685d51c295c89c11e467953b2ca3385e0bd8e3cebafdf5e4ee9e0fed8cabc9b40d5864dbf6522984094bad08d7bba53f81c2eab58cb5ac2714fba830a1da9e8c8872a128ff4a8bd5dc2ac40e52cb8b051b05898d5d461ba71533d3ec0b2317c6a8e6c6f65c631b02d3ba7eb745ce78296c527085119249667241f23123f953322690d1bdc4ecf87a24135cdc4f8965a7c6214cef93f16eb334220eaaf288d00be3e5de3fa39979b044a40ce8b7ea5662d7f6629ea5f6a27b905e770833ca43a8207e879ea84f553a74f0ee6842646add3167c9a946626ec3227e53a4df8e01974f9659beface4e18fcab44e23022f13efc4acef9332e1f6736cca117d1098d255db97462d4ff00a744d42e2ee55b8ba4315da09ec51b252f7a56ca43a3f6b726abbd0b900a71d720546f364037eb0d7b2dfdad6d63feb2ff2329d1f00187506206034158d36082e5be8ebf57c6935ba0534369811ced27f0dbbaf78a46add6e9b86c894b46a20df1715e5164121de18d2e6efb08a774a3124046fd9d34e23dcf1935e85dde6a8e254177f4f5aa77a7ea60179ae33ef4f25403007df59ffba1d5de9fffc9725af695c1cd8a1cf277082d84882ec3bbbe4f52baada6ab7b1d77f8b282ce797d80f25b13c5317f139516f5059a9899ba399d3a57691d8022ff64a8c1637202ac0bea6cdd43a0d6832cc32e4cbb049e9143159d0e8e808cef05cb965ade62911cd1c6fd1a5f4e7dce3b1a80bb60dfe55ad0e760b287b92314b64a4091a747b0df4c2895a1d5442b77995eabde859a28fb7dc5806c528d73c54aae371e59ca049a0e35e7ac16dd990907f6ad46a8c2112e7867f61cc59df54e29fadc19140dd463d8b4a0fd57324e17397e15cf5f90d885f35d780419e90e0bfbc3a6ae74b263ea20e76c07bc9cc3bbc5d54daafe017927c6008760fb0b86bba5e6ed632774ba1d7081760da4da25edb69d83967d323fa15a9afa7009160d65ac15abb8bdda5dee1f3e64c2587fb6b1c33a4f2a4a81f5e8ab41681172ed80f1c520f99b584eb9dc0b936c6903ecf45605e6c363023f0a857a85996771c1976b07b688ec4a11e12f61a4b54e65265e7fc04754ca56ba3a8432dba84d806ce52cd2ab984952fdc025a4126fd5446f81ab2be854341d9982cfd76acc5e005fce91a83d4b3a8680b6ef2a9c88abf3a0877a05b8a6ebd918a1486659e6641ef230c812cb8c42c8cfa7395729ddcfba8009435769cdd1605765bc0236e17c1ed5db0166efcb00beb9f80287778b4e80c5d476ff99c144b41922ab764713624ede53f7b0eca28e4df2db1533a10f584d4ec5f35967dfc601c6872f0fe7241dd3edfcd105d74ec4f4bb7722598df14ea065dc92607ae5a0c0802bc0af5dc9f48270aec17f31851d407023ff40eae0a13bab5b9218ae777596a68b97cedfbcb0b00ceb4757d4e627979daef4e35a65801793b28abd997eea270a8576a59f4c71aadd3b118196b41b6d0c9d55b6e824e475aeff21f327780b2229e323683e17015fa831ac244191f9a20b87a025a20b7f01de2244864509fff908690b6bcbacf0c712b9ca86ea5be724cc4a042512e72c3c111e6163d00654b133fe52af45eab5f0de5e570e2441b4205592369b5f61fb9b27eecc28c6e1f34426705bd52e73a4f7ad3a150bd7d7a04b517bcc27fc8112f3a59cdecaa27d8ea87e65cf25aceae079e264bd23c8938f606d6c2f06afcd125863b0a46cc3996e96028e2f61de9e2fd9d140830939d1e9d25aad07e9b425415e22284204c5a2eeb053bd194b86c909f4eaf7fd5b8ec3e79bfcaf5b6a1f9d631c98520cd2e1f9d4f2482f5e74307098d5391040333d86ab351f811850170f3cdab3210f03365d6f973235637f41f7703beb1fc2449c9db8db3707d61beb9c9aac33e0f8c4820e2064c5fe66af432f51e805fefbb0e92ddbd56d676dea2d986a4801b2c08440df910dc7aeaa02b89ed7a6ad241cb006d098efb9bcfdf7830abb56668b912c94f0fc6c476e0d512b1a8b6010b96b6a5f53b6daf0ee9fd82e80823fafce9a5fb0963dd084499d1f727b05e05991e771f81eecacbcd2d674c2c0d0be390e2c926a2510304afc39294a7e0663f3b48ab7899473ca61e2605149fbe53b39b9830a7359c7c47e68d0ce67d0da948b367d3bb69ce0c3f6291d33593faa49107161231dcd9667846c1617dd7112d09c5350dcc1c160fa0aa6fed6a683e22d49feaa27426fad8e966e4ebcbe84f478f95c2834db52ce9018ea0ba5e31d424ca129a6c814cbd46d7977c155cf3902de47d3899bf5fa55c80d6a7ff98977395757bc54d36f49c0dc2d4f6ec8e5c7ebad92d9a70db4c27b7f6ab2effe110cd5a16ddc404f4553507dd0089614ffbb543f138e7a79c1f1cf54df1b096b46641a7296f86515c3f0e7341574ca4f81c7cc1f6e535eff20dc6c335e97cbf8cd8d777c2fdcdd14c608d895cfb8910811034f254212b10ea6b1fbf9b801eaa120245e9132fb887e2253b89c37ef415954aab665ee97fc99c2dbb8aa24b88c5f3f520d7faaf98cc79c84d1f686eabc2d3e5d4576e8eb4c7964b95cb8de175fe411955d57da5d01b65a73d5011eeedb6a7445401833102441388f375b287351a189e1ebfc1edea8e20adff4e54138d86b6bee6f3ea61642370f29b9121c7bdb5c1fec1270dbf13cf4184b0054339e9505cae7d2d856e40476f7bb59e655f7910cfddffbd6fe92d19357b99e4df946c0542fc3d37721be0942e8a7fd93c6f6a66c1b3b40fa8d88e68d188d5a9ebafd37888b0ea31995b27d7f93d58544e82fb6a063dddf15eb063537372bc49d1c74cc43dd7208c1e94a8406efcfd5201a48cf09f00117b1849655c1cd6dca3df6910ebee0f6d51f44b13cf362054210939eeda40aea9e3b289414516c8b50c08b2338fd72dcf6e12f25c44cc583cc9c9258effb7a3b185fe99feb72fcca92eda3a7da10280b7da7c681011501a522f2e9ce792cbdd385aaa432c622e24fd09b3e9cfd6d0a6dede91aa1d4b6da431f941dcd5a14cc8e7efe07849b1ca6ba4219668d7803c45d8e2f66de34ebfd0e7bbe6124aafdfce6e1100263188eaa16723377aad548bce07f6b1a633203da213d255fe83c8409abfcdc30879a449701efcbba27d06342db8a3d592b6fc732e71542ca6623d70fb1d2a32c9230f28dcb5361b56510c861d23f8a73204db1e1bed6355112cc0104053b9a2ebfee53e187aee55f5daca9e260d81edd5d474af39351d1080d5fad81838426dcac153f0788ca036341e590315b1f2f5ad6f61ecf7567f78db311da57588bf77aa138cb8d0e1a1e92b4c99bc61f6bd964af9db415213e13a140ff3bd67d9d440e05451d832a5fdabf39a2299dc28fd11210ac0b872ac99061c13d3dabb83c7b147ddf27ba00289a7b8c3b26510fcff9dfff32ea04a4c849428560bffca76d43acb51ef0551a93d9ea9146a5119b7898e9ab292c018fd39d508ace507bb965900458ce3119c23dff9cb65e752ec97faae2bf4258cad1c563119925abc68a84507ac8264877466f5ee4484de7bada834c3a6a887e2f2f77c2667e0da2518b28b7df9f76faf0a3a58535e88bfe553c68511da1194119638f32a154b97cb112a0de6bd5e698e41ac597fb5f150a207b648a7e0ca783332da0236df1ac4bfb9e61fa78ccd8c14564f7630af33aa11d585dbfb6b8f365f771825c399d702b4bf9c9c72e5892cf5c64b9e0e35add35d3821cab0814c13fcfe2fb3d038c3e32812dd8d8b3c234c3b76e6a47165bf33a4f4de56e829b9468d951dbc8552fd303108d03629d68f0fcdebbc440ba101c0891b957cef2a1d5e2a6ca0e349e47d8e4b89b1b177acd965b06c49b782c1a045a00780598368863da5401347c8ef4996e7e58b92b2a8088674a10316e7ccbe7ecc9fec04446df60bb71660f2af8954c3c53cff3bcc008408edcb87d31569533a14a3cf49634766c5f33825e762b81ee63eacc96c24cd54274c239f2a08cbd1a8e40443216e7f7a20b37d5a0481833e520f409c8b5af8d713c92623069799fc8e6debe41ea9436e504eb4b838ed3aac7650ad2c7f9c9ea4bf7e89c83bc8abccc5835f376d9e1574a2cf2456c31073be8108d8369289a01e2507c5f64e6d411d339c8fbad2ac7ba84856c5de3800d68eb25507dcb30c9555e3177708986921c9b74af24360b764c47808811d67cc119ef7046cd0cfc63dfa49fff0f4b78aae2a5d731ecce1372be85d69b6e3aad53d2823a736609b953a07075057ddcd1c68d36783277dde49928e4c21c2807be6c388e33b5c029a757200da6fece85086096f38d50165ff3636cefc361fe0fccfcdb361dc476beaa8ea33abe512a9ad8a8f7c8f76ffaf59ad53dd4d0db105199a6d163a92d8375096553d09b20b412df71bdb4e62ec79acb86fc1602dae79264770ba04595a0b7793cc11a15186d8736908086247aad6801f94bacc2f192f84aebd5267af861850596000493e5f3f2d3ffd06e66af7f84c77fc48921e56fc7684d5d24ac9313bd735a532b0936a4b9334878827883240e7ca04d8937fac17281ea149bc50c7a8c211348d85554937e1638606729acbaed7a8185b1a2fa17d96a662f13f780266f36fc9647e07ee932c1f0dcd0a7c2df292413f1593b790cdeee0bddb33a1757a18e45ff06b33060c39fd50bf4c3eacb7e8ec74e6ad9509a33767cf36c6ca7fe85429a8869f6762f2a489e93f8f1fc5b8b2b9c5c9ebcca147;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h13a1df9257836bbecb912b1cd2bac0341cff309c783939ef887560c303d9efcb7e46fcb85a8f177b7015363e7192cdb9272743bc622d31a9892119a321af27e12dcb2cd6f0a3eb52a263020f3abfd58f4dcb91750f71230f8ff4fd6e6041fbe507aabbae8f31e5b3ab2e5942017f463035d7ad32090d355766ce1a2ffe10ccc02d2e757c137e15489e35afe34a11df9bca530d6bfd5b356046c84c68f2650125af77e157dce8b865af2ed21b41444ce6c4bede98b345cd898bfb86a98024c2386dea7bef575831a0a7aa4b7ce32332cf4350afc96f4d908081771b41bb8cc666e7d4d57a930113ee09eda6287323bf5e515e7da36f4e26df7e525851945e60bc3ce902fcc6ea196d1104e369ba2cadfdc620313c9123b5bac3405df3ef2134a99ab1ffad29f2a7fcb53c522eb183e40e8b7686079b2f94969a46911df20160e1e8527519c1d1e1862dfef97eb007e84c28cf54e21682e6a38a4d303114250fd3b52fbbc8021d165deec239d2ab9ad175cd36abf60f46f8d849a649828061cc80ff98642527d396f039d2a2c716294b5be718999c8ebefebc1730bdd797ff32ddc137fcb6eaa7f86a2aaf54263adef15f551a3f5b668b4744894f7d3c962871cf7af74c43a77f355e509304eb64624d3346b5bba264ec76f3d0e63c5e89d471f51098288bba95cdbfef3adc7c5fbb8cb5c167d34444af2dcad5016b9d134e074b29cc0f1b8f13108b26bec1a133b0b51b2b82e08e9defe47a002ef6c132434e4e936c8d15829e17e86e54f76b8af2142bb9904acd8d55707679ea92393a9b982681bc9795722632391886d011727579dddec7a9992e33fee355030bc4a9f5e588fe67d1d3937518fe65b21f9e3cc992a5b9b0a2d61632a98a304c2273f4fb2e1421fb8222b9e4574dc6083aba15f577feb61a3f51674c48ee037e1fe2cdafd7a12ecb643a701ced1bb645319617181ff9f7abe29e74e33f3974c8ec3d4384a47008e9e17062c18cc63effee012d851a114b4baa33e129a3f8790350a7c1c1de8394e1a61143ed5bbe4ea9a5eb757ad71db274000f082f0159c16f4eca3b10038d4d2b56ecd4782b2b760b66b9ad50b9fa785bb46cc685d12cf9e3446d3250ac96d768a89675e5f7d675cba4bb8eb804b2cb83a159330e642a4f70ea49cf77654ba5c03356d06c5da15bd16088a8744d261dd331d7cf2d654f8e0017afffc431d887678fd17610ab943301c30f83add0cb6b343c215642c5a5bc2ee6a634faffc9f4b0cf36ee38097684031cc5fde6cc2b796749e46546cbc7cb7b45d7edce697753786e4535e83eaf2db27392202f1c436e0daf9af2b2d2e1fbf60072c1282336a9fba296881da115124aa15f0370d0d7878e21134b3090f11656acaf80d9a01d77b22aca68149b2478a1b6ee99e8cc091c690118bba24d82f85b17c51783d90c8346818cb288d377d3c91a32d64f78c710fe07713d6f77cbe54b2f1f566e11140d9b857871fb76230723966a1caedc26c16cff960571443fe9ef44f395e824633c00cd74e96ba071243619ef32435ab19f791d5c6b0a04b01bdb846df7d8e1d67e4c041167f96622d8cc3c77b12d1a52a43e607bccbbeac8a82149b08f7bd96561ffae1a5fb5c74666389b9fa22d53fd989a29a0e8100232e6bd9265959a8a84f8f2ebbd04be954af8210bf1ef4171172efb3175dbd4337ceff0900491d76ce1aacf9d75cc3804aa6a31bf074a59c4e29ad26a6e4a5202bcc1a6fa5993f83f9c1a5d7ccecab3c9b54114623c8d099e7d5c40d7d08ddee5349272c3a6136228ededfa20c683d5e66dbeb82021024433fbb7cc78d6f7430994c96922560df31d9c2fb86a7b0eae5a86350ebe1177fe8dec753602f50eda8bba96219fb2e6b102537b0387bcec0828bb4b6befe047a0a4df19dc758c1e452ef30ba504fe166d05291f85b3825492745d59af8bff5ce28871be36806f8e6b3be0892a303d541786e59ad112efb8d56395121ffd2a13c3d24e78af79472e04f12c811323bd8393445fbfb3d96ff08422a9f14e8f03f2f17a1dfcbeb679ab7219bacafd2a7b499b2593850ce813e7622b216240bdf4546dfc42ab6fa52199db993c4c8f3abd01fb590bfce283c017cdf4d748f1d4ba961d67aec6f2e26e866067301c3dc2ee839a3e01f6c4bb4f08e90eec35fde98447a5db92fceeb0b300fe9d24a9542e5c806131f8897a2a19bd9edb13196cd181876531216f19257b1c6818a1716200e7716c1ec25a781eedad12ff777df84935826c6560a7ebc374ad393ab8c5ff57baf876d2bcbe45ed66159f8cf0e766946e62b635830f6659695b9282215acfdc18358c1b5cf1fd54d2003029f615aefdd6692ea6abe00b23e60477107574fa753194146fe60791e905688cf37ef5ed59cf406c5ab32ecc59973ab4e50c99ce9b22f57ca32b0b5a5c37eb0f501c2e30414b59822cca48d40e1787822494cae6012f3bcd39d139b3864fa64b51f75e9f88e03b0ec5ec66e743db7d88a19557d4f71775652838f701e2b82c8522749d9bdc4c2f9af154709999e23d99598b9c04c8eb89d137cabdaf6df0a620fdcd9ba6bb9f4c5d4f7d851828b08fd1d62cfb4f848b40b61bc22d1ef87fcd6dfe82ab30aa56f023f2bf791f16586f71c850f9b5a787f80427964fcefe1afb2d9bcf4640b9de1d9d2cde41ec5f78a66b6b88953f75d057ff9f9e77765645b215f875457a2c9f1fee4f809fd95bc837c4313e869d8d16497a6f1c255bc6b017936f06431cec814e9f9d3a61dafb069e1a3896bd8bb60e44888ffd9c4188a61deb8de4aa1c5bafefed7c3ba713e481ae88afd4e982cafbecfbd11fe6175dfc0187a88ad4237852b8cfed031effe24e7e998dab246fe304830f7a3bbfa93b47a6656ce04f951aa78cac4ca60980099f8b051735464b99d00b2e9dca2f29f327a6a81a667f849f9caef09f7dfe6e2530025e26199a09c4da0793e90d444decc4ece5de79db535b4f7206a8c56fbdaec6420c2693b2bb5d53b957016333f4b9c9b107340c09c8f6b6a0621fe69a5823653e394efca540fead57ea58d4fc1e84ddc7544471952068d6a428a18b5f36e83f415d90de7f459dedf68e1f68a4803f6e7cfd0327a999698ba14631739994afe584c6865c7486812b6aa563f7ffaf0534d4b2b76b60a33541d2401124d53b2dfadac06194daa52f1374dbafee84a3c1f737cc70d4ecbf1bbfc7ccc3908ca198aca7d4f448cac0e083a0e2ab23303cfbb5171a42824daf27c6e59e7fb92cc08a3e403e1d8d3549c34cedf8e95d266151a6dfd09361c92edf201a68fb6c22c3c5e22f8ad3f6df1def7e9861d18fff34cebc4c11d0301418016a7a4c257b3090717c9860ea4c2b43a4685fda4e37790a8b716db9833c0f22d2f7d3ac75fb035083789d8417bc853950b65b31fcaaeed6ee63f31de633301a10a52506aa9f8b859f3213a4f8d23b43ba76daa4f3a9b341d112f478b0ef08679df5a1cd8c81cff092f3f67bb842166f8df575450693f46a0d5d5f16880ab1b65b5840d4f8fa42d8d0c385732bd8cca63cbcc5273e8b79165755a919d02b9dafab4e95757dddf224d60e383265ed8549f6dc6d9ddf3918a640af94d9de62e1ecc6ce98df69fdc8026c6b3871606b5eb55159efb14b914e8a09ca1cca45f4b0204bf1dd12e593cf5fd6c472652d0b0e405b0a26608c5e378c71d0978b3e9fc1e7d45c83fd458def2e68887467120449543ffb75203d467cbd6f186cfe32cbbb4fb23fc39747b93341011ad358302ef960eb6c4476ccf4ef06f6a86f240201b7eda442895b3ebe93c354522b1843c76e719f9fd91672fb7444bba59a58ecfc1f4bad8e4a95ffbaf0afc378dd721012093054aac1ec6d9a76a3e198c12394f5fe4ed6eb02030c2cb32457ae16dfb53b727cf1af1244820edc6eb11fa30b56017484488cb369be4648ad618f00564b56c7a84b2d112cacaa23a879a90be56fab84cac4c870e8a4ddabb142d9a8e4a1dd1690d7e29ad7aa5f80a1969d085a48c64daf60abeb93d979e33eabbee096925115b633507b44e68363af2da9214629ac2848ee29a3adef9f9b6bddd6b4b8bed0ec9703c510ca55e2414e32b65d7fbbdc151f3ff01554c491fa0b2bb6a288638f549edfca55579346fb6c9a2f2550538fe875c576875d4d2ce8eac5fea3c6e04c2744e66bc262d443c65e50e69d6c73d820c851f8babbd5c67ff2b4090f93bf0d7d035a2a884d57bf1afe0df90a864466f3de21f87fa753c219deef7366778b197065758481c115ae0a0e84a270153bb4e81fd6b2f3bda1444c71d47bc01bb7f3c0d6b77c1f64999f301a67002033c3ebb0fe6f0270f14b078987c1dd6ff9643f83cac19595a4fd3d80bb8ecc4e0daa24f84d9fec0e2e9da38127ee2b9d9fb3183cb9b18c013e23017a2d4bf3d0dcd8e3238f0c65a4249c67ef32f3b9192d19d992b6528dc128be2b9d78fa0f1356bb2c06e08c391c47d54ad1e3718f139c769f9b205a6f32481362f47c386e1b06cd426850c4ff51899f70e4584a1dd78aa811684edc9b26feb5a2a271196549b1b477ba36c7dc995c7a0ddcbdf8c2fec31975211913aefa798e936b32406e8ffd47cb8da5f72b5dc4ac50a29333ee3f34024ee97d0133501d5b4e2afd70a921a2c4395e31ea977ed12ebcce27348a56b17938991acfe4325fa69c6baf0a49a3cac6e275ac9db0c81b53175cfb897056dcc7a2f01e1749b8c3246d2389a2870ec9bad152579002add966fe874ef6c8c88c68c0551e5ffdf2efe679262b5f73fd58c106959ca4178c19479260e8d2b2d12c5941cb30bdba990979b39402f24668c1227cb84201238901af2d4f2bbbb25545a17c8f63e6955add221a046efd1201922de6f45acf552061ba44633f7474f40b7cece075ea4566335820d6e78b7cf9e53bd1609385fcdcabccec727ddce965dc23a3e64f52c99633d5c0708a1366bec480af0945a01a23979f6f8f0f3f2f721ace593c19b7150d3d725ae7df822cf496fd528fca46b1169ab582b4d1a99e7f6fe5f729bf389fe8cf81daa7eaed2643deca4df7a9ca1f548797e66ac46526b67f6a6c5f1e2c2051a2741f82c1bdea9527dcdb1fd3bdf8156eaac201ef51ed929b4bb61586f8012dab503b9dcca2c8e728541374adcb43921c651ba41a902292391682f586795f84d3c026304cb81d0adbb44b4d6f59e4cb83b4a4810d8aff4d955506d005968d5b27f05f4a707d14ece5070ff18a19e200362f5475922cceb03812e7f1f022237cf8a7f1dd4a431408438c949ce030bc70e88ef5758f9cc37f43a06d8f7acb8863dee4968d0f5884df6a48c5eac6690edbfe332305e84fefe3cb534836bb5d262ea9aad7b6e9a5619abdd643c08fd20275a75137de5901b17a2df462fd628074adef9a6ab54dd1db276947e619a356721e3a45db3ff6c6154da2d508de8655e51b61e9cb8f0c8cab9dcd6d320b4ee227b5500da6379b12e7c7414ba5737ef85661999ffee086686e7eb95c7131a3febadcf2f5301c2951ad34ef2be376ccbd000666e6f25a916b919d4fd249e3811c51f0bde3bee7a84dd7ddc9701380fa5e8d844a1ff00140fe93d287b5d2d23fb9df170671252eb9c54f1ca6cf23330a35c48cf530ed54567884d65102a39af8109dec119bfe46942e4a88c48d9a4d5057dc875728077a9e9ebe1b4594c363d3df5d82c83d23e892a217d8b2be4e9815321d526c1fe2b1e11e1cea3c9c025f07b46cd9e5e415b46c8a625a4e03e17b2b3e8171d2061f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb45baaa73f29c3904ba78dff388c310bfc1137dc7cf6e472ab31c1364f830768b6407f141f5dd68e3c24b280e804b973ae5e1bed9748ab9e2f6636a601ebcca8ee77f5ef36fdd47d292f7503e48bad712f263c4c99df3a665e6db3c1622db5b910270b6bb90cc8fca51bce2be59dcdd58850f46d6f7b0ebe5a25deb66053d74bdf67c73b999b86e07409fae7fdf632127e3075a4abb28b2b9f24cb89451b2ad877467d1d6358ab88c38f6007b888f1803149ecb01b2fbdec0b3b728b22e173062f4c7fa0eb3fc338a6c0b951362a22ed1dbae9e97873dc58dff8d32e0a71616fb26da71227dcacc8ce5259a5097ce4aa2700c5640b109c3bd4eece347562d3e454773e3d24010d36567c53dfa372c5ce040bf09d950ba60a3b0fbdeb154162373ecf74dcae8205dabe9de7c62dbd0cdc3aefec8aeeeffca658908d60ddabe56e6eb623c548054021d029f8ac8368a353cb3ce5dbc49ddbc59fe7efcefa7f0efa5a5f41bd9b42adfe8efbf15bf0e6c21c16065d63710e0280881d06fc8a26b116a58432f5833c93f08c3508ad91a3b2c6847b1a80fc7f0708f493f77fa5164b69c75ee8f23105109c67269c6f01231168939446415cec7d11c1ee5d03f0ffa9993154fc56c0df3e275c6153d38a4710fdf427f90dbbba7303ab5618953a3ff10de94be66f5a18f1dd3165e3433fbe2a494cbd229029901a1da576e9fe7d63a80145f76ad7bcaa71ad71e934fca465792f7525d8c55cdf4086ff5bfb081529cf72bb4111c05e487e74e490c5c5fcb85bc79e14fab867e7012519284ab0bb1907a71ed323eafb719f78fafd0a9b7949adec85739d9089e9f37519b090141e4e1cc8867d95f412c0292c19161bcf6b671ef8433aefd0e6dc8919810d089fbd1603771a7f9f4b4ea43e9c2c3d14c6bcdfb8e85e64e0632e4e614547d225e9b1515a6c111af845112998dad0983771525426f2d0515a91fed0e61a29a3d2a56e71cbf8f2830f70eb4e2b27526970526cf32851d30dd398783a72ab70f13342f5a0bd46b7c2c52d2741b9eb8a427108f71b08efd51f966880fc61fc5c07e14e4f9e0b37fd63e7544beb47405881e6e0f69cbc52eb49e44290c2e347e7b2d2058a15720b2105ed436c8aaccdb3be11c1febf816ef25427621a5f4745bbbf8cf53cb5ffd9f3a9cc1afcb0963c4e4d7a903102ec17f980c0437589e30292a59cde00e7e7bb154b64d7e58922be0ad93702d55eae7563dbf19ad66139ecd604abe36fc72c396a8e67ea03a61ac0266dc674866491b8dccd2bda73820f66b149e55220c399a0f158542056f20665c341da57ac06401505417cb8ab0b9435182ee4f06c8f08766fd66212f60f52ecddbe5f32d14dc74fc085f60616d01ab0d1bccd7bf727702606e8f97652cc70083fd019080a343d5ab84bf185216c5fc9add4021d3c83ec17e6991aeea51c4d67d0578b14b471f40e712f8800c2b51abb40ab194c3d4315c7c8cb735f4bf3d0f93c4009e0b9e374bd9ba08330f920a48b811e60047daaf48b061a540f979885666d715f6afbc3f916d2cf38088b4a019b4fba5cf51c631d1d923f3fe2985d466f0ab707eb359aa9036873b405497b06eb9c2dfbf98e535c646ed1f69d9e1d322ecef87599c47e5c8a6733896a40fb0eb708d7cb794743916839b100b9a915f754e042d752643750f359fa82d1f8fcde531fd52893ab86aa33d1b588a374b00ae83a1ee69df6f69bd8b0b43a2ab9c62efc4d11d18b85cd3283c491966756a8e4440ca9bb92866926e3e4841e05610707acb2db653753ad4f2ada00841db822edbfb2c7eabcb8123b8b28ff87340183862c34d5c6cf9bd5e0ddae27468e84b67ada18dcf3ebdcbd42f852a5d15fc1cea32bc2a969db0491c6a5fbb4e372ae5395b2e7db03c5a4a5a4b8eae1a900e7368299cb8663f7a128786923394e875c7dba7b2b08bf135c2808c250778b838771c56dc636140e67e8661bb3e83a125543421614806edfcfffad7172b6bbb273f3b8decfd54e1f1792db97c83342d9adc882e4aba89940045669e5b94f60a3b3290b57aebae3baed2c9ad3bd8b5a7cd814cf2403a8d6cc02980aa91bda6d0575323ee468d153ecfbf89315bc95555c806aeb1e35e939ac8cd854d249e4e446eaab7db8d7f19b882475a09f01e30374c89e2758987716b215f828e41825f1d2dac09a3f13c97a9c4cc8dfad5324fdc3423f5b6bf989244565ad14082256f0211c7291babc03ca35360d88f51b807bfa3bc9a8f1cc040433a1a6209133ed7cb58cd3c053b11856e202dc019419037ff1f564d50a3219a17237c20d5870b5d6be29cf0a04fd962f06ad4b3b8408e6ef8296552179cc304a0f623812ae1defa489ee2f7290cc0dc93e1125570e2e704089bf0e12e1a878704b7f54aedfcd6be9bfafa69105850a4bd53616318fe58a875307e4420f84fdcd7d7211941a5ca781573b36411cd243c160a2749d56f62e44ba108b55687039ec08638c0854a7193417df1cb6c4b5d16e651c15ce18a2cda4dda153d8859ec466a200b145a72f717d8609e1f1657cc1eeacc3e8c0467efbf19838ba9bc9337004171a9dbd1412545e16a1aaf0c91e0563a0b74c60680025e6ac3f42d12487b305a7a3b2fb9fdd151b616e2a239aaacc0b3b40051209d21d195913733c186a2f0fca581ff8a1203a997661e678dab0cd1a1a0dea99c2f11d6f49c4ce1d01af07927d592aa91bf4b1174bae8a7f9995680c6270de74e587ca25654a1ba1d7aa08679bea960a36892f0a176e6ebb32dc8f112fe83618a917628fdb7c45a234977e066ecdc3621262218a670cdd1f138e8dd3e19ac20e482a199901f2f5740efaefed72dac9ea2adf0046b8d0e016c6cc07e7f05dad5e7f433a98bea333123db8cda484fff9f6d978ef71767038cd42c7d7f9e52cec5b4e5cc739b66bbe4f0ddd5fb3c2c4ff9f7e79b33e3423c9b93da26f051d572ac50b018023f96418311158270be593e778f37da683f53a788641218a7fe541a2b152a68c6fc459c5f80967a1d9f1148c87830d6f735c7461f2e6f976a3d0f51e09489abb67da3836777ae9f10a3179bc10bf4e9d9b330d26a0e628bfe00b4daac07fa003d069565f097a1da6db189cca0702d7d7fdd92489be6753475a016e5718af77cc850965bbd20b909f11e8ca58632149c20c65e8d7be3402f946f7551aac3caff4380dd4e2b8ef8801748380ae8188ca3775447a1c243fe842793cb6e346eb51c6b947470716f25f9f27c21c75e748ab4b9667420a996a351466b89a0de45def5f2d4d27ebc2b3fce8333a372bffd45a18a4f7951e62ed7360d3ee05ddeb4f4516e2e343b11ccc7eaf8434cda88acfccde21e8b2feff6f5153737e24c9610a03857b187cc2063ea6041d7e26677e6284c654dbb4a20c697ecd050ab6eedc09e9137c1e946217e385fd2d85f2987da9e7ce9a61dfdeed3165e3054f07b55d80a9ba7d935a20f6a1f65104f665679375cd00e3aa85e6fa0e75b50aa511fd98cd5a0b84e43be8e44886a3e57907a97bfbcdc1ac838535720b642f6e15ec1bbbb494dd4dd42a107678cae8f829c75cdc89e4309ec82392bcc49ca6062441e96334789323fd728294b98a883b2c868bdc65b970ddf532648f486195a578873112b53b553717bc1135fa6e6e193c79dc3eeb81ac64ba9099e7185f36ad71b44c8e7267d039efce18b8f21d95e5e53658d7690edd68e34aadec3266dc096be641a710a851e68a958d12accb1e0f9755b3e379781169d988d7c2bfcb18c557960830bbe9c998ea83ce8cb0591caebff3c5577406f2797c4a13b3d407cf9e8a4ed6a46dbdab78b45bc108ebf6a7a93543c7265991f011d0d9c1493cfa5c573383d69c9fdc718ebdbe92d736f9602c65fd227e06ff0a5e6a482b146b0520d3902fa71c595851323f637ec14448d7710d2260ae5e4bf1d5c89455bc94dfe33ad7ccaee5a399436e0d33a25c2c3c57ac8ad6a75c61a0cc927181320a7f47863ac96fee68dcd4b76739dfb1a5fcf9e892a04194b5235f771561e557bfcd0b7358eb5a11f220eae27651d34587097aa8f48364dc33481ce4bd19bf57a40ca981f5807306d4b7b068565f3c6dbbf46b73386de9ffd135f45563fe6935e670a64a04ab7573176b8492d167ee15df3a210bd7a556c99efcceb1c7765b53089c68ec5d1c4b47e43b07c9d26bedf607aa1327c611d4f0f3011c741b3f77af532127c112bc1e75edd566e2111ae87183549948a5eadda07b960d0b4e990a5e90868920436c039d2cb5ea786633182fc872a8fd0ac558c4cefadf094d55b7d31dc38f851e6f5595fbd4876205e46a86bd3896f4d0e30723e3144b7c55a1a7eceb82dc11028c1162ebd4af9bbfa0967608ad91cda158193150673abaa8f9a767120d77bd5e470365224559aa2a24dbc912ffd63ab47effe8a8301299db9f98c5c3d07cbd3f02765f9f5743caf83b83117a2642b9ec0a654bbd350a6298e3db5962d8429d8c8abdd1123771cf061414bf21f0140adf1182cb94c37bc147cbc60475c849eff0dc4ef132567fc442a15333bb019bc74576e6b244cc965d056785a084bc8249d32787ebada29ad6e1b7deb31f1aa80e15127f1f57697223664c064484144c145db38f1de045650faa44fb9090734b9a8bd8886c14e1471d8d01319b273f87c6aa9d1ea9fee45af361732880950554441ddef7b4423de23c84bf465619fc1f5fcbccf3acec0e67a89c719d7d7db01b9d0581997c973ccc4729256c48f574524bc1b6864c92171b082da52c89e3d5f871e7f4df185d7fcfd768b5a587903d5b1e9ce3c2fcb5a7a0a5830f54b651e48b75eea418e8b51de7f9b8493d22fc56c11244f9f00e9a383f0d21c71b030cc82c133e2c4a8b31fcff13e363e8780aade7e9413429432f16f0bcf73bc37164f0190b8c2c099823b9e90dc868797e4eeb9471f81928afab19619c47e97dd5f301da4dfcc7be1bcfb4895a7e54ea83fdce769c38bb9a943fd84d151e76eaf5af0fd8c7e5b04365662106c4e0b04c36e8d2d75e96e535cf0cb6b32bc086d0bdf5183ef8c0f67e0bf717b82ee6849f21e30aaf1570dc378e909b93ba06ee7b96e9140c0a722a0f1544df231770ce936c084f388b272d239d2969b1d4393c2c4bce458e400a891bdab7c2a5f120731a2ef6c452a0b573b6bdfc06d3f507eeba9e9a3c2e7fd8fd9c5da6595c69e1f0b8a9b2db511914bbc4c530b9ba8603838c7ca3957bfb5fbbb43299e4d779311908e90bc67015d256ac9c036092b42ded6a96f629a5d88f0cda4dd8d66d07dc60c95fc2a81c633b929766f7508fac162c3d5305031316b380f0b09a913df452b616745b21733af1fd0f4c2abdb4aa328f5566896be0b1ae31bb4a08d889b1f4ba5492421f1d23a9d44936418f053691b9af6f653ea4b5661cbb73da4b55b5e4a40cba983e11e1caaa03f2463b2869f640eae1cdebb62717527bd1beef25bc9961e302cda0b1aa73e2c2348765d9f3921bce0007bd05867b94d035dd1dc575ecacc57c1c0a8d77743a55083846507240d241ee9be9a31ba5cb135d85c6901254e079f4c506f3b4cb62ee9d99d1660c57ed27aaf0064a72695754b85939beee4e9852d3040b81a902c372e2853d5263834498e77d852d656bf0f42b5803059b28e513bd36f1c379022e0e836734c6fe5676680844c3537d3d17faa4b8577b70f92b6505e64e4c7ce27764a4fde426713580dfcfe553bf495216c770fb51ef1191d6a34034deee39f8d3f898bb30;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h548f15fdf6993fa328dad3ca41b01705939acbe4400177f7a1c6f7b166df1c6046f065067acd646bf6edd81fb294c84dabef503161a84d8f9e6f976e84cfd18d34578790a68c00f6e50572e8f95e95feef72c405a1ed2ac99b72030a3b0e9319ec1b23f5ba565b37bbb74f952de05a1cedba3c07bb7476dd19296cec514c12fdc63b51bb3bde7cb3f46c8c6452bf7a99571816f6a7d6519af9e0419075786d7a719ab25f00e4e171efaf79c2a80f5a403ba2fa5f71ce918c926129b85b17ff4b4f52118523753e864941f3af46daf5bd02fbdceb5d6da906a014e0c2a7c3a205fc8c65553e1559d98c5509736037791fb45924da1f2358f8fbb9d83ec71a4b122e09fdaab7a67fa8a9be9df9fa6fb1807401fa6838d481494dfa4360af0c4852016bc8b78589b7b04db301f18bf9463b19ae5fd4bae2bda8d48db38b406bf68ada613987ac9196754bab1b0d396bdb7e43dce7ffacb2eb445346d010161919628697b29bb4014ac1ab145f43898792a7c42b3dff70518df576fa677001fdafdced7abb01d3188f5c4b5a1ddfc752498ca98cb6de619624a209794a0f2735b19eeacbed6370711b1fea2f49a5212b51bfbf295787d9d26b3244517c6dc58b19db527547ec5aa05ab3210641bdf08d0bfcd1c4062307222ae405184384c8f3aa586c6372f56d1c9cb21682a8d6f6f23a4cd4ac39aa945e616e758621fa0189ae48444afef33e4a7f40fb9e35de3c796e3c7945835194cc781de8d2c8a0c0255e5347239bc39c5c89f81e73727ded1454cb40d83cbea5bce10cad3a2874bc3cfe9b6edecc0f36b4ad3866d15eec9a7cf3fc4f6420a7679ab7e132fd419121e4da3c2e1fd4b356ff17685e187c5afcc49a3ba322007e80366e7c5f9659b767d5c895b434ff7b2c751591e3a34c65680db3bca6a95cd4c121a33328656d376ab67dec35d2117f9e6b764dc69aab8d901cf6e508a4a9b4543f851900c2fe77c3a9dfff5aeaa9515defaa44464e49e9f12af507d48b02314acddac4d7f1669f1d8caafe85d3ea33c28e260fec6a551e28ac05c6465125edc26d4ecef950c195a58b2289cf6c2a48a096615c6e42db67be3f320972c3d6c5363d64322a5d602b9240883e2b437b86d0ac416c3ce9d59ad81c4ca5ce33bfcc7efc879bc7a364c264647035e6f3a2d7ad78680f1aac7150ebc2632feccfe65449e1b3a9e95f0ef9335d579090e70416bf2c642ae4232b3db0fc3a97ecdd79ce242313eca31c387f9fe26af27935db0692980338a7ebf9676d16178d4939f7cd6919bd316a789dee1c6674bb2b24ce6a7a6b964ef8e2bd74655fb3576349cd85d9fa2bc4535312c83618156651e477e8aed1df661cfe67141e177bafe293fb527be64f99226f989f87e5ffe9ef9253c21315992a81a36b51260eb6e781266f3b4e7ffb3965e87dc514afc279d59be7465c0ebc66a565a4f88e96aeb0969330ffebae7f26f0ea868835f9a38dd2fd5579fa55b9b9fa8d13eaba21f1c015a561685ba603ec32978cd8140f69363190cc93e4507fae13d2655c432bad2e030c2d29c75ea0a2f63b7132628a895ce280c1af8d1811f57add1187634ceae992870ddfb2cd496c203ac31cdf0ad26bb206d54f4b2250062079eeb1f4b0511b224ba130e4763b963bf64a80af93862349a5ca4237e2d1d6e7327949fa752adf0f4e6f6a1a628314c305dd60cfd38d02ab35dd5e30507a9c2c5400ac85c3514f8c47fa5fee48f6e9881693baad4d66c00d3285be71ff59557f967c9dae7b1c939073207a94cf53cb91d57562363319a1f925812d66ee8526980358dc5b5b92d7872a60e63722b97b8c394ce20be703c8436c438024bbaa9bb96e41bda566982cbd6b77c5cca7fc977536d47626caa0df42e3bcf54a2b1ef4c203c4294c591c3152b1763cdd2763f426df21569d409c8fa6142211496f209a4811e4802cc6e40d8410e1b554305bba2e3a2014296c65a4614adc021e07cb8a9b896d756e9f35f290300711278968b90a02f2a25be11dd6906c6c100ab6493a34fd2e64f1b62298c1d7f7c56840745f58904af65069eea353c0c1f0ff7e4994e92b878cd0a9e8df47788e9de29b2a6feabf027e4f80f3a71d0eaaf0a3faf6917e7f76a5abbdbab2d17287efe4dd13bc1af494511b872425c078de9a70e3e45a78aba7325d4b86f3f0d9bcdd9eaebf54fad77f34544c9d2d72dc9b067947e1d3b222b7cada8ac0165f97698148952fa8ba3c7505632f70a3a3779c5810b1e3550bc83c2db409169f8af79ddbc99d63d5f7c673620962fb82b327953b84308123ebac22263d01d1aa5afd24f8174afa1da03bbbd274a0df30ee454ef47ad8eb820a0a5999a0f66dc56744687422655dbc4deb027461f6e19b4ff23728abccfcc5f3db9446bdf2a7f982118598c1996f20cc6fb416b2d87c50bf1c396f0b6ed7ff7cdd5ec083108324066c51409ed401a9c42c904a75455e5e642b41887adb4bc0bb34cc389b5f50e91b7d83de2faffe032b72489469bc99ebc7ca413892ea2fe4dac8bb373d1f35a113267e1835e980e632e2d819915d5a229da3054a93db18ab29a386d39a2b13ea3cedb82c7e6b09ebe499c15cba7cdd4c05d70928a941135a01b788ef5fb00a1453cb45deaf2745fb26bd7aaf74786a2d21ef920baaed51a97de892bfd34fc8cb75c2d2bb9f49b7cca07cf8b35b2142970f17dd8b395741fc2802e7e1031e2e6106115a3dc1d8faba3aa80304732fbd96a45098fb7591612c8df92193812f55267f6e6d87a5d606c6c332b65059aac35f8ae065868eda61a6703e808fe66c4176d10928787c422db668446562cf461184b32171b03f4969131f629f8415aadb884246a15973f010a558b8f71fa902531750bafb7ff0a6efd7e5aacac02df1cc08e3a34a8045d2e0bc326adaae140722d981a5cf9d2b960b63f5a8197f5795ba55fe716302b0aa02b0cdd5f98f30b4c9eaf393c965738709325dd96a80cf0c7030d26f84c4d353b4c552c46d0a167921898879b26d3d08a08cf2ff5ee70a9720b3e05285cb9630bc9d8573950c96005825c22bb961423c34af7c4e8c8f7ff5e9cd69f69e37ddb0d81ddb96c98b3ce8742150c96f6a0105f6d5067d5924e60d6f2c25cbcb1e3f497184b078a106ad163faccc7ca7fea526d154429d91288cd2802e33c9345b447a69732322695df7d84d4c19084f4799087bd3fb750c1eeaee50cb4f3d786befef8df9f4286c82a4572b9fb7070ce3e9a062358c19368d6278c805c1da3ee8637335bf4f96d4bcc7d0c15d34c69e78ccc12194c4a099e23836e1094a2ba70e21bee5043245aa971a8d361eb9bf677a4edee010ae9c462d156f036f02201b5a793c1770ecfba2a274751ccf7d5d1ac67d680db2fc9cad67cd1f149350627a94ae3d6584edb7a33580c079c01618343ce815e86d0bd02278196db4191912f1e8d97c8890cf732c65b99b2de5979b9c96ed3f3c88c978dc71829f1c7007e724426140a01e51048b2788a3e8db2e4f16a28d63de6f94d4f75a57c2ac64649edfd735b262d0c911ad64299637921a0dcaf5c17e1285068216376d839f71625d352ee2a722c3b7a45ff1d5200ae171519ae0d4d51207fbc39aae15d4c657d6f7a03dcfde118003b92d1af54961f60c6e769077ba8e9087b0d95a82d1a0c944bbd759bdf6ff5466888ea43959549ddc9bb8efc80b092510d36d28cacbfb4b5220e7c10f123328000e297e13d0667b2970d2f259d22aef656d39fb53b165900825182bb10f6884cda923fde23c866529866e0bcfb880730d3113844c8d88e91adb5bb630daf858ea70b280e4ab7a22f389429da35ff6938e5ab61d6dea910148f19e5515198d3a012e2a7e0c04a5c542ea353b6fe2b13deae37fb10e21453c00db2e8ab85e36fd123b028aea0a8224e82bddd2fe0a034a59d0855e0e62cd67433c18eb4ee920d6c38b784c113f7b1a25aec0de7ba516e081b37aeef3c049b155b1d83466e189d419b2784c51d5dc65ea1a3d6899b2212277ebcda72f406855db1bb859e5d22768c31d92050c43ca89e2568c812237bf8aa356958de85a403358fb1b04857ef7189aa8880af9ebf21fe36c5424354df4f8b80c0e2014d9b5b82573792c8cbde07b27db703297960eb96a088619245af37c85270d1431d09fe4562355c02ff7f9f4cc7ffc4134d6d3ab708d525790b33063ed96a3653d568928fe243f2d60adabdda06f23e632ee9dda0932362ef627682a7b7cae950731ec2a7e3b2613dbd117a5f6fef47dca1c48af23399a2156abe3ef5a72a3afe0a7c7cb001d7aac542cff43d2262cba25e38d74fa355325a85e404c4d7c49e73001f8d9d4fee1094735e498d649d1d581b6ffa22c21fb2766a2496ea95856a2acbeaca0679b4bc4489bff7d26bd985754bb52f814daab6145ae9a3b9a68a5397df8a55277c2350d7de77da7c98a8b7b90d6b1117923802a5d334b64a803b87265389e6eba6066c29c2f94816023fab1c982fb579cc06288e7822a7718ba5a3f6207566677a57e82e60c4d51783a347bd547dfab83833b1832ed2fb7fe385451030facc175a6d81dbae3e86aece00939c76a4824a393d8f8db178e568b183a1cc4a056033ff8d42cac7e40bd048d5afbd518075e3220bfe8d9c3ae06f0424660a18e107b891bfe1f0e05d0e2493c425bd3d204c1e4325e97a8e34905431820912dd9f75f201d292e44d1c0d3f8828d6ae20f075c22c11471651c9736d0bd8eeaba79aceb5eb311424a6eb7bd7954cc99562aaade2c62a28f0f8d6ad5b7045d02d9fb9333deac6eab59ab201e16f6e8ca010b714d37e4b2318dbfc855862756ed84b6ad413cffe53efd85538f2f256a0d91b68afce93663cbaab5e54f08184f6bba1e950799c562c4eb966de4d108002c8ee81805cbb9d709b784dae69638fbda7a89a87a80aa4d7967128ed70719155d91a89c56576a67bf9c187b07eb3ee9bc3cdf7437fb7417f15c27daa75cd20ee754616ffe49b5eba2f8033baf99a1c688284468a9174c72e289b7b45e0b587106143fe76cf3a29a009e7b9264a7923f40f14ab02e17490fd5b8723aaf07225361688395b1184141b263c08df2d1d613b1e0eecb7a9e1f32710a96e1edc0afcf2dd2299b75f6af8eae192d2960835155071208587177e6869e3780158c28ec98df3de93214300a1ea0c518edaa358db10930950db0c3fed0b739a8befaa2c12e36980f4ff4b237a0876009ce0ac192b0a78c4f992af339949b00427d5405415f4f3b2b875cac91c9358d7597ae8439268a33d16c43434d2f5ed082cc15a5b8f44f91ed7665c522d33588505276bb5cd8a33db8bbfe51008abaa6069af12469682a9a3f2daf651f08c588ecc0c7910a8e8658060e91785efa9760c0bbb627594bc646630f65a7408141a79fe2564347de6538ef6abf74d0e75e9fd1cd1ef304bc70fa62ee9ae4b68a66a8feb9289f115a3f66c55cebdb49bad3eefc8e7b20debc4f763375bf4ef6c4aed30cf94309ec8240fa468b6e3050e97cbf5a6bafe8103d7ad6927acf68ddb508c736be244c05f1433411a3b171dc13cff6d7a2aecc438edf1bfc608446fbcabf4457381a9c1d2d088f9e0d91bd92c0e955aa00b71001204a79b8994e5000e6e2c53e6cee37148f16fd096a7ad8bb1323e5ca79c52283cdb8ee3282b40dc51c53b1e0e2d6dd7c3946c33f24a5b2feaff47d4e934b784612a83ab8785560567e4b871eb5debba87c9acea7da5c6e4d480edff869fbd1c6019125fb52;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6021570dd2f87efe69b37c9d6085a17c1e9ffc4e3222f7c539328619c9d32ea38c848b35dc12bb70325f384db01c361a93e2137c10069921decae319e1a05f01a6d936871f477a66e738196b106fe57c51b3a7f1f540a8126666be63d572114b9df23d537ed439755119b422a1f6df4663175bd095bfe016876c7d4f94515437fc540bd48fb8a8e0695a2bd36156ceabd6f8913fbe5d8a6e1a8ed23b387fbb962db47600582bdc3748ac9b475fec4a83d2e7f09ee1142072aa17081a0466db7eef42381dd04a56bf390792317d08397c59519a946d2391915360573f7ba0d684de2a2e1cb5913819c84f98673b2aee73495da5ebb15c1e90f85093799d8a92a0a28036079c9f50bfbc14ca67baef286d1ac247ca915356cbb8d42ee121d7935d622c6ac3a890385dab9433731d5de26a6a0009b343aa75eda591bddd1c9a60126d6ddd93fe92f40451c8972675adc56bc2f93e9e47461ee628311afef16c2ad068abc87ac5a503b0829cbc52fb7bb2dc85ef363444963468f17f540fa659eccd628dfbcfbf4f65c5a4a2d5a160e19c172929d301d63afa1c446fcbd2141949381a26fa68a16af7aa7c8bdd26d3aca372aa1d9af739d267e3e5a6a550e4f4bd669f0b94fc33c95c898857e729c0e81dc953dcae635e11c52a13e620dbbfb5e351eae8b9097d09a295fe945bedf6469ffdc4fbf02515c40d7d95f9bb3b56980c84783947e78015b72d94e6c98e169d0ef5c8d7b1dc62782ed034f6e4833f5cb05e9abc33dea4af47543de126f4ccca826d361e79abc391208131de094642d1998f9cb5d92361702fd31e267875eab7a24d39f76ff77696594b327720fea0da24e397e0080cdc51212e9c88e60ba7252b54ab12b892978db9239709dabb7f8ce7f55053ef31c0ef7b1eda00a5458478048d94f2bd8dcb8e2765ce1af52786a65796df17b3575f75cb64298dc932b781119d2d1d6aec21f357baf65961f3271c161701c1a1a32d7f38265e272aa1caaf48a2925a9b44614810093ddda27c2eabe68fdd82ac18309cb00dc32d4fec5eedb360e3f2cf7c685754f9bbaf2b4917747404166213302efa171217fe066d052badb5aba4e37c99b5cdd0a938977ba35202a6721ad0a2c490b82506d961342e4e605b84882cd8b3c685a4bd6b253c41d06735ba6ebf6be14ee6e055939ccb636ded9f9a1318298d87e296b9d1a10f480a7c35957dbd3f9baf9342170b506b7ed7d397fb0fee1f3d970c6364afe098ccee65315e37a9a7cce4edca8a4bf1d305cab79ef8672b64ef174490610268dec3a1fa823c4d252bcc99f129382fc6ee536ab6d20f6ba61bf2d6d15a70b5b711d735a69413e597b1e1c2cbc04402c2b783e4bca39879eea5ad89c1ef8c206e114cb089f1714c3279638c040adc8d55022c6301993393f77329ba55f01ab9232ea1c6f38a12b51b81ce5e4ae875051aced82fd698fd8d4dc367a94e1e3d52b9db38a901c3fe426abb0d1a6ca92dfc8f23039ba389d112bb79113b6954ac31f80676a8432966f244167d37f00e02074cf6ba0515820ee2891b53bb19e66b0ad9378921b66582596b95a32c73ac741e3da03ecb6d5b63f478ed9aa482591c13aa448d2ab146311fb962aff674744f6ff39fbfccc56678795be1f9f47226a06182b449e7ad2f7c6e4c22f9086f5a496668e581e2f7fd8cf077ef7d8264da2cf0ed0f65f955c7a8067205ec70f98e4a3bbfad2126577e4a1a218ff700aa3418ef90087fcd090362d06792dbe921647f67a2672eed4d6e294a224587972f9a8c0c5a5470f0af5fe3e632f7b4acd6b5f6b31853ba81e633fec1c8e136dde169421ee81eb43722efca64841397c52fea24382665c34a5a49c8f68a11b9195fa3b56861630ab2c86db0e75c91aac36a45acf4bb4512e1607edd5333febbe58f911dfd7c8c81ca491c9508dc77e7a278717491611cf3f2269d0e93a05beda7db4193784d60ade1670aeaeff7c0a3e1322ec688b984672bc38a95c3c9549569dbae16a234fd33f86bbb71333319a863910b92de31cd62d610ebf592896cfc87dcb39caf31115932ce07a9049af3ea4e4648a8b12bb0a967664b8d10ff0d1b88c2aa044b4b5d56ec840bf815aa5c8f4b992d18daf64d372b6add8c31870d0764544228ae33e00cd3577e0bac3d9a0e3cbd9b0c744e00afaa6717ef6ca85a660de118d0cc48c7ef68a54ca2239d0e2f39f82535994e9292a0f2135c3204001dd94f9240911f3599411e4f496fd936f2fb9c807bafb44d636314d56550fe7af6fc4a9e50a1250fed5708ad8d4fc8b5bfcc5340c72e8d467d0b234a3c40938675757f565cd38c31ba78fb28dc07a9e33853667d84f578a41aa6a70369741da4758a1b91abfd42af23c3c67d97d1d10075e8b88dc62e4b70b5da30f48c69d966bf782503b03718f66e0621e64d611cc638a312c685901841152036729c18e6e88a8654cdbbf7eeb91170e3c51786d8cd4d38334cfe300178d0f8cc87e538ce9a860598e4072a6a09324ca7381b7b8b0bad9bd575ac68696944df3c9b78009b8e9558a1c5454916dc489ed3a34d2dd11d23b5a92520e50f7dba21611cb1defc358af4f8e31fa56564af22b500c9975c4e458f065268ebff519d9e8627876ce4da58b6fe8579846e43059cbeb58d8785efafeeb5c44c324d25dd81947704eea15e37261d1a3ffb31a1df7c5422f75bee35936738e841fbc3e8a6641d563f5ccc381e1bffcbab8d198c7868f6799d38fee756aa7579c2bb9d68971e1e1d69de3f08b9e4635c07b7c225d146ca0f647d6798773e2dfb903b27b18f5ac753131d23af4cb8b9592b96bee9511bddcbfc0df6cc4df31dbfb361a8706915f42041c65f99acbba3899a5ba7b9c108f585f99d77b72699406c0e4f2037ec10a5b95a5ab7fe350616f9fa9a846cbb26500347a7229bad567ce467d941a59579133c20fe3ba957fd1cadc88dcba218782f3b172a7197c69e699533bfb502524bf06527b9c92fe95a9740cb777f7d106d810d2317b5d375ea50e30bea05c37101d471dd49101108764d1d721942d1fda24b0024ea4c1c26e7dffe19e63fc3e51869aa031b3dabcd20f90646b99e5b92b9557cdd8b16478b4f26a3795468203ed794d10e348dc86c404a0ad14f169bb7767ae657262fa073a15168795d874240257071a2397e0f62e712bd8f48ae8b689f4fbef0d09706b4c53b74c3e2141b37d54802bfc54b69fd805c94e42be7e58e5cb2830953aa96b95c40e947371d43d140fc2c8d2d05951c2cc02df11d76a4b8dce85c3bb9ac6b35420bbae06a6e69bbe12980ea52bd1c580c3066deb2c1b5392b3c5077a7c727e9474935d9abe059432c7c66cdbb0bd1cbcb48356e7a77762fca4bd3added871a638c6e65f0bbe3166549df4f77e2aef11f917f1234e5d7aa27e949bd1c187c8035d851c65f1b630ecddeaf92c6b5cfa776bbfcdb1ae7abdda0b5c0a0c02341d73623169e2b3ddee1351a7d8631018c89b0e2601ed13cfe9de9ccee70cb604575f08848a036ab3cea7392a5a4be82282cfaf9ecdf6efa75e15776a76290268abdc345774f0b3ff6e8ef0501580de5466b7baf8591a6fb527241287409a054418986f9acab8f50cc1bfc15e6310251a58fe90b9919d4ffaad916caf07621971a905da67104af6efd8510aac8d70621aa131de2c20b480687872a1e68dbe5576c97ca541d87ce82ed85b384b8cde4d0437566cf3e7bae61c134ceecead91d1cde61f19bd2a4fad7d8e3b38f8148b14b0ffeafe1a95bdc71351dab08d30926ffe06c93568bd8d48c056b62c7551171c3f60922ff6199c93bd33bf2c2235d1d5543d60d285bd6bfaf80c657d81adc291dd60d37d3196d17b7e41ad4892251c6e80d5e5dab196bcc06ed71d33d314b418cc4af5a456701213572dc3753247a32d6c0d2040e448cd443f4de11f6ec12efef238e9bf5eab412674f5aeae00c7ff5a8497bf73c58f97f569098a68c33ab59c5c454df875a65b10923c10492c992b2796c77849b1069b0b1d6845b0122701b1fe78510e9acc61a579a03901412cf00ce69e586ce5b5176f2da484a5a5faa067a13af6f02d8a0155746d25643c3f9ff7535611d502b7173e719cfabefacdc8e4bbc6476403d369d6913341dd470647a0e94aeda7c053076eaddb59842807b2cc6004ef85a805e29ebabc6577f878fb8b49a1af84203203d826c014edf668bc3635f0ede721deb2310e84364e4053b3c0d2e8d5ccd274708ceb2d39900cae52ffde9a8ee6afe35ce731dfafa9d9a770e95b550174edf3ed88f73a9daf9c245bc9045c6a1e03d27b032c0f5bc96a4b3d44794ffb2df9a348d0fff84eeeaadc2d95998a2421bc30072b52964f54e59253d8a81262cf83568b740671e62cce213b041b317da674b31cbc852aa6cb9e02021711cd5a249a35f84d0c4f16e2aaf6de2b770bf86c1e0e58d43622e4f2346e25ecc402e2391ee47c0c115a3aa80dc244b3137af4587d3283a65b16886fa3a7463e0932967a380d9542990cfe010dd4df44aab8557f0eae0cf16bfec2906dd6d563af33fab82cf657f1d353923652e15bffbce38e42b30628d579a62e580400d7ccd2d8203ce34c7280dd6c37961b5466e78d386e558b8354d3deb4de2455d6e8b946c79f0b4b6f4ac37cc561b46e57d3f532ea713fdacd8c33bcd739b381f82274efa6868d9d250b5068550130e13780c842842edccf565fe6f57faeb6b31f10b2795762750905d4a878fbc67434734ea83e1fdccbfbe09573973c6683bcac31a32081c4304c299365241d506bc4e8b3c3d577bbdabd49ef24e807caa05171adb5a5e47768032db6a8ce321fd99bf73dd3c87d943ab70768cac4560fca6fe2dbe86a98cac6df0e724edf704e6214cb896d5acffa8fba6ee911432db8b4eec5b81abc0d2fd37f82545aa62bc126098ed8ecb4d2a3ab099ba101b2086ff74c28bc35caac8fbc7df9bf09703a134972d5b2fbe985e75eae7cb5dbc228721cb0658b3f44fc4e1a1be62d0d8a1ed54a3494fe40012bb271d0e0783e9cf6a658935a317c541ab0ec83a9cfbda670bdec83a6faabf4a543e5b81464b75a34db187d9876a95c26b83b7e8f08e464a66a1f0229eb57c014949805217950b696fbc592d2791ae11681084ca9f59525495f1ed02c031e57954b87715a126e28821cc41687fc751312e508341f915d1b4cfe2636e45a966a6ba4ceb7a310b9be86ec3d3168d740e2f78502902a462027a64005e73f424ca7d608e27cfef78257727d55e27bb51b76ef944d7aeee0aa8b2e765a5ee907264e7bd2e37a98fa0611a1defe60fac31eadb378d3f056d191bb3afbd053e1d7c0b6942dfcf83f24938a19ad5c9a8bb9e97c4766a377594e6f332e1a5028283fd573fe844e1be0307918243bd4ffd48b171d3e2b9c258d9dedefc4be0a3ee49c830a879fe12d87003ff106b58d96e7576ade59c7dda5fdef1e5bc81f20099f0a111a43f2eb51a93b1714afbbc8a77deda04b783d5c91d61baf042c3837f2802b932094d69d024b161655e9dbefacb2122f052fcc5ace2881887cff33d271c3228b410968ea8a86aecd2c50ab8b095d620993d83bad404e68b3c2cbf3fd6c2f71c638ed2c41e2dfc3dbe06325ce118252c104aff9d06a0e5443a9fea7b9fb76e34a3487c2742b8eef27cfc56aae9fc68f786325fc05eb94c771cd99bbd436f49c493a9f13cc67f8cc7177a731beab7b8046c7ccfb8be91c75a328d68531bd55c83354a26afbfb8df2d9a1215e21ff7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc8e3c4ebcdb30b80f64db37f74d8d0156a0d16420bde6b21a811ca819d0bdd4a3e3370510171f04c8992406f3203c70f04f1154f384a2b9513de4b6f3c17599857f59f1c6b810a0b9248308d2ef2b30886d28cc900479ec0e82caa8cc44f4384eb49f8f84b8e2cf605488dec4507e6743f113010fdb22a294bd88848c8a3ad3964c95f50cd6dbdf49d27954ed07655ae351564cb857932e78de0ef6936a29a039603efb199223fa4fa99d4fdaba4500507ad9278b7ed61d62c222e7833d6bd39884d2fef6ae5ee1a42aed928a321c784435e1b72b2d7cce188af45f753ff20e1d53466d14293192505c8cf4945a5e3078b5787244f92b734276a8075bf0ae18662463fa918cf4661d19c586602bdb1e378bd3b1bf5683a715ab42f2b4a6fcc84290961e1ecde945155c6d6f37db18270beac26a6a320f962e20edc8cc005742be0da2cd5965ccd5a026ec5ef6f0fa8417d748339acd1f49ce19e5877b60edb78ad2ad605bc3a8d240b431ca2ceb3111d552de154c5f4e00d64638003d775016abd10193904abe0bcc4553082c676a634115f3a738b80f724edaee96afe444ed5c071fd1c3e85428bdc212696de6d201ea16557b54e0d1004505d56e5bdbf99c00c04ee19bc336603f0f521404f20ead5b96307a250404c753c19d4ede69ddfca6382c69086665170ec49d1e94b383484ba46826f26806dfc533094e9c829d4516be1e233dfb9ff7fe45771f508bc7cca2baebc6b5e8c4d21de2e21debc8b5ee1393641a1f716e607615672c381eb4a55d051e84b1a1178fb37c510d63593bfdcee4afe6cb76c42ed0eb4984e4dc50660f8bbd24883aa1c1f1c8a088eb6eae954d24459ba153aab3dbd0c87925ff2018445f37dc679e2738ca8d88e2be631cced0c61735800bb4b12eff51389da3a614c95bd6c458f0b23bb764827eb7afbf75a5bb6174ae6eaa10af1e9e232f2512bc3d3dee902b611f9bc21506187ed4114d6eaa424f1e29db0be393e43292b2cb4e714655ae6caf92b9fb18946a06125eb4fdfd944459af4c1a871604b3632d30ead5f1dddaec465a0ae95d21ba4f7a7e4cb9acccc918019c9f1e6c35e80662175f3624940ef52e6f871d41648d2c77e455ee69923c66466b453f9d4c610ed25fcb93b14718f540ef961a49ddc5214a7a5f45fc3c7c48bf1dc8aa5db7cacc0e27abcf65dd5cf1b5fffd3bf8632c583d78e70c9383fc2cc8ad95b0344937e111fd1bf056ba57a890e1fcaf0b2f89b5dfb8365b8c9ffc5d6dc63195f636bd71f6eb3b5e83c08c393121b88df60f6654d40ac8859eb500b006e11b5616872b4e6fa8a94458c0acc37bab25867e5f535f7246a9ae20fdfa2cc44fc5d837180e53dcc195e4511d3038ede92e303292a8c39ba90f2c149c351701a089d4f30e27f345339477b3908fc72c86a80c2cb83969b023eb71999cfe23b52015a0f0f4281d59713850582bc91eda2beaddd1482e2e07a9555b9ac9a4754152735a7208b3b0bf807564f2045b135cb2107b2394cda8f1bd2a34e3fce57a7237ffc8eea65d99327fd3a29e35314b8514151f5f896c65b041d374a2b58a6ac281b7e0e68a66e60e3fe8d9372ed1b3b84fc63baf9d98044f9fe378cd1e3fd2fd4da988232d5409a95987bd51a970543ef0b01086a24a7458309789c9f19750f364f58f745a8b87e2ff46b53f282fbf4d2769839d297eb16f134ef4fda86d74ed0c7a10f544babdd03a32aab8d68845c8c2eb9c89426766879277f526a16a96f52d2630ea6b69a53ce5012bca5ded205eab4823a86bee102e2107e876e1aae0c1a4427693c411a0fb56ec77c6799f5abc4fee5f326215f7d05f903fc299b323faa44e6371e03e91aabf216edbdf63f5b554dbbd2f58581c89fe1ea16070d8c7c69c037f960671b1a7f2d35c35a1e791418f0d70545bdee8778a6dd37be9da4b03b94e7258c8f55adf0966b3c4b78f50f6ce3bc0de3ab0e12b3e51b9c35605eec3508d67f46a6f995cdaa4669eaa3c656706d4fa94250e286635deffacbfb81c0b981699e52db49871ffa33eee5bf6f9ab3e826b7b8faa25e98eb06c85db190d5ecbd092f52841e6b4ca914bd4c6d019fedc0f1c6e4d936e67db11682017fa740808bded0151315b8afaf4a5cf4b1cd058b61d48859772d7ef1a200edbf00523438ebab2e721cd3933cb49ccf322acbca7cd0faabd49f63b1d5c6bfff2f5849a3ef62f5998591db64b9634f90ceb215f07b411724ea240394ea06ca8694d4e9a01392b249fdfef8a2bbde42c5d717b0bc870923bccbddb58d27c1bb9594f2ce938f98044187450b717fbc77b4a0725ddc64128eb738b50857cb114ecefde13372d2e83f0a7747a686fbf46c03780c3e26f51093c696b3a1bd0bf9897d3f5cf581588c8dd55bbd3aa26a074f6784f0c4d5187db4adad976c468281afe6b24cb77680f049adc2a95b2ceb8bd7d0035deaeaa6e27c66f35b3b837c954989028e2841450d760c1481e97b3912cefa5ab6e503a801db91b403a0386b56a8f6371936e9c2973af02edda7e8957dbd58a5d28bbc10f3175f1d749c8c247d4db85eee9d7452e45958236f55410ecd65d3652dae6402303ef6ff1f974fdcf36d583fdd7a0a2f15c3ae4e81ee0b9d8f9d20bde198ba7a0bb799fad6c4058362a0df7c4b9b736f1b59cbd4616498758e019fc2462815e906e3ed3c9802e3bfc3d5e2c05e3411dab9c91a8da589e1c77a31e4b921104422bd71811b72c35aa79ecb7e3b8d1eed63d38d265072c840edc3415c06f45d301a1de19dc375117b9d6425bdc65d14a8d9c4b09fb2344072be28718533226a403e812ce4b1a33b79f50a5542fc1458398eeda13a52bec19373d5b56cbaa75baa8b297d9c6af969156d3e078c1d06bae0429733d3f907f6188beafb2757564d9d1a69e212874708186937fc78ce82f8c9193487ab2d0c7445e361ef2a8f5ee9024fd637578a21da71d3c25d7abeb0f8e5daa6cd7547031aef93b84cd7af7ec131cac5a84cdf0f734cf355144ca8865084ea5e5d2bed3172268be82b3cf87ac329137ef0987be648d367315f7b15d24246f5798ce60a0b7a04c7b3833b41debab1c7ca0771c6bffaac5ec3bd38deb611e60fada9c184b3a25db5c8f6d54dd8fb466b8a63d1480ec8b03146c4f5ec7a543c6b743d224639768f32bff8fbca70cf7f911309668dbdab3d06cc8479ef6b728d73d222799f6a2d111de1d86cd559ef77323b8b301b21c8f899875a609da987f58e320d8e551c2d89e980ccf46ae163741c908370671dd8cd74b8474c95df9030bfcd1957c8fd232a8228cff66007b9d1d07ebe3267f165367d02cc83ccd394103bf29d92e7cee614a267ed34f6510daa3c34356ddefe89e1a0d1d00e322f5d1b75a704c3f0408c7d25ef7601270ba8f9bf19fa6ebc93df7d6b787e7d8991df33b5e6472d00df2c541fc7cdeb6c8a8e0861d1f4b9e2d29a3d1e8484d7c15372b9fa34406498676df21b767c1f4e22181a6ec41284f912320261dff1401e244797288518128de48c91c0b851ac6b34470ce6297c00d5c3f9b5b2a49129f285906a8998d8669df7b3c2ba966f7a8939ee7775ccf4284e24482b7bfb46077d0c06d470d71881f5f718ccd756654b9d78d19692560eb3af0a226ccd0ec10b2b929793ca3a78c35c2974ead056737534865d71e6658bdc383bbb8f2903ddaf07746e953c88cb8866f9a38dbc887754e82882ea5f67d5b3cb7d513698e88700c08e1abd18ea8840c1fe53fc5e087acb6560332fc5ceeb4583d53ecdb873e2054072ddbb2ec2d5ceb64ac479d1ae4059853a9194b1416f6796b322b417eed689d1e0f84430517edaac6c8a550078b0ed2e6a79c0c920248e4cdc02a5e5f834760b48a0be4cbb65288c3753e8b30be68aa5cac9d0f24d9bd5e1b287c9cff1f5aef8b87c43d0493aaa40209648235b26d22eb69d6ed2610139b64644fa7f360c356a911dc0ff236246346cbd670cb95be10afb67b63b5dc0b90c61d38ee7fa649459b026f16de1cef74c0aa38ac0d190eb220cd1ccb9b55a321352d23fd86ad9de45e0f767e5b1ff07d8cd9b45e7c33496995d4ddec58cabadcebf26636fb0b0273f733bcc4f3561b32e3baabd51d697df4aaac64944117d40d727ed44464d66b55121070840185b727b56c9f97879bf4c44cadf3191ab73cc2b4b2e7d563a1a5a00121d8fe1cd5288bf06571062570b13c4c96e8282de4fb6bf035a01d5761b155a4e8d901b9473ae3af0a1d3eeb187d34b3a3199fe19c94bb912d2450b21f32c55c6af78a34e9112119d42958b7c0ef6465d72b530b574a31343b274a4485b388357fb9dedd43b402971b71066a64669740f7809b41b5ba181159c53fd866b980e340591dd57b967633fcc4da0d0f63fc588f1d1dc09071a4e8bdc50be241a47dc0e000c246538e7edad538a46e642e745ee34dd5b472a755198fbaccb7dad2f5e847aeb72decc93af5924de7a29876e7a29767b57591f2db90cedfba83c91aaedaf820ee5d662ad1499136e2de810dc36438b126e6a436bca5db8c864edbd4cc903f26403e6e11f196978139eab5e5e4949762938266a0739a07d69bdf61d44754833b916c87923624cb4d174f82251225b3e1c66ce12bff3bf261af53fc4c4f93172e48c281ebef2abd3339913ed1f12afa455d1df5f3e5fdb68dc2bac2a67adaed3d686c7ac28a099af3eff1db1b1558d1f1da3e7fc706ead480df9eb756679b49956d7aa08520022788dc02bc642301069340ca778454cc93df773fa83a7ff05e7cd6c087079630132240858120f185dd80ae3e04b29e4e5e1c1eeb6c6899a6a55c27304aeb6be6eb8ea017dea6bbcb06927b57ee58d08900d949a2a11fbff6b9b73e4654b65cbc7dd28974a2bad41a1f188b8b9a606b271244b415cfd8e060a86adcde5270e85371cbb35fc5cd302a72d22b80e987aa3b112b8edf932e675c56fd6b1545b7d1b751e22fc70997e018339daa8fecff5c3025e5a03e93f0b9cab2c3cb21a9617fee36d6b371b29a3f9e7cdda209abea0bfa43c7f21cf457566a57d89bdccef036c67132028d2823f9f1931b3b2c69973a82bbf4441a61b67e180fa232def9d85d7f16b12c1fa86bf0e59aec25d7abe7ad527368ec06b113483614b8a3d3c5f47347bb1a3372e06bd70f3ac212d53a04cfa4d70903cf804d70b3c6f683fb78680e4241bca4c884e93c4f71430f343e647b3344e53ad53ea62259df7192da5822a50535aab76e943603da14eba3babf54370f58d29ed770f106f360e4b0ef1deb1ed16158dda519f87b74b002f774abe40490d7d01d1507bbc6dca0cc5f68ba971c4c3a12e04958c2be5838ee7e8f110f0f6f63fd82d81dfba4ca049f68a261f13d1ba39f731ea7da8a6d32a9c444bb5df7aba996d04e92034173fa47d0f7d8dbef39279d774e69bbe1495a7b2a8f6a98a330d1ebe85771ae8881ed6e17aeaaf281b72b42488ec86efd7b8687f142a674007279e0d0da989587e08c9443bb3c4adb6a5179c1ee0ca0bbd0823ca3ca69471f6f4a30bfb94c74946058ecee3cc96e02f1f893d067a588356328ecd1f486b86d314d8bd7accc95b949f72967a14ec5fbc029d7210c2c22b96a540b560ed75f2b7b45f748638835fd1ac4b79237dd04101f0f02e7f58371fbf50f96dca1643cac23191f644fe6c481b2c746ef1b1faddefbc0a18fe80a4bf0a261fc625c6d9bde864ea38e74f5b7ea681a25d704e3aae0c50d8ed8062fea10673d342f8037b2ab6b5816404225a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha699ea895f425e7e1aaca65462013a2dd441ff5e3e6462f46432c6c8ce1bba1d737a68ae657b170322ce9ecfee21c97a46468bc6457071bd1415dbc9bdc3b9fb3e351923e1c709ccbb9558d893fd3953707d64fe4dd810a8d68eb0221719bddaa26d252b9977d7bfcc9af5ac11af357abf952587fa44c60adb238859f42caecbf40d5b8d02fb11673907c2506c69c5628679a05ab9a42aa81702cd6dd61b319381ce601e3497e0df646a59436bb9c92b25ac2558c690fb6dcf23673f95775b6f6d0371ece6e864f4bfed8f29d733522072ced340d2cd34a4ef55f7daf3cea2dbf4380e281833068ff3c4a7b9ccf60cab4dff2f69f672fd4975ad7127129c56704898b13bde942609c17eb16803d9fbed9c909ab2849701177aaf5da525811679757cdb1311debeee838119d5be41741774e668a527a9829dbd0e66f40539d8392cfca190c93a008a423dc16c881179a220283f1add9dc9ea14d902cbaae0881d6266b908d58c3af7ea317c7c78e8532d4d97da082ee7abdb73e6c6b20bfd487d8d330e44c94f15a9d4739f7608808283798ab8514c78a5448549ccdb554d24e35e37bdada48e179ab00b6f00021d28d039d31314b6e9c59f55fe8c28ac11340d39b6a7c0be47ae0e987cd39ea353935aa4129c32d9f67d46bda5d350c0f5d051aaa4e9b8cc13041e6e0b1271dbb6cfe32a694223909a116487f0cc79dcd959e8dab367191200594610b15e420dfa9d272454b442955ba1cf8303690e8e71f912456ebec906b1529b22a48daf5c609c21b2c98954386ec2c455c6c03ee4e474bd3f1d8931b008ed0a5eb2956f4e0d95055cd08a37b8ee5060642d5f7bbf7eb4fd9d0cfd811379e2f93132929e2fd1171859fa02414693c88d7c9b2594301aa61b42895e833cbab2abd172458019a347fbd864317875e31efedab6dce22af114eb7288b1a34b644ddd9fd4ba24c5a7cff8ad144680fe325c51a2b18891b4ce32f6395d75721c5f6df04871ad7f3b61ce342ea14da2ac9b3866b08e678db57fd674c8176b7eed67976a6ac4152c8058a5f5ed2ab5e7ec4d9990a1d23feb6acd7f7466501f569f1e61814b14546969d30847244824297dc60049235dacf3e31382007015b82eea19d4361c83b21d7e2fb11b4e47224e26de881fac06573e51fe51607e68cbee8bcc1cf8ddb90ccbc867355c2b799e767f2a15ba1eb2d223bc97ac57c0fa795d9f0715d4035b3fc9a3ce944e2836d74927104ad796668168cc469128472b5d2650c3e8ecfb445e0b97b3d8ef0b7d2bbf0de5a4d1bc16970ad2d5afd76d73e4eda0ba2f7c0224894a52d4d59d225fd208d76c2212eb50457e13fccef5cd2e1849b144ffa284dbaed27ab3a8732ae85e68ab79a8e9f025e91438a3c7c998b4b7a2bbc8ec6a2b67beebc1dbd3c5073c86e11d9a2ccfb9ac09dbf74c5fac99772e41ab692e6bc902bd2134f95a614b4e8724bee5d1cf1d7c5b0f164a7b325a3e31c83dc5aaadf8731eaaf0c69c44c88e9280a925943922401b26817cdb76f0d9e8320e58545e15e930fc41bea032f9ebcb9b479e96d61f3192b713b4b42a86a1458b1557e97e22aeecc858ac6caf152e051ea8efc3af6b67ea0fdc5dee87d9fe317b84d11215db18d56e24682dfd3cd7783f94c360031459c8fa45ec84ec8aab0a4d42be8f9046785e2a2c0971ce72cdeae6b3fe5b78c888fe3adc9aa58409419cc57e497bfb632835842464c2f97402b1d55cde23e9c66f90bee7d197f7f8fc31c607b019cc3e713a72d13a312da23a012eb63dd2ec5dceef0b6e9873a04ecc176d57ceabc1c4b1aa24a3218c4f14258b2a2d1bcf83a83da5e8527ee39cf4bcc623cd48bdcfc5fad317537344b5dcc27646c4c0ab7ca89d346ef377da2ddaa0b579ce0daf8443d25219fd75852dd3ca009cbf5af98f6619bf297909954fda2e1257c60609e297f8cf2269dcec6724eb08aa47545cf40860bfd9cfbcc95ff48d1431415a5999583bb0f0f9a01a40b07635e2cbaee82abe9348e16da7113aa01abd2c5c49f797a481bebc887909d8c5ad50438d7ea76dcfa307777ede077c41966742cdd18f3d95b1ba1eee1aaf2eccf32f07144db1aa966c8051e5cc2ce08b8db66a90a5d08368995959d12ad4fcbec5f179dfdf009f9ff49515287769159b6b26f58e0ddeaa5aa8920ce74fbd7ce486ad29749d68039f96f529214555ac1bfe7f2f0ef70f95758282e2674371046c499a376ccddcfb5c587367144c1abe16148ab9691575323caf3181a3c4424aaa3e29765ae97d3f4b89125053cee169851d6624902cb0fa8506db65b72d604607335ddb96ecea1fa0f854b527c810f13e17601f68b2f04cde9061a5d430c3a53edff954d145a720d76a33fad4a78e54ffa858738944f2de38a95610fb853f59820a281b5cf65d8171abd608ff1559d6bc3334eb2f1f2c04fd60ee7fe926af48b54f32473fdc4cb89e24aea04ccb304956fa8af5fe6bf70ce2ee4f9b4749aaedbdb149845c837f0b4b2aaaf8c9c222598a01bae5a4c41b70e53e0992e0be25a987e10a6c13be15b945ed79ecc33613b83d3c24149ae195886884cebde0caca23b8cbc2e4d894ea7db3f7a1a3c70d93138147f81d47aead74cba3613243eb0ba14a44a56469ce2412975ad72cbe1a35aaf69a0ea2bf22838e136fa3cca499bf525e524b9c93c2c74be83f212b178a4b151279058203ce10566aa33a35e85a6df3ffd4697b3c8c6c9c90d469c43feaf119de8359214398cbd67d51bddefa507cabfc8cc096c4811f00dc557cc730c6df566aee2b1d41a70b6a5f17a93d9b2cea0546e6e224a812769f1b98a8c5edd63c0ff9be22836b85745f867c9dea670d97adeece4ba39db04c849b83b29a46c86572b195ec798046078add3fb55d40a3bb8685d51d6f8db7500e27fc301f29d8c52ff5479b6f44b0578135ec217dac1e3f50cf83bc39fc5bff884b53c3aa00106d6b9605a082b9273c9346a56bf0ad9096d4cef7d8af4e071d84761b4be096861604709a085b2b0eee0b9d1ce9466b2c49bea849e91d7863c0893eef9a0d6f4ac695ef2c6ed05141bccfcb41d126e55a71cd8e2a9dc5cdb1557edb07bbf65ef8561a31b3ddaff8b56bf0262bb41c3625d34f76d4d0817c517e4ffd409a314c966fa391c4ea2c26dc42d31e09bfa5d9d9555c8e6fb72644925b6ddbfc7a049e8e78fc0f839cd01c497e8d358d6b9ee2df3b7a5d306ed929246d8f1b3629efc2eab5f19a9148169c6eacfeb9d6cbebe2e8b34d018345997d5d3ca865106ee47ffebc004b91b70a35026888689e27ec920d1c3f3d44360c9e0c218948c48d3aecaf09aedf67c20f54a86812ecf735184df9deafe1a1cc917dfe906f5c15fc072a776230b14ccc2afb39eeef43585993bf87ebc7e421a99ded82c9fe2077924773cbda413713ed8d4f703f85d1a2c0999ecbd96e3137aafaea945776485cc41960e00b333eb33eb153a8499425d0343777d6e4ca5d089d68cf7c0062826f34f5763c4956ceb75b226c04c6afce2da44eb1d3c53f718482ca560336ac95951ec67d652d68d9b83ef9c395020e0ffb41cff91f24ee91c9b326a43888f1a5bef0b1ed4ae92270435e5c94a3c73c6986d9912d3a0a5d5cfe818e16a37189d1b606b08e7c1f8ae7597f5d47f7683a43c21c33f64e74287e85fdafd6b561ed48d80a74bfff7ecf37964c2b54d1f1e96dc054b2b7a4d0b30ca1a5b6962a0ee95d667d1f60caa3119dea64c8eb900ca55b6165bff8ab8a9f59ed01f2c2788d61c13c172768ebded81af97c615210384201a7f6c6f6c0f3590c5b98ec5e8314fb5d894be71a9d54f0decf878dcd8d6dc84a27cc0962635194539dca4530705b47ee00c16d3a4c9874a657254b2ed8e02c3e1172f85a08c780145f262f2f406120dec9dc7a4bcfeb722b7e5b47084f4e647dbe4842fd24a826a486e0646c43f93eb72c1faad8295c062442c7a0fe882f4a271fffc15996d450d344c52a315a6a6d7b5e98d30b8fb907635864be89bb42489d40c59d2a16c040ab88b88920e839494bc73b6451fb0ce1169e6c065d3ae110ca2e6c03c11fc1347a8ed60f1985b3db1eb3f99f4a352f9e4362a4c7ff2ea444648d0c0ccd3954ef154541aab4b2778ca82512533aad13834eaf09c80a97fe877ef7e7ec6e2bbf6e22a1d775d7fa8459c5adf7997644f612208aef363e1f37b1aa76e8829647c8837b2a76eba66f2b8e0785b1a1578ee7582a343b7e385647d951fffec680742d06f2002ce6d38cce6658e69e9c3d9c345d51d6eb4bdfb40585fbf1e3b0c197e3beaf9da496b00cfc8e9ce970d616007bbd0f610abe29737f3a13ae0a731a39872f08e5051c983f99bbfca43580a2cb4fc8ea314341b5e5c48ceb7f66d79dfc7a90ae04f89e4010e7a0d28e525400747c9332d456af2cd6fac57aa5e39607e94fd16cffde01622537c637675ff2aa03f02ab568530bbbee03484a48a441403bffcdd2b98ced3cf4b8ba588bdc6ec5dbeb59485bb9b8d4901d7a4838ab2005aff64b84ca2af51e7801b22a6c83048595991b4a99d26f1a7a5cffdd3dad1e4c9f967b6a3d19bd87dcc21a9ec882bf17886d27f0237c4225cc985b2df4b0daff3e3250363cddcd4498d3f1d4bc69c0b6d77512b1382a0f315ff2d458894e54184b02994f15ecdafb99128c4f2503b94a5c617dbf5f95fa3cb414f901cf74ab7e24403c288cf8c7bc2a8cb9a622f0be1e0bbbbb71f4cc878753dcaf76021f1f83d630bdc6c696cfbf41b231aa468c4a5983bda71c5de187836f28d05a4ecea8ffb1d954479218908d608ea79af84342d4d1ede6f52409d3260ddaa664a790579f1a1cd9a1c3b6fbbd3d18a469489a60e03681bff7c194efe58b5b68b056055f6cee7c464b92a09146175ba19e096bfcf4c049473561a078ee25fe88602bfa2481168965909123dc8c70dcb7777b19885975b3bcdd434b3daa6729251a5499484b38d4e6555f4738332a01196a8aeb64cee481497f0e4290b645c12fd585c1aea8576e8e4381dd4ce60e19689da59e5927b4f2f8d589ac49bced0712afe10e9614c5fb86682a17a373c9aa78c6c69ad521b515f7810ec0a775a7097f66753ee019df9dcf5cc8cca38f6c27d37f21495e70268ccf6382bd173b81647674fea431524ad4a6a7420558c453e6965cb1750e3ef9a54c6c78d8d25a0d22560320863efdf5338898202092b91951c23c26c66d8202c74b084084f514a0883ffe5ee509fd0d71227d3a7d08f14ade88fb0f9f55f31f6ecc2bda74bb433c5ea3607b68b403b0e9b035a84208076ba0868ef3c4dd3fb856e55fb38d84058c82c5908ba451b5dad26b80f16b2396e8c8ddc18dd7dbe558b8435143d9115ba2411e65a89869da2bde79f47b67aecdad5322e18db55f0e0db9f4456dd9bde08089e955b9f3f972387bec8c3e585cc252dde7d13d1f2e1846d9b2fb7e4fb276147ea2f830dd7be4c96b841f3853e8946869d35b39610081cc672b0fe429148c49a891c16c1f4ba1963f765a2320441e59681e79bd8a4caeee8184b31747f48319916b34644e11e2c8b6e8ff423c189023f7d45658d24ac8edb5d7bca00ec9e47b18c91e2452ddba6e553639b1047ee650b9c33e2e64a659da9c280415116899d724b73b2170824b25ba2c0d4d0c9039cd0290ce63656a1eb789ca81cd6e5c02d923dd6f01fc10cdecddef70334eec51ccda85e754422851381d8301f90e7a9ea0a7c593326739ebe369818113bd4b71b05740398f76b383381fa1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h24d8498106f1cee0dc19501f8537f2f804851dd614a21a1b4de9e505451bf088c1243250fd263bf9ec0112b2bf239459ababbb4045e7d9fc44ae1ae8737d70b7b16a3c2acd2e62139c3281865dec7e408e5e0bf77055a340cb791dcf082c770da431e055fc1b5cebc3bc70ee6f4808f1fb143bb16570dc57c7001cae37a45e182b08b4e37a46735ddbdd7157efff7ed490ebb6b34ea1a2e64fbd0e5f1e697680fcf67597baff7f5adbd6c9e023cc1744ffb1705c47974e5afa09c636f6d06599bc3e7d16ee9cba9f4cd5670acc390de6b3d0bb075972ab4a7b32033763c9cbbcb4f15260b5792b35526b9175951fae503ccc143f7beb1f60822c359b7ef83b6db849e4042aed4097cd3e29cd6da00191e3277bdaffe9c0f195f8e8f01f243dba120a724b53ea455d1aa04b22b18e65cb4b5595f9afd9a77f810113becfa740fcef9aaab24aec7d9092b8c4e289c43577021fe67ea43fcf46f3973b3354dde878acafd8bcc715e575e53b3f1ea0b78479c224e5bf6ce2d3d5982612c262aa139c9b2485ed2d0ed9383d6d3b2d14f47ca012dfde40a4aa7967535b840fcf9bee50da95b711b1dee41cba59b6ca6baa746ca6a49871d6f59930e21fa602f89caf94cc06030505961c1a4a2d62bd91f27b401526e6afda326cc5b4b6c15371519f2429aeff443b269775784aa7b9533727e4e1ead29605d6a759d6e68d776534edb38f88301d5bf17463efa9e881e2b3d58702de27dd2a729d7b1887a6831acfc42c329d8a61d5b98c561135a418673ad066b7532291b10159a87cee0162047a30174dc9c128f0d2d90893c63ca4b8068e2b490ab61476b3ca0706f84460b698b184e4bd9c122dc18b68d734a91b6bb5f05e45d17b1c0d56ff6c5c7a9ed8019fe717eeee2420b9cb9cef0b4ef4b9d6855b9dfa8b079dedf21d23219a895d6883c83ec916025f73accc74048bf2323591b7894103bc57010eef21f67433406a2a0e610c71797bf85c16cd0131ae0d576899c212e5b40a70e77005f14ecf3587dd0dec7bcfe787c0b426b8f44baf9cb42f88b8cfe2a791ba95aa4e48a53995979582a7266fb4a7e0dc32b9af41210750471af26258abe9537dcf357cc1bafa7c2f4556b2836156f205c8e73c92e29c519bd0ac682924f40212ea205c1f82f63d7c23d379e3a8ae111865a53d2ee090e06fd8f836567532ca3eabd3cb0508740328863f1b048a3ae800d87be7db8d48bc77482afe14cd584ee999dceb07a2bdc6ebe2595f0acc7bc235d6e2c41d70aa741addf8fed3286b2c4dda3d3a891a1041f7a84bee4d2c0b188e8a9d914d6597ec8416e6bb588447e3f4293b8efe32a459e70651d91e5c1bf5f94556aece1b413e0dcd9d8c21096ddd8ada36f12af18b8451a253222f429322b2474e133017921242a9227c22cca15f16e8cffcb26ae3f61a81c197eadc51f8f18a2fd26c5dc2e7dd90d310bc4d49cd913ac26a275cc32973c11620ada398537651bedaf706cda97e01fa4a8fa582ba9d35f0204992de68b30e46e693c76e2c9d0b42aeb0a7e1509217bc889b39f753449fdae20f2f65fc30517777803069470f734298266b2a289a49b01b002c85a970d859233902e79c4f90ee66d1e50784e2a35e65804415f5e0f1f3383863681902829a7ee91cbbf4b43b18b3e33ca5610e1fdc27b537e4e2fc1024c82044d32a0e1362bd1fa92c88615e73a61bc242d4dd153f34d92081981c35d0f5d923e139dd8defdfc524d98d26c34e6b432bd410c7bd6122b62306a1e53738960a5d6b18da0cac712bbb1ba8b9b9a56f611f07684a96c02c8550605ca6fc7f17331d0a8bef13ad1fd6fd019ba762c0c3701ce0716c7f0714a69c28e4f55a1788ed54a72380f1e0a0c4e46f2825b002f09af8ac364022b9247ceb3d6e8edd97de5c8b89eed71af14b5516f869e401dcf9ff527968d8052b7087a651a2d7a6ef28aa57bdae375604a4c14f5f31c62f9f9580daf086758a6eb921b49f1a0c26d9043bb7b87733843b997df91568dfb964450edd1dc2ba1d84a0a504e3b8936d5674cab4085b096c9a982cf0acb9d067a62ddca5f47b067394ce2d67d9341576d6228d26ae4c4a5b432ddfb166ac092a00ff216dc7cdc88ad1500b3ea939797cd1c88e8918129b8bd39c830a9ee140b0805af03918d6c92db9742358ed9e55afb24b9a93625158a0489621e4bc634e687a5a19a1a741c72ac4799a7e862b84d8daee164fbf8f984a4cacd70d9f6fdac6bae3a73b67b3f4efaa65ccf0ef2006da8ac5c69a61846844cf8826b5d4a7dc0f4fdaa6cadd3fec251ed11928f2999162f699d46b5fbe8e13fb43ca93ff3ce04134d5a41ec03feb322d8488e4db72998840ddb3b5be65b668e8ea1c08b26eda69939560e63f886cf71c030f973a2830343e756424dfa5ed80bdecd9edc225abf5b76862e45e93158417a1ac8dc2d674d4ac82d3ab633e28922d072359bd023be3d92e87decb3b51acaf1b18dc80bb086cfe7096c958e4e1beda30d7f8844497e954682eb5b3680e93a414621dbad9789ca33ef93bd0629816d7e54264ae37dff3534c5a4ae806d015732a7165f1f173ed103e42068fd9c39de60859fdace4a552ba9c22fd2bbdbffc7bfa7cb9a8b62388f00b5fa2ba2c5612fa4f7e08d05e3a57917645c899e1bad43878450f00029346ec04f795f2cd15843eb18307945aab8c8df42015b5b392da844eeab0213720bd2b9f52ffdb6e133df7e777d6d218fabafa2bcbd6ed860865ae7ae255d99c8275964d4ad81512fc5d55be2898bd0c3a92b6e16d574b3c1356ef2513ec83febf6a3dcb3ca046923e01e31c203720d376330847c180c18519e502a2f5ebbcfc560f6237a03089d29b551d539d12b3ae460429824f9c24057a49851c07a98a76e53fff2c5c80a6a1c9013998119bda61086c5ba24009db6e8b4f37081b4dfd1ce0ce7423cc43c941a2f9743a72ab396f56b7a401d7e5174ef0cae972c76a3b72424e593862371c5a789a3e3e2fccb3fca7fae0d0ba7f67a4760ed78bb549679369476d21c132f3cbbee918f29a544f9e84db784d9e713a07a7382a902a6dd051a350fe1fe928ad1453844a10ae98f7ed2481654ffab2245694ae0f8e6714e2e6e3d4d3f970d2cd5ab5e8b38feb935f9065954fda3b867b618453c064240856894c7764782e55b4d9fcba3c35f49aea3d131489ff1321079e6c1a7312ca4075e7253db6f0c0fcd266569953832af61a5c5766229c53a815d75b03650eb5b230421595fa5ce19fdf69502cce3b0a41f8fdda72b9e9ce40fdbb70115764346d34bcb99ddb3268a43261689f9a935d1b2c4369bfbe5b3f362e69d177968f49db3bc41b38ed97d5bef02b0db7c90aa63c52a0181674e43873008bac05cc8fa0a621653371df9cd3896d853e36eecb69b64468e3b252d007e03e05e98fcb363154638fcd43982e58b7d055e08b17a8acf6c782382ae0be75dad158fc7928471383d836e5502b978ecb7e31617a44767db0cc61aeb2eae7978be335f8b103185c680a2011008655e74c3cb97e9add07d34b619eddc118ee49c6512e7d68e5a172945b033ce25992b85b0fd6a7da6ccd2c10fe2a81c4fdf14510b946893f0db6f79ec8d4adc0e4dc5d140cf1748e3a9240b0a1e4ebf8ff31e44f63c418a703e54b3f1849afd38c3350d5948a988ace954b9b11ee7e9495bc39af4987cebfffc1d7b42566e2e9bf6e8457da2f54e9f20632e958c8fe7ba080224e936a06f316c3c1c187590a7b77ae5efbef177ec6ef8085e860cf2ff2dafd240009a857e47d55524d48414a08516c6b212468409ee40657d44fe45be991d03f25c126fb6f794be4499644045a71ec9d68f4ba2c11f569824badb88a3a99a9d02ee0b0614829fb9ef5170f70ab90bf84c05e899a44d653cf0514581d9b313d4b5ab93c612f5c95b5f9ebfdcb0a7d536c1341f65d8be985fa3e3a6a287f9fa1467329335d78ed26082bde76cf895c4861750391d7db79bd9362ac55147d7bcb70d0fc1d6fb7dcc1b8a7e5f015ebed23e6c18e9ac2ac10c27b00e28ae1a3cef550f2bce7401311f63eb1cf6debfcc611100d27f19fda6db8ec94d437ef52c7c4365cf0908ebe9bd8b1ab1dbb770968868b113e7dd3d42c0920f46add75eb3dd7c2f5a072f6cc59468e36002cd05ba1b1608b47c5c85726319c7e6763e57c81e024784c20fda2fa52aafca723bcfbf87257747f50fa8b445325028895b863246d1d1a15fd7832e703dbe6a6bf3cfd2fce64bd6afd23ac58902129a252fe4c45f8a41cace6e504a30d11d5c83dd0915a4b922ca03f4b825858e3649dd1f20dfc6f2f3ca90bafc1715f6c98adc9944b5ffb619590ea6e58f37e9f7bb56c7865e81a9bb072372b6a1e08026688a2f8365c3bc1b04b8cab49b0673e2e77b83fb9773ff993df32cb9bc88386156379881f4e753e26a010629a17d00dabff25320f1d33d164bee2ded4d0631be34807ab5bcea8dc787d44bc6328648c73de9324fe83b28c82244f0477fa84fb34a73aa9a9bc659f71760287b0a718c12ffc373cf7102fe9e4167d0af3fd031794aa906212c1f0b243bbbbf18ab82863977de025d22f7393545c8fdc875380908b8810acbf8c15515edcf411f60c90451f59cee177a2c9302a9f1c4396ffe97d47b1d22070dd2db6c028c7459b845f31a407c3b8fc2022b7ec44b230b0741f1c877919cbc192cdd3fa8a3ba7f5752de6819e4138add38c4a4f9fbe08113a48b4d43292fdfaf4ab53d8fa343b162a4a6426081663c4032d092e4026424e283ef5353cd3b71d9a8b6fe3fa3362fdb322601e3dfa296322494d3890b26faabe363750f6bbb9aeeaff7dc994ac5d24883fadba54d57f8b96a76a3bc24bdcd9cd978065500218ae72cc05782b803513304dcc06ccc93c7aef9de05bb0d958bc8ee72214d6834c394ec94ccdaf1f58089b854fa5f84798cb76ea3efab772b4a8f9e28e1f74e54c1385fe2dad78deeb32e4cfed98ad21bf7be41e6d3bd3f4cf179555fbbe5a0082549344163a8b73905ab921fdc2a49a924b073ea8a1e0390a9e92e304efa18e797885395400a0939842b13f464c364ee6d2c4b0bd10fcf6a59f8a9abf0cb94e44616b3c68207eac633fefbfd26f1892bde8c45a5935aa901f95e92ae55a814daeda1456d62c05da776aa6310055dc819703472150b01e99eb19d132b04fc3b5f33228c345cad7ff94bb99fd6b280a7de88773607222043fb1dec2f4b9f771aba3c6d5715fdcf527a7e1bf08eb1ca16121ed3d4778266bea8ae109f98679b015fe5e8d896ab05516e8c98d8c5025a59daf0d6b64103c9caad46619e39d3ee01a01a95475c0d77b192dbde49ae2929dabf57b5338463b98748c481debf396e252fc3238545194eda14b5cac9dd442ce65d6609d59ea4d56b50373102536890b4a9e6d939ac9392e95d2177fcfad8cbdf1af760bad5c8c3bf12798b7b3e417ed0a699848ba422093959f3f4d0465d6ff9733d80111bf3154e5eccbf26a8fc7708e2f2c7952a04849eb4cd9c3a16a8f9dcb3387890af38bb8a3f57468c524c1da6dfb2e501ae08a4b3afcda26377ab7bbd65070576293a404462d9bba7e3ebddf5113aca9392ad17578f11650c7d973e1e048d52af06ce96eb0a73faf14c5789237fd994e1c36fb9959ccb8ffdc7d2e610a57b518106ce6139dc91ae7dfcfb676f41bc05370ffaf885fea8baf45ac869372ac99de9d9ba7b7e0eeedc3246dfcd8080ce76689433d89a2dd4e98935af0e6a5c7547a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5462f400895e646b431a5e7ae42f947ce7a8134cd55bca2341d70aa63cda61b7fa1635a05926de8622c11b78a149063ee2cc191f2f01a0b8c88e677ab2e268af4111a99c4240a1ccb00d9d0ea4b967f10f6eaf8181236799a7a1908856c3336c95c8248e3275493d19ec49b5a0d326a6d442aaa0776334dd071dac04c2e58d2066e0dd34d724632799a6ad098d609b6716d0c8532d2e75fa14e56ce4eaf80d4b6c4722d56c60afb3b982a2a84899f58b10544a6c863123cf06550fc93663ca0c900b21ea5f6801f01f0b16c9745f442c5ae57fd3377f1b0994d6659cec22ded220f2090e35e4d2e2b05f4833b940b0491564c2933e8cd2703b36c14388c13d9656ea0dcdba322cd560edcfe7464469242646823f0db810cc3edcc0573a0ecfb8349aaa540290d2febea2f6f8d93d8774b3985269e337a6af9bb67242b8a18a206792d6e47994f3965c85611a417511a8f1edfce4165d51436db23ff902a0bef1352bc9d927c4508b17197eb14e3b292580bf36fa1673cf508db7584b0201e11dfc7bb1ea0ea8856d98a9c065772efc4f0acf362e61a7d79e24f1002dd59ab69c57ad46cd8ecda7648eede6c266441118ef8eaa8fc05e103b21d8ee19906235165011f0d02a1c76055e802df243c653e00efabc6ddaed1a3b4b050fcd5c8d36973bd656d1b77fab3c2c2c94b496341ec1de15f077c20be0cfb745dc74176e6a23d07320ee9078b52b533d2cf93bf0694cc60d5244a3e4f3aead1f93e2906ac906106152a1b475b48e4acce1aee9a54216920e2146d7bc67aa54da0d2e032b9727e0789862d36a092157b3f35196fd6c8333b6ce8b9f8e856f754c9c590af68b218468273096cd66c2626d4e8dc82a4d2ff98b464a992450de9e30c07901e26b482647c623ae9d12aa784686999edc39dedaed10ba7aaa07e98e0a039095ed8382b3281fde828ee27244eca2a79835191a272fffaab0ffcdb6590efac5c934f2658ba3bae85504a3c6641506ff040f0530eb75fa912349abd790112f4a1b6b20e2ea36148dc9e36b0e7d466a334b1e43b63dbac45f08cfacb53c9733c5f1fb3e3f91d1d293c56e1eba909fba6fca5a8ced478ba8c38500069c99fa8dda62cc120c912f7f0232e00d5a07c3364e8eeeee7afac4977268f9fc791418e9cb26f485f48199aef63cdd0b20089221c06a1e2c417e0279a460cddd4f5f502f8ee1bf0605350d4b363d81ca49129269e2b96dae07294928bf613645fa72b3aed1a8d12b2bdf75f7a17b9b9e02f6f86c5e8fe8dfac7fc4d0d9de59ccae42e7c35caafe9e17b6ccb9c4f1c94f9fbfd60d08f20d9b141bce7d0594a3c133876fa04fe7f94375337cbc88b6ac77c54c9779e38a8c6cebe1efe7c1b23666c44b8dc1a17c75ee52e7f4031142fe545323b8b4d5cb8b61d6925eb83f9cc7ff5c3ed99357499cfd72e3c0a8244298727f503870f704801d5d2ca03769a9249c1878206f4be6f7cab298710c3f7bfeaa4444f68dc3c1a6021c3ba387ec14d178976b905e7ac2c85f34991d7dd61ac9b095f1a35dbd3792f0cf998819c7c820d72d701335562cd36592fd3edf0434fb15f81c807338f2d48e01fb508d0c0179176f30ee48a00c904a14a01e1bc49a9cc26f2137788720915cc58549acd3eca3965f387dc46bb618ba87daae003c0290906d443431d4403e1fe2b16166b805b9a6aa79fcc9966d9662dc8ad8e55ab562122949f0456fbafcd58a95158e4a4c0bc59406f0d14191235edae13519cdb124d8ade2d76aa662a80f863b17c297ac2392349c5566bf968bf947682c104efec9e11417811fe4b784ebe67a048bbe8ff526695c71213b69c72cbabea25e597d66aba509874b5cd94af787a9d4354d26bc3d856ab6150d320feed536de3196d2f784a403d094bb55178a777f7a7d884482a05770c89b4eceab1e98ca092835282671682e28df3890aa0004adf4961ae9e32f9c7fcbe098b57d4065c87394f5a9c5f17258843f508a4b9f5bbd931dd5bcd5918c6fbe8bedee96731d431f200491b1e07b293b0b18e881f05ae3c803c4e9bd1f92b8e204410c45e163a8567755363c1b3e19a54ca290823a00fcd236e6934d9581b030cf602c34e229eef8d933707b82cbbb5e6875db0b44e99edc1dd911bda4d3d4bf70eb514e4bc353f4defd5589e1b3cb8562ddc8ead0649449f91b876b4b6e75aec0466d988044e28341184ed00a8f6c81807802fe0dd100e6af17dbd3e176f9bac8c444e0282b02096d4366cf0279d16b47e72fb83a2afbced7129ad43ecf57268c0fabf2ee551321d7f89b188c24af6415208e01b7206d299cb23ba87de785c5e2e51476a1b7d5d09eb7061d8fda0386d19ba8c163c0646bb194a6db7d2065cb7a175feadc2dc131d6062d1731768d90542ee35702223c181aed391a9149edc8ccb93df284d244221ea6081e4c1a508fbbbf6f4b3778a6ccc480c003aa0bbf6b3ac0402f0fd8bd66f5febf1204b61b81558a35d3c71e42b50e3a3be714fc826c4a0ca69f17a27ec06a6182df0413aa2fca430735ecd57d106d97ce0fec623520db80f94112dea71b49469ff4e5a01eb69a1d5a87789f3c3c294efb87591ae2b8c96dd1c2f43e9d9b18a32b4f225933ec9831c19dde275e3d13632b23265b3b9a734fee120dbe7b7af03d2a0c1266522332917fc6d61c2752967a8b371be1ecf50c3927a965fe96b48a9256cac50b169d49efbad1552f071b9f8d2f8396faf6209d2242bb12131227e0d8a2f9fa823d5378de65f4e45ec9ca24af33c0a6f11570bef1c89bc3563d16305fe2d7b879c4743b558e0d7538fe313b194ff0362d19e1c765666f72e6f7c2e8e1199234a43cd0a9cae48c188f107dc8fd20bef3c547fb3c832a03df4f6cdf27ad9764fe2fc8d36d7ef279a76c5bc1517fca40a7875c636687aac5fe0ba38e0b04bccf2a8aee9b0a75f5bffbb04738ec2cc78cb1652aea951a7126cef36fbf0ebfcc608514126c78d3dc7ca7df149b588fe330c252908ff79fdf4c353713dab613dc7d99521b9c159efc3ee2966e526c9d3230a219ecc3dc45c3cc23eea5bfb0ddf79944a143543f1d8b506c7f0826e43bb02f1d21f2e33c473643ba476c1cd88a88eedb4c00690f57701e1049e71892e6be69aa51a32a3a140bc0207e6793431a83c7353ecfd1a3ab8f8b70e70916b24d83a0ef410d31433c4bef9e6e842734f94e49af0ce4b483b9f284270451a63ae8f0d6f1863117139db1dafff7d6202cfed26214d5aa2cf37adaaed09eb01a7d356f0d6ed39a58a38b9b3cba08fbfb0f33dd32f851da1ea8d56bad6a84948443db2bbd12bab9ce133a663b63869522a9e84c8b81ae7b36deefe32120bfb9bea4ab27f1375f92fd03b137ae50d09b174ae81b9b245a66c357eae92dcfd306bb06946c2e8d7da541f0e3edab9b123d63190e0871e73764539a3d3aacbc1b69e96fa118b055bbef7340da6025296b0a79f58fcbf83d9a161afe411bbc0ef50884cfb7464398a547cb834c824e500fe39259dfe954b24e38f661988bb714f14d1cc7c2ebe5b19686f7a2d7d651def0ffda8316f594e2518675866d70b809e160c3e6fc3375c2215fb9785f625f6736a72816061957b0dd6616582db3f207573eb12fc539201e4374c2286ccd3d3d4d5dfccefd326663cced608f2c270cc90814504424a1a6cfcfbcebfd7b7051dcf6fce6c1673d47a720ee2ab2613b769b0dbcf8149b4a31ca409d549950fe021963133c549188092b55041697f1aa8612dee5ed3b4d488799d76d82f5f1f966ef4d8a6e7a859c9a86695c341e5e0ac3a63b072bf57198231ec59257c511513ff1437e29671fbc1b3bbe681f2d82daf3d14839f6a14e64d16e2ad963e393825748aa91ffe3cf09d5bf30cdc31773bb815fadeac8c1d8aab75eec95f0672ae8501339b94ac6b483524d7d03137cf2b95a12bba3c011ec9e962a981a5d7b204e68ca71325a796e85e149a33247a6819bd6b8fc7603c4bacffd621d4872e39b1d7ef832a2bf2aff35bb42f8fc9b2bb6ae8eecd053639cca00d9cbb7bfedc1c9b7dbac031fa3bb8a8317bc73e079b45867e52c468eda3e28a2c73a6bbaf9f8b10b5d54b0f8bd6270885113b2d32c93992b7cd6ab1b98b77dda18e8ebcf169bd5537e01135a88fb8b5a22c250887220d5b3c40b20de6ee874a5596f1e5b6dfe566782ebf46026ef80cba69e4cdd5efe8992bdb9be46d45cfdfa32c9411fbbe0efd1dfdd803810aa1ff40b3b9d57fb481b3d88a29c0620253228cd2244546ee41d66b00039288b6ee99fb76a2d1c2bc2943ed690c8bb50b15f67142d16045b995a5f6a50f0252fab0a3466c9c7c4fb359e3ac179270c3c028c90532338e41b9d7a67c513e066cc700c168b42f6a8ca3ef09605b1632a57603aa6954c7f8f453eda14d5d5fef97a9745c3d08f1efc529a8f9cea9deeb0bc96585f48cc80627c42dd70d61ac18b6a822498a39707eac390cacd89df866ff54bec4cfbb5278d0f5569ad57b85cc082ecec9e61cb8b3b302735263d02d738973cddd7c8bdb9596905cb31b8ba3d149f323be2f1bc712ed02c6d5a32d23b7d1db7de474e2e3b1ad278d1af70a5e10e6685d507874edc6139b8f34847666f6221092555ae46d7eeabd253a57933314538b05cd2a437d85fc50af64027de417e0ba550566d80ba4556077e747c00f9b1b4bdb7852a5a066721e5e26ee89b54a76b2efed87f5bdd5658cf17e837b9b207c06f9f2cab45bf500ae987cf43819214695444fc414b23804fb0bd36b437e4f5b56a0338dcf0a7b8598239e3295d860e6eeff8c97aa92ec65b18348f2b1ed964b21af52ae482b59c99b81c4c75dc6dcf883d4dd76f7de7eb2844da93440bff8fc37f668b1b1c7f7cdc19f5d68b66235fb3f439e5918dabc31caf7868221e98725be812b5c9b45ce8d8c2d7b46417728c37fc3b577ed5eeddbfa8d5748d003cffc637476362eb0d5ab73c03294e8f2a47b1d67edf0d8a3d9b7a4dc7ce5f9d9741fc5521d3c6228e6bb1d15cfaf7dd467442a1629499ff8268f57833218d5b243093db405de29f70ca771be2a8c65b00e5030abaadb7eddb2f0bc3729840a5cdfd49b71a932bc9af737009dcca406d3f52450bd4916a9012b2cc7a47472ff0a9eeeedda7d1f0c5d558ce264e04716bf85de8f9c8a5fdffe55986ead6e70f9153441d03c34628e9a601928aed3026052f028a9618c77ff0877d3065aebb00a898228e1513fb396cd4db5a6ec49aba7deaff0404a6c6c91f401527de0d470813e3389603ec71f96772658c43c287ca377fd456fe09cd242b1256435a4b8345209f14aee4034cc50c7ec5d74404fd15f186a60b3c31a23be62ea089ba3da692e9da44f4f6852e9b604a07f84ffb9f4eeebfe99d54dc2e9bb7ea0d406ec3f379a1857ca5ed18d545030f031bfcc3419d8ee1054a284f0960971d286987567fbf6cd881a3083aef2c88c91bffe000d39d68381b77eeea2f7275812e59290042a6499030bf284f12865de2d7e1f7c26d3935a28e194d6eb4356b209afc027839682702a58705bb7439cf9a5c794af9894ff9bd1a24ee205dc474094dd607547a7827f0c381f90ac0d0b0651e673cd62a60ca4aed7f7aa11c57543431c5380c707ea33550b82f627e460dab32f9c38e540a50bc26c78ee43e8446eddba3b61b24272b7ad9cf3e6702f42ceb722f76ba0bc450b506f11b7780862e21dd43f408241c48c2b886cde90fbfad26f988b250f0473175492b46381368c839a7cd550d29078769;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8857062a3e21a12977964cb09f60db3bce5c2c39b85caa0c6a3d1929eb4201d37ebe0474d05fd4a69d8e1c7988c7d3d833b33d3a8276c898e0a2171f7109733c2b58f73e852e4f0aefc5f2f015e63804a44e09d006942e95aca81a042ed1e9f078466f58562f101040be6b944a553a7384d8a815d200c05abd235581fb72167f2ba7051cb53e3013e937a9bc35b2dd28a77bc0cd6bbc976894a2d132c4991a5b053271e900e4b9aac211d4b5fcb434fb4f39e129977289f297f641d7d532de2c2ece1c28c7fd25305f890aa09f2eb06f52400a6a4e0a2a349c35fc50cdebf60fef1d5619dff3da7bb848c074092bb8afccba232a9610abe39d722cce64e0b9c186d5a49c101bc740f7a6a38397cfc59376dd907edba0e466ed4b16f7e9dbe0707e23543ef1c85670d357ee366c09265f04a5ab8c27921b6303ffc090a915b49127e12d67269db9a5dd0f6c6ed4c8883ef74c4ccd739e475bffefd9b90cc3ce81666df1695a6cf303b2945489bf459276f19f7a9c9f424a642a65843e2daa3ea994c7e309d68af1c3846594394aa067fca6b8b940db81d54238f1f004651e312301e46162315dd7329596cd7c3f66a386f57c49519a3dc69d5df4aebc63aec0bb22e683870e24e19528fc6e978fed2383d4c76807f16dc0e2eaa83491b43bbeaf8431ce09d23c3b20b4fd19dfd89e6788ca53d79074ab8e5ec3cc3594a96cc7aea5840478c1516f59c8f510cfbee51d2bf65343f62ab45994d00d5fe269c8dc7d614023ee56f18f427881992c8bc342c6b357da76aaed587acf30d180542db6c989ffd70930757dc069b4a8513567c88a56c9493a727db56a9493952cd44453d174cf0997eca33d719fae190ac69bffc8044c2d8223f6e7577adc9d5fc9c74a33ce58be6b1549e8e115b6b62c7e73a5057292c8b1130f7468f85679d05933e85d167dc2340d2add8bf72f139e776ba6eace1539263a596348b7142d98f528c04352c5796ee513ae7a87af57bdaa3623cab027f15829cd0512c1f88ff1fff9b1466a37e0b26fd308b3a6c72558ce53fc7fc8d335e932446036d437a87455cdd768f2551bcbb107d686cdb2decacdd90a912e2dfdbc4b6e730a4a8ca229030d4f1c75b8f3db1187954de8c9158344c455897fad633e706fbe529927e0ef6e659460ee8472ecb2b239a46872f26c33aa5a6d0aa1134ab0914b8a2c2d2e25f582af3767fff7cb21e79d36cd9282d8f5a001e8e415b15d8df60b0431bf15e131b03dd3b6b6d3b7782ea619b0b81c3f6ad40826ab8285d6ab999c3bb2693a8f00995de28d68baac7ad48c15b1584cb27c6528f73ccbddc3bc5447e2a0efbc446b595a4ab3126e745840df9949b6b5a68678d3f8a3ebdd3fbcecd04d1bd127b96c5e9dbe1c60188863dc8b050bf8fb37ed0f8fc9ae697af931134ef1f1ba19cdebacfdab27b7d1c37c988825558a37559aab93bc90f26f9ce8d9c2b4433b323ef2998278e9b3f7db40d6f81e65d63a9fda31aebf9a9247b5e6e1250fe22d4a8db22b503d3000874f9502789d9c0ba2a91a9cd904f205d82fffefa7e61da2387714d57d03ba0aa3535b1351ea7bd92cea8cf34d85cd5c6dfa07884cd857ad61a85fdcd1eedbb6edde877ba8cb627ebe349dceb7863554a2d82a742ef2671691781f101a6498b1e6f5f8cb7d0c3a9864a0d140269cfb22c3324b5f6203b77e4492084c1532292f6b53c8253a5e67d77697bc960045700f835a932bc5709655982258cc08c9c18f093af5fa3aedb2c6887f427f1784714588e8de8f937afe7730cf3b83a40f9bcc9c9c42a9a757c805f5e52eb5fe92c5a4bdd5740bf53968533f7ed7e2f94db07eb54330eb3196115352292df1d1e4e89e97ca91ac88e36b7299ccf826f1cf1546d471e26d34286d595ddcd1c3f904e203a2b1033a33a3dbdbdf654a82e51917128d5376feff3d82db099123212c0de9d45da9079a18500115e419af5c12533ca8dd12bc179efaba61a33abdcacf9a48d3a506fe6d0f9ad6162e75771c8dbe31133793796513b2430234b5870ca51bde8fb386b2d44b9bcbf7bd2bf0c5c0ebb1b6a4da56864d2e316ed2afe6162e16d9c89ad0e84d22a2454797a385f8037c32b7164c6e2015e2d1eaf8599ab4bd73bebe24c5386a3b75239d8ea180de15cad834f8953a393be1dcb80d8950251778d820901c4895bf5dc354a4b541e15fc656b5f1c64f525d95ea6c7fda93ac75788298c8484f031858f9a5218f0d4e6f10718a93318e6e6ffae86392a7c22cfa48baf9776782f602e8ad1886ca1bebc27484961f11efd94a80169ae5fab3f9ebb8d10b8d757767003033dd77465defeb1527e35f71d5fcb54ac69c532040479068d5ea57ce9dc38d8f6eda794f49fd1401a648220062aa741bf346ace5be57e2e4b04ce2857d413112a3c9fc389cdda7e7d96a65f925d354beec1515d6d51fb91541445f34736ca40ef067b551060ffde47361455cdaed87f7fc434d3910f138251695ac29d880c26b369b2d3cbe0319f8c8573e77400c3b476e991bd176828decd492aaedd020c87de72394f68c9cec760f1e4124bb70c1960e07959ca04955af547d4c07ad33e288e81e61b74823b18e773c2d8c5919aa1614900c4b40dc5b9c3a2ccaab950d3035560072279c55b531371f594ec80633b3613880c381732f2a9ef00c38b3e7bea3a6b80e2e8fb33ff51ea5661b2d20f15bd3b3a931ee6490f0d15723827b456768ac05a34d4b9fae6f236c0b4fac78f24423423a7165775a79ea5512e0dabfce62cc276c51e009526c5c1613c45a150f0910cefb5cb83d1675a8fe9a59063ef15d5aeca5f433c50664594a65d6f14b714a0de419346d6ced5295f4418f6fddd9e854b632639fca6dc698434a949c0cdbd7f812b0a6b476e763fec1d8d6fa42e27cf6f489100cc219e560e0d71e731744ef709a1cd3c4129fe4e9c584cf77628b354420f17f4f4868480fb94ce0197743c1c2a12983e2bc94f28d8f74677dd5f7c88b9cb717b5bcacc9dd783aaae64ed634b18c76b2a448dbd006987819c7f84b5f3d98c4541d30ca46c5f5adb2ee77b31e78ca65ae268e87398bf8932144deb717e47aecd1f352438c5ea67ce8084da89a10750a50eced9deb1d772053e009a50d3bada56f2ac435a53a9a0c41f9ca73dd93a8d3067935be0d0abb3e40c02c0361462ddaa1166853d20dbce83426f3f084d9f5b22ded581ffe27c965580fb3f2c6b097ef03b113f53c4cb9fdad48537c1dce23a5dc3a611f159955dc17c1ff1efb039e0d2bda3f7068ee7fd7930d56d00da528aac0438d6f9f9994908b4823fcdffbd5b69c4c1168e1652b76779cfa5b98846d0f97cb6a58617871c117f916d0d4539f768487831a78629b5427fd7aa269232edfb75c37b40951b23de21a88d575286321305e62d396ecc4dc3ae0cbe0e47f21c76ab0bfd32baec67eb645f1cd257a2cfc25f36cd41aa471d80d1d9f81c0238781b33967d30cb3555d798f80493dcf3e31d91689a368012373f45f3750dd9c7100f09323a90f70f04e679b910669ab419d8ccae5b8c0c54815d2db28f81011c13e4fa00de305e28e3f5bb8bf59d27218dfff151a905a3c3cdb95fcb4a042af7a23be915b0282c188f122d085a918fdce0169a8b281b98ec472417bd305fb14bdbd37172e7a0da8ade0516d4d0a461907e07a715c6982b7771b36e2d97ec29c84115a134ce24929a9d998f2cbd64248bb73135892361bcfaf006e1424159762e5580ad42179298c108c47b4fd4e43947fd09acc4ef87011e6662927f0bb5126500070c0f556b613b78f237f3cb7bb9c6a435aa24ecd5db9c6013675ad03527efc436158b240842daf9251bc264a142a2a54afef6ec8e2e2c3c9b4e5a2aff04cb9f8878e07ea5354e0e2172ebacd1995b7456de088f057e7cdee03f514b9b9a9fa92df6ee7e030216397f4b35ee7b46e1029fbbe3043724ade97800fab65450b435b3491241b0047d2b5bfbb6cdfebb413676866cdafe00fa2402b4f04b838bac53ada9e5defbf9ed7d382c8a61a1c97ad62248516c44b84278a2193160572df4fce3d157e66e9a52745a65282609b9122417ae8994e20ca0934810057fba5c3d2a5eb663ec50c0c8453c465b2621a6d429ff7c240f60489e27b22cb08dc48a124f30d96757b02f894fc793215ec769ab3d1a020d63ca698c56645441f7ab8a9b1320b13fc5e6d13adad6026289b28e24f482eb8aea7dafefb5441d65500607fc42fb4e2821c855f202c14f90d9b4476bba35a5d18681881d125509099c6e3eaaa66794b1f9c268062c56680df163056e0ddd4d47391d689f1630386f81eb78a276659f2184b13bb023bfb43010e04aa487fc6dafd52ca4e4bd9e7a4d6b429eaf7e1fe3f8f36a9de1124f315da086b85d9a6aff7a3a8f096b7f2f0e58ebc11535153b458790a48f131d54d06bff135ff687a6992ab30daec299f47d6f037a7f21cc4384f355d9f14ecaa32f41bfe6de2d02159a2ab7e139213dacb5a643d1ea1e72a6e6ea1108429f1da44f9cbda80b7b2102443c3f090f1c118909310064566c04817913c833ab9c7133e36ce7f2be5dfe04fa5d3c43a33feac0ae17a6f6d7248b0ae95aa6f6a31fe1b78a13048a8fe4debc45aee91331f3b61a902c2705678ee2fcc1ae21ca184824b66e112058f0f68089d3fbd1ed1bd9711ac001be3de1ff690f1b1e9f6f1983d13c95e203edebb1af72932c1016b59122cc2290591bc303c2eba0e595f57ebb8e9d83118a3536f2eb0da01b9ed50fcc22b07cd92a8bf8217765e096942875d35c5b0463a5ba217b1cb5e3ae90dad304f2363bfa75d28accca98f90d5564962277a731252ff4bf340dcb706e5eb9c64002bd3227c37f6ba922735f33ff19fb309003ca1a77105a2d834fee0d3986a4bcc738dfa9cfa00a17104484ceef34e3a8ecbad6dc6778349e2be424b44375f1c68b52085d01ce9dcd1741203b3c6bc27ae8ed4a25e1651e5dab91a185f08b0dd09edfe02a67675cbf7572bb9a8c39465fc5b12b55e70432a20b6aaef9bec8cd8b4b54841d20307e47f6b556c9c1f426640b4300b206547583b4aebdca018985a15eaaf5dbb7468b0efaf47b1037f61754f873c39810ccf6ef5d2d8050cead996356978416d4447744c0d226d5529e5d72249c89a81940f09378af4fc0939e2d0694f9b844fb3c511c8b996e03637ded2f69109d9a63e4a3737784bf0040419d6253b3c17783273ba92a81617ec4384ba6adf94d981e1d2931a079069519662d00b834933e75ba696a07768428ff3d629210bf68a221fb8f6416c76622000e31ae4287cd0c637b97849cc60937a408459056ab5ebbb46a9ea8424c3640eee9a222a9f4f6de7ff1c38739737348e32431570d191201ccd6a647243c94bc69031a7a7f340ad29439928613f362df8091e2c1f89eacbde38a1b3a5c1a933988c0a8137149c6eea41b3209ba461e8fbe776c5540d2cda4df3b8099b8d4724a4dcd16e48b5e8d20f50cf76cde7fb3b69bc7074bd2c357acd2762b1fa7819c811f3c03e03f88a70b648fbfed17444fdbe637d653c9a6911dcf1055243e23c73d5d0ed90fbabb7c250b15e30917456ac2a5c6dabe8b29ae3ea4ef17260eff6c94643881f10a80c6827b67399cdb51ec10aad991d5dc39f54e8389b95f247508acdba98ac25e04b7a4e4a7cfebda7115ebbb8170be730b987f32461827226d6e06d13f5e3514d1d2b07aeea0303c55887669d91a887997ab2c10c4fa2e094678602b4a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h40bbd17c5f2b25072911e77ca60bbf8eba7293c92076f0e3e5c62bcb50598b76697adb6de7dcbfaf6c1409c1fed30e5d17802c19669efbf79d5d89b081954f9b23be38dbea2df79347a66e85e613a4f7b5438126c7568524800d33893b1d46c4cc30bea778b7ce30fd6afc1425f1758eefca34c53d9f1a3d1541730d01a1945fee53fc8f7b6cd582d08ab07a36cff8a7e6e9a7666190bb2b0ddf896e1034654f928a5baaa413037cc6008c912057fb6f3221858a5a919efb25cf4e635a538925d55d9f3998cf302e18f0dae5c6619e9a072455f855155b1168ee1db94f4e9d8e5d9f153a23ab3b6c642d636319508cb464ce791d3a2f4eaab9a412c24147a2e48702a9982de36d2f7682e6100a97ada199a5574d838336c5cf48f399f2ce886c181761dba15db06df3f4070eee50bd2526cd54661104fdeaf96f8bc37649e99f93c6807c232fb1479582c3ed654b628c7949898608168a6cfa5f6e9affb837a398b5ad5ed2d20f00ad260c0bcb43ee992cc01c623e2649b1766244e4c3abd18b1738554cad5a7c3a1f3fd842686a4bd72267489fa9869e25212c9f69469b63d82e4093beb17f0e2d9610fe34db88a4a4633656264238f28225b6c4aa42285caadf1a11560bb8aafb6ab463522491e355e4135ec73fb809a427f000ef3cc39d22fde9dff6938d330fad217a83ef4d05cfdb6fb6bf5d5d37fb560bf6e3355fee1f0200396260217e23453356f0e919ec8d5671e208ec727640e45fa6ec1f7fb55b609f5863eda44bc1abceb2f69cab357b97eabfb7dcf6b21df63f8263578a3d9b47b3a608428c6770e9936ab159472144d1ec31ddb7074e309df874968457d7910a921ce7cd0f2cd0ece3a524a35e0dedf25c48dbb203b4d6738f2195cc95e544d85c93713c000be396110fa0c5631d2285b49cc4c092e83a7ff439586503f043e052df53b4f63af67168c6026ee31f96e3d0967ef10fd28985c870ca07d35776e1730aac08abf7014a0a145e1aa6dd63d7b08b653c272af30afdb51d2af5b76708de78d0a7f04f0c44541b26fa1c7c728e2248331685aeddd545e0785cbd2e48e1fc7d81aa7b14c86fd86f9c13bc19bd1bc11eb3a87002f01b9ca4d21a5ace13f2ac474ce4ca7915902c24143d199b0a3068df69c3b804d6b9db6c314c31df050bb6074e447f9bdd742487dc9bb61d991954e9c08fa6830e1709eb49b85f895fae279ffecf4a049ca6c2752750688602bd39510e93b1e240f43cf654a26fb1deba37aa903a8a9ae24a6fe4d4c2c112dd02a15468ea014d897cfe15b89698c4037345ef986d78099cad65b2d6a320def618b696b83ce51786c93678078e734416ff3b87f581d0c1319f927e57ff2f02db1f3f8696424be03087fb4b8c0394668296ea1e0cf824b2cfb400827cbb96c3cabb3c67aa1b2c1bfb01f71838e62702818d9539d78c6b3453d07c2ff0e919c71e8b515cbf324e71409d46242cc9d4466584f38cf1442eb8b698607667de6d444628fe5e934f4cda8a2448d1cd6d6e9b1b0f04bde3c6cb5b657634ac69b25d265ab56e2cbcd39838d5ca5831e6f55105668de6e80c6aae0dba658ec3d23ea89552ce06fd661640274bf7f3882636702e5aa9776dffec2958e18d5e5e9149d1725888a859c963348ce7cb8a0c4c1126ef5a252d1a810b0feaeefb6b900d8f155922cfd189714b17c2790a3d372a132d94b25c9a4b184d49ee59d4fc0787268c89c407232e68cd32efba322b06e2890ac5747c9d902fad32c02abdb944c331f64e8c4df6176d8950751a3ea2c346a701526bf9eea356e4fe89da1451d3599f3a604465c2713b270a7837465643887cbfb25e0ff2cdecc50dbe24d8335375bf668621f646acc3660607d67a94bbe85b6f05261e627a18934c85574da22e77b42ebb23025a327da4e6378a551d62c2a4527fbc6df23f6e1bfce0bcdfc15ea0ebccb907c915e3ccb1c69aa3b5992a3c623643a8324ec7e77c9eab35df7854b89090622782640313b76347735f65972e60692e9ee98fa7959968dcdcb2a045a89dddc7beed58dda321dc64520eca916da586d44fc2c6bed3f32edd78924ee36086bb1a51c6421c37ccefadbe1ab835ba271dc2d3073f2f9139b696ccd334257615f468b58cac54a0cadb578b65c306025824a4be8eda6e7d6d836013ad7ab12cf4535c9a63dd5c4a0dd450d57b9c0ebc1854d711d937af8bff6642bceb617c0e05b76f919b6f12504eddc15a2397c1d2d998e217ba988ae68e925a95cfc6f4de8f774fdb3cdd600f3a196f3f73f6409491d5f5edcd7702b21368f304c76a807b44da9d7ca347fd4f0c734cf13a6ae324687af517b3b15395365c8cfd34c5cb8686737011c8cc412077f8e138fe972c30902150b79a92c7dec53d906600979ae931000d7c80e75079a59309bad74957cf9830b87a5fab721f7424fd0e6379f0654dd346e999b2986d6ede4f3da224cd98d08490210dd64e6fd49948a3c5317b42b106b963a2bf22eb29daccfaa65a82f167f80f9edbf08226936014f15606bde3387762380bb6194ea699a6ec23760f1c59d623db5015e33b6989ea0c2a40546c6020a17f6988d4b8d0eccd3b8c6d0cbf7cb18b98bcfa7fc2838abadb75b68575d20ddba3129d66bb0e36400bcbfadad74bb5f9ca5a8ffae8c060e523fd7075213151853e7a382b79c612de32c0ffd500f48a644cb14595712ca87d911a98ba24134cfb92cd81e6b2123bc4c197b465320970404dbe4dda1be6feb40d3095b8b420113b027a7dbbc3739035aa2b6091143a4e34b3afc9af1dfa52b30e0d35ab81251348e1bafbd8cb04e14b401d962806202ac29658aa4d1a4e891f53a4a466e2a05f5340f197d6cbd4404ccbf4b455faa16717387a73f8f93f46be81fa16db29e448f9196d68bf7f74c8390cfc3ce8b4cdcd92f0b4617147758693c01697ce0096b394ae88ca1e80e7f8f2ab984189f562ef7b6a9096cdf7d95416bbea027b37f6931123737ff9bda577612ebcba40dff1b3447771226a64445064c554b0d784bbac3d5af2fa3d8fe67795269049ceebf41cabfe35f3212d047bc568b32b62b83602238bf932e5d6f13df48d93ff4b228d88f5dab88200d2bd299e910b12ac1da8ad203b1ca5b4803e229dd902aa61aa144b75de82f98a03983fd11e74e8121789c396c3f6068a4da75a9549cd7eeaa4bbe1fecdb884642fa847eecc7db939a178c8dd935416f802312c3af52a657d0a8cbb19cf267ea69a907de0e2648c61e74c98764e12b36edc48d96b89f6469557538bc8de27e7cf89b9275a4592effc70a31a9c16cbf6143c93eea3578db1fa4119c9676ffef2cf2aee1dffe7a3be25b1ecd96fcf9513f7331b774020fe9d5f2566899560d5fd8378fbd4f3097934d60cb53b34afc596700057d552bd31b656226926a66688e5bb08d06d0d5d122e7df00fddb26dcadaaa371eac5dbdeae7d3a4328be9d00ee5286facf477e186835fdff295259f6589729642455217c01825fb455b6c285bbc53f5f806d8f1053133db0d2729ba081345f817307d3c75f27b23440cf69864fb1e364d3cfc385d8fa03677871114e3846737794c239649f6b766bcd176ee06173b9569d1cfe81b7569df2e3f0eadc2188e9aedfc2e75d2666274a19b0afc300b4673d5c7f30c45faeb106787a98c2cfb9f7c9a34f4a5eaf3fd8df3d1e8e07c5d47735ec08cb50eeb06683d1712dd0677fd0bf092db6c4654caef12ad2f126abe370726e0a9a9a98e5c291e7b340954c2804bcf1948da993aab6565041814a9ff9c98c79f7a3336a2445fa44c7215f0d4f4e51d1235622d7f2994f7af2d20200870d3febfdedac32c743ee3205718a5d146e0b8a9b3b9760213f430d7ac5c3d65e722eab11c0afcc2d577ef22df344a6111d400ec32f7a0f1773f5a3bf66efaf640429f9e596adfbb4147858912bbb57e14e7638e9ac542efac500b49c294d60131d8e639d5ea75a24c8538536ec3203584dc7c92e160cd62149894853425447cced67cd0f7add110368bb8dded57d101136a2f72a2fd352b288080bb652dc4718f4159533225b2df980478b05450dc6ff0a0bd75bdc46c61d584ff7e8e7395a400bbef0cb01e1d3581c9cee49b95c61ae50c8a123902ec4d01ff20f2b2de669bd6db3ccc892a310dc7ab728bf667aeb8379f5a8afb11f9678a5ca136963c57a578a2748029802c6d58848763565a991b297729ac570cf051164811849aa3e94e90112b46c3ff7017eb6e4c2181a9fff534a917d6368e0aaf35a352795c057771e8660641c9d0ec7ad39083896e3733d53be374f87a8060142e02ef9bb85191dce01eeaadf68acacdd82303524ca3e7aa89b4a8b6162d649a0fca03c58f752ecda0111226305996b17aae7d6be9ac422ba231f2cc31382bff62ca3f476e01bb03976fccaa402204edbbeb178f96aa7e064431fdc32be3383100a6e1f27319d4e550aa5e0d547bf8965e85c389dd07dd7028c9b84876818d504a9c2f1e44aa333fabe92192272fdb671a1ecd7e7c7d12c3de89be91b44f99f4c50a06b1c577b5112198d6f3079241e0e6fd2f50d3a33e5a458f3c1307102e22473b133fbc3a0e1d3b1efceae5f0de90692afb5f7cbd80972188964e3bab48167f161c01ca249ef8a470ce79508e8c151e2696743e16a9bac0f4b6684a889d51bf231ad49c48a59b607272c8389e87a17ca3bd20a9e38a59806c1c6f2b86f10cc75d7f55ef6c43806075e958f673bb3dc4a330b2fced2057fd6bffcbbb971897a478824aabf1e3af442d03ab10722ca18b633290a4f91bbbb501390392130549a661a4c487cc1da9a75af34b95df86c50804afda82b4605b288348fb41598ffd4e5a2f015d646307c7737198990c36847dc08e9dee4809505286f8cf892076053c27960b98bb562eb57b0d9d2b61db92364548f2b9ab5df74f5d106340f7bf35aad99d159fa30afcff1b578f02a3efed43f538680c6f542ebdae725c299b59b4f5fddcf8223ad3224c8b03104327811c0276e3086d5b89fb6880c617399d0f6db9d0c4d9cd3825779298146009b2951ba788c1b03e086de2367e86d15c24bce5dad8cb1170018899e25864a3357de17014908606231f3a8a5e4cdd30b458bd70aa9b3da729bae26e1e1403972887ffda20cbb96c9988c57b50b4a3f7c3e3e7b7a99209018fd0b9119cfbd3507d519958ed41e26dda33a12c3016dcffb5ba24a603a64dfecb0d84179b45ddb889f8fd4b727ed4aaa1dd150f8af7d9a9930bd21ee5bbb10c4fa3fac45a0c9adbba9a48434a00e1197494275f07fa1249eeb1185b573688bb66e3fa9170c871122adb7b789df145847c1568c627be12dd01baa8e1e6fa69fb927eeeddeb385facb2291b956f9428d2309a9562c59f7ead808186bdab1c413652b9727b1b1d9716c5d6f736f16b9b19397aa81cba7d6089261341d370280b749d299bd470fc8fd076a9f9a535a70396dda7ba552da94ebcd4f2a7d40fb6df3210e7ec1de542b29e4015e7bec676fbf97392aa444b347f7f8da824e71ea73f087f8edcbb4c21aab55ff5f05fcccc22cc8cf10f6c6aae7f83ea0c145195f4ec56f63091fde0e4b07d2403a23704642067ab52fd16ecc0384678535575a1e4d905012c2e51789d3bb3b39873c5136d05b25537b405dd196ddf040cfaae02a1d1ab1d4986c11454e3fdd8b694ab278d25a4626592f7c542abf1d3605755b0a235ae9701025a3cb45e0c4f23da09221216f8e754b00570ef3b3371d0d3351b01c74e7ca6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb06b4bcca37dda42447fd92c2d71d956bc5939c53e75a1beff5d50733ab56d1278e9391fcae6681ea83c2d7e4da313a97bfe21d73847f420f46121ad20f3f5909be86015265e30fe7711a0b8c68c5a607394f63dbffd27ffd1456f1cd465cd8704241cd02134d994eabaaeef581b5a3f12d8bb24de97ca46bcf7ea28d915c3f349221d54e7970db5726b058cc19bcdc73ef884075394333a6a13f229e27748d06ea3012f2fa8cc31ca5d063e0439d4caff9f2a7bab7242a0580af943a77e2985b679f05d719f8c83f363b8c1a9d3d13f0093f44f1ee8ee8f3788ecbbf2b3fbbe69999a41545750b85c80fdb6fd79cf5d0340b6c6d34dc1cf96acdc88efe6900a929be3ab86511f6ef99025e38bdb13d57c10b6887977d3b7331f23710962d7e310ffa902cb7744b7cb629273798c4062d0f70f01d64a27a595bfd76f4b6a6338680b5e4a69202b6ab7429596c5330544289162192e4a9999abbebb358c0bbc0a5d52222a342598482bf8dc31c5c0be789a2ae4651e986631dce3797a993acb376d94dc93ac8895cdb80f2a866bf6a08dcd3d1fdd475b9543f02228ffd0ee375e676526b88da5b2750598fe56730d193d1d4a477c1fe172c58e63f92b63fb4bc5ce89f581fb6ae80bd43e5d2436ebeaecc890dd4bbed1740782f190d44dff56fe7a3fee23be6d12aa5559ce45d6e07a53901aaae9260d53c6d63346987367a45054f42ee05aab888dba6b259c06b53c505cfcd0de6da329929e7fd11a0fa52e2fc8c6d0168676dce7db5b19669fe70d14d9160dd15c8375034222e955f8af9ef236963ef383aabaff1372f51c1c7b32201ba538a0f99ac292eaf7de40dc8683c164f4f2031b94d35acf816dba7c0cf10901307b4a3d28eae2a2a7f5ea0135ab322ba54f47f2ed6e14cb7275ee3768574e80ad32da650b5e9e10e5bbf4310aa9633a70720a6fdfa2dcf2aa317c4b14a7e9a831dd3f40cecb2c4974020d84b0f3a432647d9ea2b7c1a8c212d82e2e8962921b4b25f48362d87c53108502d03e6c35ac119116010543d292ae7376c57eb0f4b692d9e3a3b26d4e5914c4b85ee6087337444a5396d7e40fe5f976a35e5f2ae82540cdac39f956573ec841576a64ea22c2d0b07d0e3351e58a69254e73581aa4d4c57ef70b88271f6ae4f89b9175061f3294f7de212d937ea3f175c91f9cb551459b7623fee433f9cd00b4c147d22a4a94d6fbd4ab380547ed76b7619dfd312663f177e6e9884d5f4eb891576d76b60b1fbd5703fc470143589e3c8e7e291d9814ac88506c8c1e792bcbf400c8b0108d55236fc2c808c6f81dad79133359c33a5f15c966879e04cd3738a13ef99bc872a8c11b78c9b9a84c36c19bd287774060fb873ac070902ac34d2e2afd2613db43818571698a46df686c6d3eb474276a7072db02620152ba8e9cafb53a84700f63728d6e0d1c13561d12dcbe90cd50fbc42b527e98804702a986c466283f090d00adb91f8639cb72051f2cf2589c42ea72be3d9e927d1bd562974a9a3db737723727ef0f4b419ed28acb8befd6dbfa732091a702b26c357cd22218bbc0284c14c79a09066854d491b8c20377e382c60db51aa233231195a6a6b02aff2016d68af007ce4fa3a6f0151625b5acfa09060643f5a7dd667da868f0567f613662437f718ad05598e18831bbd7e3e8c0cd3b85254ec5c8b8c6873a384ae68c2717c42fcf5fbb5a2842b1b76dea9cb1e1aedb089d5e4f305ce52a57265d0cc92e4fc8410f1fd1d2377645a412325b72dafdfb08aa19d7f2d6c488ed6d6c0036b2d402605c3c00ef38305a729197f96849448b033a211c5f6b3d1dbd08643ffb617b6fcf66eee3d162af0dc028d391eab89f41e3de3878068b6f52c02246a8d58833202c683e17aa2bc897040c09631c585e13deac071df5f093e97014bacf69de18a5b96c808a5db4bc0b663817467564b3ed6a0e30d20f447c64d505d5e88e1dc00c917a30518b38950070609c8a28749b3d6add159f32652eea11c7415d8c5b71670cac9298e3a225c557e7087b3ffcf9e2e39d36962f4ecb5cff100dd3b93fda725b8e945a580fa6ad7d3e5afe6732338cd8e24302c2581988c72a2616623709229f11965b7b3c4af3704aedc429b5975ba280948bdc1c6c5de89ed746a823f92177f3f41c415c3a5fb6504d1021e5a3f9e1d76e4c68ddbdbefc623325137b29e332c5809564787f001912f926ee62ad1ca895cede6c22912a58895c50ccfb433773dc6824bd3a787faa5012b3d5c7e9e7c2404adb7f9c4de92289a2ace48ab631175ff0954b30a174c7867a9eea6262c2dc7c01206ea680aee7178b431c0d17706820bc38615ca3e255980405082d5fd3dc49b619975e0454fa3502c4bc2d46718ef0c1b58fe6ae94515ea7ac3ddb5eead522c284ff78b511ee8b178960ea36a012e4c189248432cbdd05232fa30b38fa677dfdb2eac5a03549cb55a76100a92982fad2b05b8a1b717a6ac2ce1ea458f508d5b42f3985420d512c5ced48aa3cd04193eb5e31a6dfb25f5586b6f3c084cfd332ff8b5abc65061d4edecb0f6a32428a28c7ec219f560093a0e003f67329eff2867832d270576518b2c68b5583dfb554684f5aa1ffb8f41ab826d198788b46a7719470d5403c159ceca427e53defd978e0aa44591761f951f0fc2f24a835629b786bca62334b5b8eb02a2aac0caa6d637e87ab6cebe6181c9d38c351e7684a22f3d47cd5d1ea6685b628b9593ce7f3f271d72abdcf650f070513778d4ef60389b5ee323016c3d46b5890af36696d383f130c3cfd66377c2db5afc62e301042445fdd542b2c9091ff6c3718aa0f0cc33dbd882c9ce4ddf2f81988550f873c1dd8d6f15628da0d4a15a40803b6c3c205e544ce2c9823a72b4a01b57cac68f42a0e398540664f605fcd33a82525785e3bf0945231bbc05415c41856830fe8d94a1dea1727e5fdbea2de80cc9db10bd3e65953da52d873ce5501e5cfa7a0992403aff06bdbe0cd43799b80154b71783ebd76fffb2f6820a5fb199867ca8929a55858cf2a13c4854982728b479196eaf7712be67d300d9a6c02c4841c059fc136b46feb812e113bdabf2f933ebf287f4ebd1a1bbb0f9ca8eed614e0e28ebd5f5fb4d710484176391027b3e8071fefb2355c150c415b1c7b2c681ca36ccb22f8136f18da76fc3a8b1b52141097182126fb5880a548f57aa94912ac848ad4ccb78f3e7d884a8609fcc763cef55ad46549c53faa4061f3ab612e6e93812bf5a54c6aefd87b4919782e0dd090542acb401865c3382ab3fca7ebf6bfc4e7011879d1d402f0a26a327d4de518575da3f57c49ab59daf984c0912263423e62117728df710e6c83942cf28f99f5584252b829202eba64ff444b488b084ff4b4a94194e57055a81ec4a61a59cb8b7090165ea23504d380790da2256c13144a86c3f499612887c5e27139602db0d0f3ffb22aa0c58c3a2d71b1cd28434c2d9b0644d21ab05b2078042d1bd6995b5e557035da6abb5e077f9b3b2370969e6f54c8c1ebf29953136d3368359ade5ca57b1471b66462993add4e8844490a960dd9a73ac3e7d28d70eab6c1263c297ac0630ccbad4c64bdaf505dac6d7a98897a4dfacd630520fbe0d5c660fca2ae75c4830aae72436c0d811533c4b045a4589d33839131b01cb78d67399cfdf024f7911d7dba56a0b7e8ad3db2bc71d4379dc199be3dc34381e72dd0bc22989dc87c4c8f35b84a9c3cd607fbca7fab53f47c9288ac62ff04fabe52d958524201087110ef9debe1ea2426dba08c312cb826f96858c5d0fd4eb75151fa2aadba8042089c190e89f1d39e9c59de50a398eaaa7b5d3c6e595af904d8ce9714368c50a94c21919b3b05119bfb42505cd739f9a54698501d56121411597f6385bf6d98574373d49039801c6680da449ac624ebdd990e21b5e5ecc0d73c342f88a636e7ee3a2f871a193a3094cc161e4279f139343f2cea8c536842823175da4f886e658bfc0ab631dec1b5b983ebec3c38d62f709807d01210489875277076a944485adee0757b05771ef548a67568413acb9eb5795fb942a36be1f59ba814a73cca182d8d90a64fff905f0401007e8d78c047b034b286a0aeb0130795ea6e66542fa72dcc93709110ba25584419e782be7beb411e1a3f8dff40a734b464a7ccb552c01e6060dbafae5671fde14d8d60ce8a8ea10e53c918fc395e16e3fd96c0dc7164ce05e51e02e3c66fddafcfecfff489ce68718cc5952dd65a0560c4c50a04fa73509a3086b9991b451db33e91caf54593f26cfd2cd1732b9f86737950c18f1f44a0c8d043b7dd54a66fc3932dcb07dc996ce56fb3d98d3575c708883711ddbd2952ad93acf342f17c756466a9c9b5ca75f1c60f39a404a81e5b43de4c0c83fb609973d457fd6215f1b89b6f3c5490e2067b98a4d6c5aecc83ffd807490b45ac1769a7d2a35827858ae6bcad9122a28e3cccbdb05c46873ebf494bfc7b29e5bce937a2adfb1406c4657731ee47959703869ec83b59bcf5efe6d84e6451f2cc7b1d7cbc97298dfafb1cc1cb6b767543e2b3029cd167f624ba66d17eec74de73e3988afd0579facd90fc293b12ce2872fe88fa7cf30f479be5463f39954ad79dff4aba1f8275dc1a3bc419f843082048dcfac5159c75c3e19c8493b0900fb14cfcea092dae7dc083b7b1682ad116c4fa81588b9c894e56bcfdf981f5b1d307ffda9bbb7201596f9eb025fe717c765e642b8f9658619ebf662c429abf4936bb3dc4bf688c65b718209d2e429cae68e23763d0d336f191e31c0ddb054e5e4790673d6a2127434967bf012464be5bd8f99fb1b7f3ee852d94edae46639e777fd16c4fb615c7fe938774fc0a8f3ad0ecf615acab979832261ae0ae092ae7cd670fd39b3cb64ed2cbc41669f752e6879ff1471123b4748127b2aa85f25fcd4f4f229ffef05ae1b23feaa0fd007cd5006a5f2c6d3b345b2c145a1791b0e026005411a5674523d9afbdc6b27deb3d3d1e34eebefdca76342c08e580cfbef211b80d7c3fe6ae63f0f90234457c1e29c1c0c68e6dd136dd9e6c5363983771a2ab6d2be575339fad2ad532e05a50321839935b1252a055bf2502bbebadee38e6bd31a551d90bac063fe30f3a40127ee01e3e1e497b27bbb0b826fc6fae73ad6939fc9155a3c6284eece1c0d1f538ef9d79c754cb64b3a37777f6555cd41dfd1b2a4627c417d1b589cd5d808b8ca91bb652b493d28dde62027471663fad4367c05e99d28b86a853a45305c2d773b0d932fd792dea4fda7e73617406922fabb0df7146a3f1fd1ed8669390911ad117377d12277a75412efc242506abd62050ab84a8ad6c890e9340fff1191db1e0b132bd221cff4885289fdd27c0e30b59a5da8c6d16f0584cd9e701eef8e49bab3f1108cd5f6b092d5ab0ed4326c9c0755f4ec773dac8ffaf5229207c47c54b7cc71d2d33c81ad193c8633c6ba4feca212d884a9905ed3ec229209b9917faac32fad92ef1645f00a7fd7c7c1fb34d8125a4bc19de4720326616b144e7b0b3e5eadc8a73e691fd7ac75c9079ebbd878ff7fffedc46df743fa58c83c9624c3b7259ad665862605a2a0c839483e2f7f6cae9d7e2ea657e485f8ee020092b77a1f7831dec8d441a86d6541f67189a2b56f56d7aaa37f7e55d0cd6279793b892dbd41b09658c6a5be5a6786e5440defb87eb23b0e02096586ef4e12f2fb0673c6ea22169b4ba3e8a4b01f9fb01e5944ae998569025899b1842d85fde0b4ced43d2a96a6cc8edad8c35f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd1e9e01472f5229f5aa520fb073c470b67415dd67fcda3fa0e2e9797c30253fc21382a0b632956a5a34d2175507c5e65c217e1baf04b30b40cdd702fda8b0e001576bd51cca737a36a9ddc5bdbab1e272596fb7bd1fcc6da75ae79c2001e5ccfb5210beda21d80a59ed7cf37333b608b9c654d134d9651b9b787170660c41d8b80658a12fb69d86263615ef93e37dbc0e1d9afe61f8bc97dd0fd6c5490106d1896c064d30dfa8341c18b8c929b53d08553056c9445060df4def2a0bb14c61e7fd635280a850fdf3ebc2d0bc8cd77367b69d7a2d10f7e428b5646d9a25f5208ec14e748c89977382dc89e5db75e8cda20471dee8ac5b2911f4527661ae97babf7d677da49d4b7b6de82d36d28b04455ccec58b9a9028814b944c5e69e17154d6db5bb4430484ccb539cb2ad2c55530a1e6f186512ff5f66844488f285a67f61272b03149e3abd2208146c0d36b584ed75e37ab6e860d5e72023dfd5931a0ed297aaee8d6ada716ea8ffe03e2c5a05516014a4159191d41a7a6a621b2ac71eda4a98dba0fc719f0923c09eb77662b95f3e59d114eca551f8009aa0d640eb14251a5c834226ce33d6b157f2b385b77d7207de4b2af461334760434169a33c0c6327574659d50a950c54c85bf25686316a0e65ffbcd5679d276efa1df87e0cedc960ed113fe4de1493f2bd63994587abca1ad22140cb23115596dfddbcc59d361b85f46adde60e7f83323c3b5eeb964208b58211428f5d0b2162135da66e2dda6cb84364e45cb7c1cd9a2b1659fb660741fe5c3a4b0e79a2e6556ba27b56d1da24d5b80758a19fc7b6643f90a185fe568e87e5cc9be1cc0859612ada02a6533a58eeb40e6b350450ae0c038e5fc0a8fa3fd512606b744e600fe07984f77bb3de495aa79861bebfa16ddfd78dd327122fb56876fc26f98e794e96a063f37bdd5ae09c8349a90097b9fb4f3a198f9c44987eb8d529b677e20bfbed88e5741ebe89fd14f789487d0eca9029a6bd81131ff1cd3e4e49e8a9a0ffbd6fff013bb95f86d28a8ff8043f43aea10ee1f8129e739831bd19499c0248f56aae325048c8fe5e13037b7fe9034b6eeac9797afaeeb7effc70c9aba20db05eaa25cd517f1d7cbceaa9d5d0386c1c37b6de783a24925757e0fd3d7fc3ca82459fc8670ee8e9f4a2ac948d9407575ff4554e9923a2c75b9b7691312118b6d1c3bbc0b92bcaae3dd2182ba079df12c9cb2611b6b0cf97cd38a749c10d8a5072d8fadc2ecf18cfc7c0d18557334d9b0852f766b2bddccac4ecacfa4746565d186b27e779354cffbfed15ed1262d8ae5220850986878dc5ea291aef31cd6e0b7722f90b8fad175c0475c98c501430f3322dcd0a501ca9599d7acf741a1a37e9715b2f4ef7a690aebcccbf6c6feb0505f5bf2b1128769f3140d5223f28d8c325c62c9dfdb47b2b0404a12e012909f8700595c17ea7e22e07417d527115d626caac7016dea762bb4690c6956648f9334a30d692fdc802c9ac6cb41e3ff3addc88e3bb49af46825b531a46268019fbf4f3ee661854075c3ef131d835ef25fa8d2cbc3f4674d2184e846db7eb78825d3b9be51129038c22d2133eea503d014919795ca680b8ffeb06673d1f9fdb41f6c387a014e5d21ae4dd61b1388e97c5593fa41058078f6eabd022d9b663ad8067c2329406db1b54e2eeeda5eeaaa766e337f726b2616c4899844da497bee0828ad6267bfaee8f893604c325720c091006a7607c58c26a74d2cd23c8243f3f162901405676296c276990360a581c21a8aa84045ef3da06dddbdeadf1d6684ffb3daf03ee109de0e698feb21604c64d234cb529baeb76b2980aa07d236376cb26302468c0e3edeb52a7bd1cc0ce593f67760cbe421d7daf6f9ee94415fd2a5aea11d3dd6a1c5fb7dee60c00d2bc0e0c5b5723e8a6877554e53d721f49247e06dfe2eb5c7ab28c05f23e37d3e954ea1f8920e4725a0f28c754bf280616e5b3ad4de52e4663a7ccc18016db8e8424c786727d8d325cd032ad08e310565d1038f07b337db1ef13257d874f4733b41c78b620c761bff5461540124e6c8df57061c5cd654a036a38bca312fc569b6edf75d8ae5715e7d7f36d2fdfdff22ef1e176ce9f025d3bea1a70926e7e29f9aa9589ad2d16012b1b98bce68bac0384f6fc8ee288ff5df9dd3ad81e112046af6648e8c6eb5402eabf4da7f78cb202dbfc59d7009c8af2bdf671f3154ba57dc72aefd3c296d2de4d4b615bf4c8f5cce8f8498ef3668bf487a82dce569c4cf34231d88013416429892f869f91efec4ad1f122c1d8ae6fdace785e81bba39fcd14e9f7ed97ae9f03db2648f06b2b6b35145abcf038c553b7cc428fb31a98da7fe70e44a276f1ad0b508f81e0ea84c97aa544c29a0f83df638cbe44cbd8b1b2aef05cfd8d0aa55c9427877aa28c3e7575da87328c1219e1ecae96a8b07dba4017905c4a4cdb7461cee2244af273318faf1cb6c5d3c90ecbdbe46b2177de0666fb4613dc130a5c3102eccbd62300f36e463f946bb1fe5fb7b06f5e4959541f621202783926604ee2c00b59ddf8fe9118216a6ace470f0ad75db29bc16febf13df5dd284c323dee117855578d56a18127d51393dc98890f7342f2edceeeab686d6ffe676d9307b9a5e02736989868f2720cdaa0ebd0c517d7bc8c78f7e146cea1a8930f109b54189a366d51edc636d7519ee80c61e7578d65bf4a6d4af71c61991b7b27b1599ffaa20055143b0aac8c9d2b37e65a3627f6c1bc83a51d6f0c6e6014c32e01241b0bc2251275a49282e9bf25ebf680a0f463923e40ab630a57df241d0cb16adae20b1ef3d187f0da789ab7d347246dd9bd6a32aab195f8a3f4172b8cf5b3eb174ebd98646b26cc9c1df039ab286d087caa8637514cafc5e0e5351688efe493924bc9b30e7e83243d227c26d84ddc50412d8233014cd26b499aec00f838aa20409f1c5fa4f1f5a1034efc184713605a52f10b0c5eb6e27ef4b341bc2040f76d90c604c8d4cb28a7ef97a808fa37487780f9b2ce785856ec139789ce8595e9f4fd5d22a25c266270cbf656c5321ff9fed0f0b82a22a57093613853b1bf5dcd7386894893892a186b5f3217aca05ba93de32e643bc80826aba07d53d409ec43fe50e6fa6349f68b2d7c969a57d18d259795c34d551887924f8d50fcf583656d4fff45fd976cf1954d8972f0d10b6001a2ead8ed6a69d602c8f9bfe0d88bd21739698e54276f171bafe979991ab6dd26b72868119a88c3ceb48538090c3daa58ae5ad9592a0148bb854a1176b94cd5e28b8c1272e5298fcfe1b1bbadea8970fee592a8f756548c0af7e8b330bb67f047ef82dba90930ccf4cdd48d21d11b35b299544e45ef079c7c3f137f8cada6da93b6802e32633bbdbbd44c2cf11b09d159efbbbffd474dccdbc81790a2c95fd60c33a1b1042efa5eae7b323b497bf246c14ba89b2c2cce69a695eba36160226fb07b84f811b22902a8ac87feee582ec15721344897f41710bfc1ff0dff66190c0263dbd53f48568e92b143e1c6146be8096ceefa17e07e8634941f1f80e4851b1f222388c4d9998ac13b0b840afdd5b7d37dce11497971ede7fa26df5877e564af0aa90f98394fd7e91e521d36a6ef2ff8443b9354e2f41eb2c09a9f94663543d6955469f02a4f687a05047ac93e3d70fee9756eb7a6c526b019217f607bbe87e6262bd0b9f92770a2d0bcf3b63cf329e43f54132bf8dd3bc2c19e77ea05ef60ba9b3457d182acd8c8f598de6d62a30f0fc6f3f89893c2541c43a4052d5c2b87c9a060d51b54598b448b5141054dbc890410a166afada4c97d0cb4b8e1f02429e0ef0dc45541a3f57e260d19f402ac2f5aa0980a1464eb0bbf17dacd0e4905630f1610df615983d5e2754605ead8ec0fbe477aeebafbf25fac16096fd8a4ca41c899652209a567f6346108985d05a48274af5e09f10d306c87f6d45150e4fa55c87c8f88b921f34584ad5a89f799fd725a0a73917e17b3ba4a04a3b83b610eba72e86fe47d2a8aec44da8078a4874f55235560c2792502cf49938f4961b4585f39f88672e36eb0b42d736c6fd5b9dd314039810bd1501e277a3cff784bfa77b880b05238e4a58395605f5f34fddafd93c8ce95b5c416cf7daa1c9101551ca37db8f583e15fa8a87245da7a8e89fd9249d6d0a4ecbff421b4bcadb419bd252e477e663f5e42337e052e05c2b230469b31ecfc0f8239b344a5e509fe6573975163af0ad424e0a3793bd249c7796b5fcc52988886dd944f353bcae94a3bd9c37dbeee362a77664deadac1f90eb213c5e6a15aff6d1fa54dc81ca244d7a40939e7531a2e7c94ee2064d402f15fd8f3e89eed833bd086dc488e22a937cdd74b19cf5937aa9e04550c4e3d5d6c1d8f107f8e04fb4ad5a3e3e72617ccd11632e8615d1e3f6a165090c6d8a09f037992289c591ca2ecbd0833a20d54f5d99f30fcdfaeffc665d85d234979f0eda399046415f012821bfcac8c6a358eda184be0e1bb3532508d1d56d604c985cdf9e1f59ba0da2bd6bb706a757337c43f7f6975b15ef56732e1476fed4872737d4a4373802614a29fabfef6c8b745ba4c1bbdcc991b6e5e90bc33d8321f3bd5878cd4974e411fa80f9e6d578edb60244f1b43c68d36d7f84f24f780dc500d528308fa4d37dff829b034251aaa25e984e7e48903f9e9d7831046806602b7eb3f8e5f55d9fad2d3b744bb46a34d165e08e357d9b035ea3569604ccbe20a9161300fb32e70d70b8b04833a0e209f252f0ab8a14c4f820883cf34e874c92f236459a0c8fdeab1357497c71035a456e571df7d74010f67817ee85892a507cbc4a54225c4962e81205225fa658095fb4b1c08ae8e616ecca25a52682e0fcdb8ca7aac8d38e2ef400dc8db90b3278d0f6e958baf59d4bd656d0c01a97dcd81b759b32e90a24b6bbebc4cd0ee4a39abe7d5dbadbfe4c8424c547b7d5766f34806191e4aa83ee3b59cce89cece8502ae0a2069793b8c95dbe5254dd0c27a46c14df028ba06aa2a247604ba2c5a4b3cefb396e2ae5619daec6c73bda7b851f46d79988342e6e871ed1c096ce4763a44e7b4febe21d10e26c16c46c3450540f8a12d1cf7d3fbcfa50bb080fff06424a78f9ea0da1b96e1c92b8a543a78713afc64c6ff9335f8f062c81694d71e8ebc99396f3a86fd21a9edfb1fd2b117d7647e33ed5d1bbc4001e8e6a3b6f5ed46bd136d4d6f28220feb17e682dae6717842b0a31c0cc4136a33ac6d2206a1d323126a4f960846bfb3a73b1e4f52f5679ba54bbc20b14040cc3024006a7192bd0c8fc0f38494511c6ba013f4f635c99b2093ba84d1db47b1ca18556c03dfd71c2c18f930baef3626928db0e0c5e79eff69d3db1cdbfd5a04696d1d8ba0d0678e8243729b57ea220e66f2cffd808dffd9cf76e2c2de52badccc0f8433ce0c5b6d2c84de287ce599d812b0da844094e760e8c7bb785f89f50d995925caecfb880e73d5a88a006c67cadbecfa90bab82747133aae54d9559a0129edcf0c120f9b6bc7b381c56ae410e7fec9b6e82618cbe98952b51e6dbe142efeccaf7cdb43c21d13c838bd0c707da3acb0ebfee6ed1d99381ddc702326c04e4092fc8c81db6d4ac4a456d984160c6869d437e757504a96f311293b1f467f42d58b70f80456a25f6ae9189d714b2c6a3327d44e0ade653d5e343101410e7627604c1b43cbc347b7ab24316879727d5ac1dc69a17b0046d04d0a03eefa98c57d513f38e9568c21e848a58052f3f50f8fc4c59a011d7039d69a8ea5ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcaf728f76b053761d42934cf510ea748986f00029e72765ac9f191af2f6a7ab5c406faf7ee427d39df96990bf832203b48c8a0423ca764b8fcd2ea4131d617fe11f8d8f65ba097b7847cd00e3414ee1ccdc3de5ebcbd0704219756376314babce2c32e349a3a1bd4c9a66b0cc77365a4349db099c470d1dd19e2e1439bcf83d049ba2bdaf3b8e2d9d9d8f471456180c1c9128a83a64189b3e68cf53733fc57a49a02f51481e6963cd1ce63158790bd9486610a7fff4870fd38935063b9cb3d836990e1a3fb9e126f8558fb40e3b0112e752a9cf945c1f06fed20b8801ec07d1491ffc5af6cd94c20ffe6a5883db886d28e2295371e08ad698ad1fd146414fb8201acf981a8fb8bb950080fb0ed4a98745f989fda2ae53be40a5aad45b225d6eec9732911eb365fcb66b611f455468007953d824966c5b6e7365ac414e41b5a0f5dd0a6cb5cf8bd9bf2ecb05a87259647b5e1aa0145043ba6f84d159198cfeb32c65c746d4ae3795564c32f727a8b1a5594a111b716b954c20d7cba0569fb4f8852c0ad093ecc39be37316c512f5a106033287c715516c09be07ac005ad5239e7142ea0f94a3bbdf1894d2ec2852788bcf86ad161e7729acc34ceac2483c8580926a1cdf0dbf2d60360ce632ac6d678b40db813b1ec083147d8f460a1d32261d921c4ada2147b19c4084021975cbc2104e21d3e4c4fd3cf6768a9819cdb98e83a47f9d02db02af554aac21e94aa222e1eef6827a7e26fb874c3838125e77f99cf47ddd3729d4280bd8aa826197d4bf102de96f2da2b433a197a328bf6533ae88c20ef7a5b5590b48d02fe82657b92d311b15a6c3c462a3b7d78fbc0f74362305b59430325752e5c27cb0799296a7da9994ffc66f6a7d99345839e9a243206ddc305e4578f550b6cfb4f184db474728c8719c692372ca1137e26ff4e5d812c3cf2ae04535ccfdc19face3d5dcacd55ba36a6e4cd16aec8f005326e4b073d21c830bdcba5eb7e651ebce4b8ff7c0b70836dec48292d74d3edb5c217f4b84332cc9f7c902f66fb5b6538456931528be23dd1098f2951233819a213038c7be8e156f51709a71eefc7ec4278888da367128477bc1ae3ce75cf2923a263783b9b5d6ea290be165754a8eeabf20d98b7cfe1b33192e97cb5f3aae48b58a2547225a4d83767db31a00eef956e5b936afffc7602f8e0d72a5a401759d365f205408d633b3cd8f4c6ea556ac122493a82f31d3df3d85525a66dbbf9ee8b2dc6b8a65ac360e528371e161413211cf370cdc4d394dfcef0f8f05ad579020963cde9aebf816f98693711a58c2ee142076b5d95e99223ca88f19aefe90fe7256adceb5b6d501d5a5eb24029b197d6555d58dd5f1db9a5c66dab8d83bd5ecea1ebc47f36d6aff4d44a88db44c489478f55a857ff0fc47da74683b9f8e76b9a75157fb9c0e88299314615b082c93953c383a0273b955ada404b313440fd641905fb963222581dd6d11a991c4ca766d461c29515e0e487ec583e88ff98a450730524e82357b2c19455108257784380e8a38620bd9524895739390c93b73ca80f1957fe7fdbdc01658ba8382a4adfaf65cebe73d644753a0718bc5a3a509e7b2d7129f2ad186cc2d2f25d24e773ab1c2206f94d06051e2d7fe0eac3f9b1f45e5ed42a7ee4519d5339692fe226f21f31d95f47f672dd05c1ce23b2d40a71fc6fc20101cd4f072caaefc9130fde727ce20d934e5fcd8251ed7b0cef8cce035bafa041c4178463350f36f762f8e820d3ce54d2af39b4dcea3d7e9d763a4b7776a2d1acc775d108dc87067ca7e427be3fb241e922031eda4b8e6cf68dfab23e250e035d499e78ae76711702479d6673c2d01561720598e5e66531de6aa8784af011995a58be9c13f123d074239b41336c29071ebdfe75e40bd7d03067ad1948bdc4294bd5b86ad4a7e883481081003e27c98f77e3f91c2a46d982e17418a3550f2b011dd7b3eb25739bc7cb5e04e4c806d9bee7e3cd9c58746e610dea70c9ccce7c1898af2fb29f6a0fa1dd538ce4093457e4b99573ad462bb84101db7b033c16fccca9ffbb0526d93eb56fb32553fbcd8ab6fbfd03d4ac1d82519064d958836e79ca9faad12b27ba2514149b6cd5909e03b74d0e32b517a57246de1870455c535b1f6e0bcd62c4b988dfb9b218bf6dd96cf4a9630863c2832509515c8745df679797b91229c979fa204220f14bf6ed652a718da8fbba525065e7bb4d636b0c5bcf0631dc3457d70d555bec543585574f34be81f67521c592e1aafb67336ad567c23b3c15201c13b49be18e91e1798a23421ce711346eec617fc4bfc2acd4f1b730891dc0084148578af8452266ca6cd38f693a1a8271d9c9860f26d5b03dff0494794e0f83407a468b06b6d874794489c21e0a83e766941ab3d9877df931b26bf357e8e7b39f5eb70c8cd9e00108d8b5037f0eba98276170af4658e7d5b56c8ec439f236fd288a8984e09d4b0f14e902927f8d30c47bda0d68fa4e42af02f99abb90ac34bc918e4b65a146927cf33ec01a168451d2a7f715a4dafcbadfd91a89b3e817fd2dc77f56413042a89dd1df23efafc58e65f571355e7a4c366a5c503491b9e10cf18c389adaec57539ba3c43b3ab0bd907ab22ee25d37b207d1c65c1f7448652ef3bb6da53d271dd25ab5835035738473c754d62ebd55373c07ea59284faabc1e24d1664d61903af1c7576a6d3b0ba95e5decb661230626129b74fb8f312c6f560c8a87f4a6fb7c82e13d1c609a627a30ac88675574f80ce7486b606a4005a966ca5fb239af9f89acd712265f059b0857f297049f6f8256ba07a6cb84edd01692d399e7728c7a532a875a93380115ec1be1147cba77404bdc796cd9438c86fed3abd90d25244f725cdbfccf03e54e86ae7856bd390281294154d83463b6f2ad3166c73e080e7b8a2519af37345b8c87e7960f217c0fc14c7d8fdb267b3eaab91f35c5a24c44c5f5fb4e391eedb01790fa8c2a8eb85f68dd6a9ef0d2de77518a30b2f2ea530bd570fb4002a9b4e5e8bbfec6d3bda83f92aff0a88194e7dc53a3cc3f57e3c648f913a240457b3653d3b5a267911a1e506b677622f41662b8fd3789dc240d44f70b2f0bfbbac06436e865a07924755bde70ec88e5f1353f477eb1a67a5b6ea6c0ebdd5380ca78d2d8563a7d0b056d0f291273885dd843a47dd49c1fd0d64b6a4906e5ca1118908543c46ea41f2a945a4fd118cd3e64f660eb960db4b907045fd4811fc4521de92ab2d14aacfb1d36451556e5f70fdccaac59874434be1989a7c93ec619639254957a37430dfb3e40ed7fde96a4c4f53ebcdeb0882c228c6638afa3f0a695a4fb0f7af9dc91d02a28b0755025769c4ad8fa7443584f89a60b02122d2342a1533defd47e1ff8fc4c1a9d3a03d41c0d1995f90346168551357c4a72ee0ba3e5c9588584d51d8d010961d3a51827dbb2a5ed40b98d5a7e7d68442c77f47217dd213bab22ab0f8808d57484b7a9e28975d44735dc460527230655c3c050a050db173fd3c6cbd5edc4ed5c239f4636de63cad76f67217ff7d124264f25ef7951eaf19d1c4e68822cd0ec91d05b26eaff5e577e792e81c18ca8613d0de6df399450b878e9711b0054cb820ff48bd712e130d1444b92389b01b24aa7906c27bf0175285905b53e780ffbb1b1aa135fc9c06f1205c356ecaa7d48c9a1d0c71b7565edd30da4d33a0365f57940d1be554d651d2554194f2f18561f90a8d06533d031e11814a00da2fe3c09fa38d2a4733f0212cb6ad5e41ae3186892d173fcecd517be7c850d31168705de64bbcbfccf1db1ba56cb7234b544c28c2d4833a979e6a256fcb43fc2d7df46fc948eb9cf4a1bbec8cb10bca8037a2763edfb3e830da2c71276499a5c2775c66042c9fe5392965298ff083351cd4735c29f6c8a88f38df2611a8e650530461db2f2ba76fefbf4d895ddf8e35a449766a17b90496367493c2c7081ae8ff726e69fb7e53bd25dfc9735683ff9848aa61a8952163329848846c67b183056d98a567c9c49fdbd95793a201bde3ac0581d7f5b539df6851af92872ee95843b961b90815e4cfd126a0e2d8e6665104f750e0a297ca5496378b36f0af86ef907265e328e02b05840d31f0e739716c379c9595a5c32d666342d36dd83afd8c7450b051bb1730820aaf6e3bf6f8bff81407a71daf1f7a4115ee95fc1cc1f722f417ae2dc7d04db520b4dcfc1d4b540fdb176b128ef6ec6fe8b05a91b6d3b559afabb79da0dcf0766ce9767b0912ebc97347c9ec5766bc85a320d4b545ad99a126dbed1770e4f61c67d05b311e1839dfef27dfb8e38a6d217fedc5e4b18e96d4d278ceca436b0d284ebc4c762c113494953edce0aa9369a6ed09d5adee01b61b66e5e2833b11b0f0b18baf026ae039a69a33898a3d85d613be89aa7fa4dc88fe7f6d0b2dbfee6aeaea310740919ce154c4eec59fa2b76a19a0dcbfcdaa24b1a14e598a5076feb28c9555879d626cbd2b6724b2fac1eded5355edee32ec0d7c8c78f625e69afc1bf85618f768f24e9bd7c42d617db2ba92efb4e2684807c8ce5456b41e8728540749168db63bec6f29096b88e793b21eab32f952fd3e54cc4813ba050ae04ab14788a3f4db6867d3d9edaeab6089f3c237e54ad1c0c2bcc0a7a9b3ab79db34e9ba4129c041f025c8b77601228ad26e5a10a7aaf3873c48f2ea80f71f4fec0f1b20eea92eb1072df185c06873519d3b4e0f302ea503c0126c58f870f34aedf97b61b355e37a00c1efcaf0f9a9b5ffe82059eb5de53f9e9aecf9309d3f420054bdffe01a60297f0038e5e5b925922bfdd92562e83e2d4e11b1c40a0db73229a2ac2cd948390575dffe06522168cbb4b4b08ae002972d8b6b4ce1c28cd3051b6af934a0ae3084ff95dff03d72b58454e8d591354c6225fcddd659d55f1eb89adda20171a5d09f0c5ae739170e13cc85c09f4f09e62d35947e3814bb6d52e468b29937cd083ac920c91efc729059fe53b8f7e45a1969f0003375458ca863ed8dbb08a0de38540429d9b80f010efe9f23fcae2490a98dd9e04f268af0e498ae1cc3ede8c8396b57f5b8e3760aa25620ae6f951b34c5f3fa144fee07a720a8289de708aedec9707ccae23fba436d14403bf812722bbaa034c962667daaf02feff655c14dd16409b936cd922d35c5771397e9154c4587b31153ec98b0d6287e40d1d1746afe7b69a3f98e18096976109dbdb947e6a837be3a9dd307fe3bf943e735f9866976d8f4255434d56f411c40538468b06d2b5c0870c55a0d6450fadabe6253ab2b27c4a38708a9c696ab88fc0591028ac24bd185aafba8b7a941972c1c9d3ad4ca7b2496836409b54e76f910d270c331c74aaff613389d396c68046a90a108cc2cc126d4c819be77066d6ad544a41e76f5f6538c117cc8dbf22903f723f84b73e4be19cd14e4f370282dc97c22d66b889ffbbbadb56c8e3a8c189c714b7b23da7f475d316941a9870731898a7f97ad206edafdb2b2479f4fa4cbd0324206d907a041aa0cdf2f632ab083d37d0dfc3ad5c2ba5d7c3a199770d8964de177d21e1907ab775a4af41dad0e6018d4b7699c5440887ee2d6e01c824ad5927931b4d5c2ff7cbe0f8dca3a19d41e7d24806c2597a749239da2cc560957ccb4c855a1cdf3970b30463fda1660678c459d201151d483238cfd1f890c997464407ad6805911d7065555377aeb5ee0cd5f5fe060b1fcffacff8c71ee3c03f592a41a62d9580050da8161a8ca3b644faeaffff43a677a4b5f238e98b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he0ecadea8883e995eed729fa705028fb7c1d203c83041e6057295f69f795e9f5a7a78086759856b87299a2ed90d30f96f9ae952a53c68ddc02bf1e70e0e7e7789d0f96ed5a588fd7ba7c70362bbe8e604dd2c7518f49ec84c91f42581b039ffed9a305a69c080c834db0adf19d0becc2142cb4f2e2a26a2a2b619ef5958400c8eacf18597d1f64da3f7435b60c4688bab9d5ea4e2b9364a658ec71101bde67d78788d7b356088882a43cf470fa4a9a03201f7b683d3ab5d6377320235d2f905d08135fafa28ddcdae68db15ae180b110a94ccb2c40d25394f2c5692ce0e9dbfdf91953080fb45d5b23548f112332a7fcb0d3505c5896864103450859d39d4b49cbe4cbae7012708396c5a9b668e764fe7a1536fa4292e33f96751d41b9d95785a44ce51744c6a0c560592ced359bd73679811e29a8f1bd4cd3b518dd635d5ed66fe06ec396fca5c5cb290a8537abab438d3ed2a56902b781d39a3d312e7fc0f7eb59320e13c567f9ddaad988c1174869dda66ddebe21a365d4a4978bc84f3d7ba85a80a4eab59e1d313d5f001860dc1ce8c162f77745548e280b3e1fb16fa69d770c4ccf05894c1c0283d41d2a6899ce84446dae738239295104711015f227bad2c6fac133ba7159eab9abc547dd209c95ab78af52f438a9be04eeac69afe8886ec7208a84003ef1db9ea56c35179859174d8a46db089d4b5530d6da3972a476980eb6b8930515fb7f77a33460ac5031d434a854d7ded7b3c512c93d0055e77c8ead302ee466ff57bddfdb275a093a837baa6d6311be32cca63f691007ab5cbf1a48403493810a5232d61424dc792b3da33eeff4cf6a59e17fe00e01ab1b68bee1a19901ee87ad72d0e106b76e78b8f650fb8f0672fd6059adbe4b37d037e600a86d39d35dcdf0c1c24400b6c06752d0e04ba4f060d1ed8cf664abdac5ebcc5593dcf87c1635332d630b411ae6f0ceda768d86f9a19d3e417353a79cd73249e60cf0d6110d278fa44c4fe0baaa01e68937be91bd49b7109bae28ff2e80604d54fbcf86ec90a2b5cb51e550e06836555f9cebfc1bb090597b4b27debfb6c67ad8cec31b6922cb2a7f54043af914931df5486e5fff1e2a57e6c0b051e9292fd537dd6c399a5956245f1e98b99a8abb36f074c0463e40fc81a1e4ab2ad51c5502e497ec00ac2515274279e05d56957ef7e1bf94e9659e89381601ed083aa75a587d5933bf8ee8261a39b979e3d90f1effe3ef680154b02355522496f82c5673369912c2ea1dafbb3f8e1042c0396eb45ec3468f54cd1a9a52b9355b6ca43775b1ec3f82ecdc0ddf28d8d5981fcc5309c06dbb772753f29e08cc2f258d51a3c240f13c77a132869706d92d20e9c1c8d4fb911922caae9836780f1179a8ca28daf449f1d2a197c65f1e7160f30bf77e8af66e5457fe76d62c69dee3046970a06b50ed386f32abd68f2d5ddb9b48f76d6db2556ad3043378afd70359838461d3cde83daee0c9df84c8f96d88d6b126f6fa97447a41f0f6553fb9d85d83a074953201820ccbbf711eeba8511875a768a96cd82f5a91de232bd03d1335b3dcd34b798f556442e99848b7ce134d673fcb5dab067ede4b3c1fd038137e76493f6c9dca4fb10491efd1c228cb747936e04a87a70273617a7ed1e3ae259475b6d841f8cda75b57a4c17cc46e0678f0f6c9bda060095c4b2adf27b45fba3c9f1713535df5df7300d3d86a657bb1f23e2c4c96ec2f400958f2119c3db8334cb8e3246dbb7136f747a1bd3415ccc5b850edbeedef5b7dfd58aca81b173628f8b5d994b82022f1caea5f09a9010dfea4bce14aed079f15e25abe4df74c9ff085c4816656274ab6c382ea3c6f9f0f334e08ae97eaeac4bcc98ff874cf73796b5179651414ee3080474c92c906a45eaf4c4c54b59733041bba476b2113c9a7f7b6c0824a09d41821271c8b6a3633226d1fecc307a1e630ae5388724d672d8957e392f484620857c52824cbb47249d9d243c4ad65f646812c9c3942228ed82a2c9422af69fd0a2d1e3cf31b46eb2352994b7f15c72d88bbf908ca683c7dfb539bcc62598aee7517302df2a1122070b6319729d927118067362437cdbb18bcc07f9b29ec2f8ba93d68c98e483485034e4665572c9fb1e3162a1d7ce0aba07fe5de14b2b96711c34f35316005a8aa476c57402f50df5d00554624f1b8d3a950c67833d2540d5fb9458799583cc90c72a3669984e27d519b3f3b182455beb21fc5ae92830ab747397543fa9c05a8eaa703656233444c19f8a361b5805f34a7ba2adcd85f957da1c806bc4b7eba5aa74414c5253e8916d10e71deeac886860be2330cf7a4653954e77711e773badc3a72963bf6d7205b5f2fba3d90e7c7e46a15ab0b46c7de567916e728c156b202c3cbda1afeccba7f0a80991e84d1aa82e76c0b63c8763f98e702b169b3c5a2c6bb6b3df455e33ac9c656954d2d97881e9316ab63430a4fef6dfdf78f0b79d653d04f6fb3dc4375c7f58de61d0afb898e34ed52fa6e1c3de4d246c795cdc74cad1e8e31a6b4e8ef521aea47fbf555c1a27f220d2691d8e049e885615f836478a049b0cc159493eb85cac96b8b4f94f008ffdb820433172e389847655e61f19e134cfb5c4d0943d69c1b5742a4f939fba206bb205cc26a53e5521201183effab9e20fa790781008021048ebdbb527000e96415193775e87422dcbd04d3aec4169573a826a5d2b4966cc19e81a76d8ef7312215638fda2611c294b207ba1f128f6b7ee5db51fc06ce396dafc7d586c70407fed57d916e791e991ff54aca46873f657194d24ac4941306b399ec8379f94428ff9436d7a6e7e57e8e30cd6dea1a1cf4ca88fd5ecce0c2290b015f5ff937266077567fc75df444ebb52f41dc14fae05a1beee864d1ca2620da2d9e3af312c7e7523c19528ca53ef13cb2ff2bbb13835527e8ffee241a2ae59acab24441797ffadf0b8f7710cdc396c6492fffbbf115c31f9f0b2b4d3de311dc51755ebbe03a24833e3d5338ad5835c905b9a504250f38443e8dd3ae261f2056be87b39d01081f3e37ff5a7f2155346a56ecde2ca75d74dd13c99cfc046f4ebbd1d207c7858f3d7aa07f58979e79956b509d55458fbfc3c1be0dd88553616a6fd3fa7609b3316b06265871df5811cee654bccc08d93dfd012fcf27ba8bcfe24594887e05e1b0dfca4ef1886259375d2172d7b5759c8ddc33946ba6ba404dc0bca3a9920478bad8897a4c4260419070a6d718592785e4d2095f11b33bb6c3a8c55a879624ae858650e8d36ed329ef27b85e660d80e06d5d2b03e2c13b4f1165c5fd0daf1670f7d673332d720c9f597b32c9e3f38f36b696000cf2ab56a08238597ac5f70fb01ce638767cb06a979f1ca08b862c122f658210a70bb4e42f58e5145202a56f290a2fbf361a3a4ff3adeb01f20dba6ae82b1eb9ec0ee127803622284e10d8646082340660a6160a1c1760ece528ce0a427bab77f913ee86cec8dfa583032f4f9e4f99ac0da4041b0ce74657277f93a13dc349c6e739867d538e27d9bfcf23e74332d16491c0eee93c3148789b281d4a32ded817031f3487fe203c6e127ea10ccdf33c6b9f15141160e6ab28b77fb4d89dc5ccad45ed58bfbf60e4ee4f2e1dfe44b685c60a58c4e5f3c63b89d2118280f44a3dc5f1b2526e8538c7be40d18828b75ba0a172bc351a45d57d97e1e2aca32015bba3dd4512d753d48da160473be8c5c4eba9008a6dd95d142330f52eaf1de857dd4bb93a251f5ea552b0ffdeb13461df2d53db9641de63b5d438ea553eaa8b52a1a922260fa614a8ff3535b96795f3fa113cd337040ab92e02735e4eb527552404be8a0eb0f84efdc2234ab810f8a15da7661e5ef068746c545a050bfdd806dc1da7fb2c0728acaa546e5e03e62f27164d58a0bc0c51fa2eb6ff002d9a0ac58733c1ccdac7049498593881dc106b5d0ea31f8332d2669b1d576deea1fd48d9e0805e2c5d895ffa5efcfdcf7fa1dc166dfd33ae56c2be1c4a7eef8f82cd060b9b8096104cb32f047803c995f99215130b2864f49644afcb57bd3d6fda360ab77f3a0f490e798ab5954581d73128e1151424d0aa38fb2f8fe3fde5a985f489ea2cc59462300f7a5fc7bcc34a8d8cca43db84a1e1cbf466bdbe04f41eec5d3f6fe8fb8718df7ccd064bb6844e6660d01bbe84efdf84ef87a938a738d09b8d6f497d1a584e25871c7d3037ca786827cb4ef9143f9110008343199e289df97ff1858afaaa22aad4578b9d5bed7c8a95ed9aa09c690bf233304a746c1ea508f896f476e65c9904ccd186fec7df24aed5683ce0946e405108cc6521a83fa077f1b912a28e09bf6285acf17f7fea172854a3bc9b9e6d26710f90f88acf35182833faea30b59be9ccdd2515c6e44ddcd4b39269ce287bdcb55a39bbcaa37bea5f8b76b9cdac8a7b776405580340948d26631d7174722ba11ee1b002d6632a3a2cb7a12db4e97064d4a050c05692d327debe1ec5bd4b74f1db39a2139a9fa30fa7a608668a938a601460f385d1a46f45cb4e5168d0ee4b1a288782a59f198b8f63639814e0072bb2694c4d469b578b02d77d029f182442bc8358eb1015ee6b7ec362edb93f82e3466e8233f6d77b18567e4c265a417804b0bf9527f63743bce758ba10b67f279185215e25e60b29ee1d02f2624cf375b5c7992aad69678aab945885a8599b2d18d6203d8703063e4174b002c01b9950d790773691cef97db83ed872465b4dd51f0f39402631de4a048b9ece91ca69ea35005d3a66d59fe0bdf2454910bd1b82190cc60fd53561a1379d9b029ef94acfd178491cab3be8b5f81af978ffbf564b8cc80f98e2eb84720a5962a8343a407810b032e712e7d39babec6c0717dc9921afb7246cdc5b38188b2fbc90cd9ce473ba479b31f0277f6c69529404183ead38afa1a8931bf3f634f423beaf76f9200e9ca3e89d3ddbbfb4da97d2c71d5ed7816426e0900cbb7193725bc2fcd1feb50347e55fc7412973d27cb3ed67c827adb52b2160441cf6eec47ea05468f14a4a0852e5e368b0616d8cbad9dec5f51458d58f6a2f04a547529bc1d5205e6624244b4efaf52c2598638ff9e05d44daae13c80582158c25b67c71ec966a371bd6c582858441a8a8ffb85a4fa19b77257842b7ab0d542e5cf88fa0f12953a151890203b1480083efd6b2b9dd34113175eae1feff9cc6b7c4bba6b69f4be6cbc34c7432ffd0d4dd079727229df7f6c31f59c0bc217c388adba716fbffd0a9b9befa4de64b30629bbbe715c3a3a6cbcb61124f88fd71b4d7d20c3ce7a68dc1882d3878556026f7e9afd4ad3b6ef2715714482b2d77edf4c84675a9a00b28ef675ccc5cbc8ef1790cbe82b262721f7699998f4925ce1d2237cabf176be2bdcf21de469a4ab6a7c706ea38a562c05212f41c8587f809b6620fa1aa5762a8b152f4d49fee11e49ec8be326c067b0ea54f7c2617153ba401dbc1209da950d1ff6dc17d73985117b46966497134d0dd6c8b423a862b599075454436c1b509807309515f08b457716f9c28de4bbd16113611a174146d80aa739bfbb84e24bd9f285384348ad90dcfc99337d27869962b1568daa429e1c4f373098fe602ca24c7454c1af19dfe94a8c5fd92d3a51852ddd04ae2701b9168e059cb5e14a3719039c2ddc6468ae7b2840be13ace8c246f8704843c36e760d523e65445d2581feea434055c1c99e1e2ae5f54aed66b67a9f5c1c47a7a5e9395b8c9521fe3937cacada8fc280cee0ed63a4ea31256680efe396e0b67fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf9abfbaef9643993af422f46ab0ba6f59a9b1a2a640711b627d516e91a8cdafefd70588762fd23abd83d22bf1a61b13eecb04fb30eab1a9a1f5b51d7a04484aeca963a6736cebaa38b167fac7398141a274f661ee7074da401f27b6d39758b0dbb3bbd2bdc1bc40395bef8f9f62cedc1439d4130d966f8b673b75622be4e485d9ce1d69ad0e38cb87f76365605f9ee9b5acd837be7593ac68a4294c6475a3cd37d84841c76063f8d66c1a12054069b3175ff83cb5cbc2d663b085e01e16b9f1fcd79015ea1ffb600b2110ab6efea4bbb6c24b6f6f4fb9977d9daf29ad726e63c85b59e3b51cdbd7572c7586755a775a6e8f7e8b4a06006281a2ef00f7bdcc2aa73eb054276ee7b10ab83b6fa919657b8b3738d19cbb722f9d1583bbb67dc49b1a50ddf7fa72d6eea542089e4f428dfad6594146f9bdfdf32e81676bbc93f8f61032c4a609fa83915b80ad945e43cdff60f5d6603c1a9f09709d0e2cf94e99b77541ab72a7338f120c1d17476e5949c7ba0f9a95370beccbc5303b614e8fd13f3d8be718ba2d86e71562d9b7501a2546137ebf80d1c8d7bb45b26256d2d350b3b9e715e6e7c6df3fbacf33c85b10ec4f539058f84d9cafddc5c51824faafac4e119a765d0875b041e8cc9f5862cd978693b67b39616370df6b6b94e9c6683a1e1e54b49d45a3aebb9501a6357822ecf78a34b9a868ff6ebb114bb341a0ae649c7e02e06085043e5d466e60670bb609dc16d3de99ec9eb576719415c02ec2ca877a91d636b66b11890a2ad64c63eee94398256c29bf6b0863a2635fe826b0738e33505f66464fe56fd2d5fa9842f04ddab59f31b4a482662fdbbb2186cf46d615cabbb46aa282f1263992f05be69311cbec8daab94a8b82577cf24e5f1c898db96035f09028c3243495b112887848f671eff79227b3c2ad8fd150e698888d98d0f09fdf3f676710b37ffbccec80db44d82244eb1dcc9c67b96dfdffa649dabe75c4ae8c8c547e86ef7c0477f1fbbe0f08e95c7d9ea27b27bbfedd2a9ac9630e759fdf991b6ae67cb7a3562f8df42199c22b3927b551de75eca1155487dc2362bcd37327f6a9024fbdebc007b7b21fa02bbac902e73c3e65e2bd3d0d6ed60dacdf98e0362c9321864179c14352febc78039408d3337dabdcaea2e65ccf9d627162e73200ed383f3d42b81aa9d2cac89805c292bb78c73af642ba5bf09ece6e38d13f5ed7a95f90b984a3b5a2602fdc1a7d800028b4e7bd74c353f0b1cc205518e305f7bac0fdead5fdfd9ee79a68cdd9f64718517b374a12b54ba7492bf6475eb4dafb5d782f4ca07872de41538c6d74a08d1574a4673ed2b6fd83ddab0ebcd079ce58647a5224855661ec416205958be1660ecb593dd5aee03b76f983b2e7374dbbb675b46f2e899c7ab27a1a70d961e16203c48f02ae0f66db9a630897bb1e06b30fb151253f35bfe34d8f50f8e796c616c981c312485a701bea68b23803208bdcd7db1629da6dfad588de0bbd27824e5740a4af32976e551e964343da86363a423d8412fd9f62f5547955153d8f357fc54d476f8b9ab2f0c9617b21ef0c003711ee10f3923d609cad3d1c7b58e20872b40cc448b36453bcae1400951a93b757bbef940ac3b2dfbd6bc7d704c2275f3fe8f0151c063ad4b67d608c55f13bacbb50f4329bfc51147db5b154506c18cc1b2d0203589d9a63350fc60befd1c0b7a4d7de3509ce1dccb256cba974eddf045e334757ee6cf1aeab39e6337dfc45ef1695b647720283551744174b1a29ec22a3879be8c62249b67d570afa14af761d6e2db06ba3afdaf13d62794c1551a70514a2363101f0cbabb596732a4b393c60de0976f5a76058594b75737d62c4f78f0b7d648a1d47a438788e68d0176b9c5d8458a5d83af3ec82578f1efd28518d6bc6dd7065a1d85029e470b95c92112fe16cede004f511437abf62e4bb68289585f8af686e80e326e9304d2b181d07f4f10c42723c6aa0b71733689ed6ca7208a901d47dd87246ad317bdd0af2fc53bf3913ee6dc8038c6bfc5438de59bf4dfa43f1af372426e7b44e4e318a7ad257b86f2f3c45e38e8f21294ce88aeb301af9342bedb565e41c1c96b2ef229a43e75713e8b057590eccc1cca0e529cef004683fd5f8d6fa0adeb63660388fc10cb0441a62b5e2b4cf1bd7cb775b2e05a221ebd78c05e3572546690c8b2f5d914acde5597de6be86912f691a853d5e264ffcc04ca9598ab23ee636f636f138f15093f3a76b96ec18f65bca168a8ac7382af312b8e33c2a2d283c10cefb3e2c8ada7774bf0381f8b1c5b1177b6ae6179b0d054981515133e4bbceb4c9f3a7a43681bf658afb069fe9d1f39c0bdac7a1bcdd24337df186149b0ebe92fe4b9f1a19d2e7c6bf9765e4732a45a4cae43cd482ff52b0ac6645b893c9e87f9ab03673f39a41b06a716a0692bad24989b7a7b49b803ab7bca3008cce6025dbeeb123c1795720c4921d309b09cbb3040d6680d5561233c0d0bbe749a0aca7f4fd5f6e3493344956d2a31df3e001ef1372b576d4493b8d5d4b43b3e3d441079f7f1e3258c8b156741399cda49afacab2d9c773d8223bde64754457e9fd0e0cfa4ffefa9b0817422603cb9d5b7035c5eb34e8c69552501fbc8b921c9f3053fc771d1ad5b88ddb7ffc8e5e95a4c4b3e5d573aaffff8cfa594d228d380573389e322cea184092aca544e009e8f7e8d5b22b2aaf7c1f2b0b6bcf92baeb4ad1c97a4ff6eed16bcf471af83506548c0f2ef51e5791d76dc8d4086dabf02ddd92a635542aa9d9682d773db78ffdfd327a08ea967c999fceace5d41e1ccd5a0850bb847944d39a6e6a85839002ab31c23f3ede1583dc33f4808f7f9ae305ff5bf08b3d08b1a7b08d6aa5eb9a165681c18f0db02ff081ba20081ab17a9781a52d7313d224d424470c14e542e8da6b79cac2121e0b7fdc0ee0f27b9a7f10649988938cdb8f4fc1cc2d357be7674ffbef297c71328951f8788ebe2c86b0b8b2e3985106a4c3393d420f2e67d082d5c7c45975521553313eb855af54d1a2acf74877fc540fa3894621609e70be1c80fcd844ab8de2315d0a5fe67c04b1e86702a663a2bf03a36d0292e5e055ee6089f9b08cde7f4dfce6398ee36ab07ad9b8309339f75cffd957021ec74b5aa1690ebd05730a03ca0a5858a68e24ab7b90895f5f015846dc62e88387645380f8a9e8b71bc180c84c2c8fac89724af7989ad96f9d0a75e48f24dd32430269b912445fec51c643acd9f7f9ec4b2b5c4acc1b335245c5955bcf2f535d928032cae0c5d5669cf765efb9086ad21142f45f7453de245165b9c26860d602c1683492bd187fa4128b259a86084dc0868d4059837cdc15f77fd06dd7dc6beca41fd9bf83cb728dc59ac314f718f15e2ee26bed11367b0f9f6044daea65316e4ab6a1c393dfbc92318f36f8c4d50470a0d15894a778b3c88fdd3b41e3639ca18c99e100d543ceb28650733331aa4f8d76adecf70648a6033a4a08306ab25a4c5a58143e951b99753349a0d97670ff585d71ec4ed35d5484ce7ea6bd889964037ee6ac4306f18410a06d208ba75907b2cd4741aae4ffa709f3b895219d55130adc23b60d26a08ba14f248b163a0267b629097469ccdd1fbf2d98ecf16f0da8b7c29be2c132f4d847eae31b6f913e9e6eed2b860e9da9a5b154fbdff696cf73ab4a4bb6541dbc993c96ef614801d2d239c962058d764e0f9d99072ecd44ede1c9304d4cc1c7cbb0ba3b857df7de0916c8e72c54c988d86e6e3aaa85d0be622c1dfc8bced5b5be3126b347144783f10116c1566737fe460c5f63a4d9f82f328877f6e2989f12cea4dd0de8e15cc934fabdab58044fce98199999797e633c9ca2cc127fa66f18624dc2ccd043196f14b317e038a65f1afb86cd2d816b9729657c6e3f0a55930e87d3fd621f946ac23dd6a5db355cbc3aede0a3d30cdc1f0efedaca2d5241d548f88638adcceed3b4b467c340085575d543df4da101c251c994ef0c4d37cb9bbd162a80326aa956c4c7437ff541fbd6b62757c206b68ca0a35d1f8a69dbf9d16b2ce7e5796c5fa230031070de0f4fb4318ba3ef1b4ca11469d867a96d730c270becd01048c9f13f909f53e3fd7721509392490ab4dab375570d772963baa2ea8b763ff1a010de7f91f83841475c014d47d097b3e4cf73b7a47d5c3e6d914ede7766c5d2fb3f3865e2d3073c399f098624b18c85357b031b05c2d2f25e44090548586368b42da4d196d7afede5f6d3535c4dd1b83aece638454209167ccc576c0c7bce9d0d7ac40f7e3deec5a1eececa7f5b83956b331a19ff32d20525e7f798f60b3c7d2dc262ba542648b94f2f7189357a029ab5b47155b6722ecc90e30cfde7bff24893dcfa24f77b2c93175ec77f6268e6d91d5d7dc224341fde7431c67016a192e60c116a3fc34a70202431aac089173b5806488a98e54e4bc526caa3fc4cc6ebaa08c3aeed0b7252bef41f22f76d8526e77f449b5768f98c7d36510cbcfcb84806c9fd33f395a99cd5a77c268b7136fb4ab96ab7f6d95e4ceaea23c27b87e7939e9b7d7e2d503a5a9a78fec1f37a0f4d300f4a5d38f08a86e50f1acdf50120aee777657fa5a01c31c6206155583eb4947a49767b20409139dc55f9e8e24ecc94bec50bef8f527fe08c3ac333dcb9dc561f7263867f80ab290d45f9b6f0a8bf0d584e8cb9aed77514730ffd0d4e61743b85f10c95b9db3b6c18969528dfdd8e5000d684399592dcbbf11ae4f376e857c6a048866793bb3955d43dd15524c8f472efc488e3e7420d18b3307e1bfa166e6d485f0a720adc4ecbe07a880fd29a86b326c409d0942b5f429e0cb0fb289ee9bfed1ce8372f932001fad64fea6494d3f72617b84f88fc4ec51696f004cea0959bda242d282d6ebc873d5ae1f2dbfc606b9f0d82c59daeaec43348f1356a15105af373dfc7add8793639223d95e7f6ebbfb44b531092392e530ee6ad8a4e7f84055b558e79355383e1441d658648826315a0c870bbbe1725e5f3d4bc97fa2a8b1e74daaab74ae67d4012fbf1a66e25f374d2565165da636ef3c7c132c069af615ea6b5ae7febff86673970bd7712ec34a0c399c342dcbb8ad8c9a67f4c86da382af9092b925a25c2926d2a4babc010145a407c192e35dee7490144c3ca112f15d927f2c542298fa4a64f2aeeb6cf93a6edf2f15e7c60ba576ab8ab0755aaba99b4f226099ee385d9a9f7abf396d35333edbccf54b3ee026bdcb4da75fcaea342fbd81e4cfb2514c13bdd7d48cfce9c19880faa914d49a9dbdc1dbfe63601bdfdbce133b095bbce5d07276cc54f2443dd6ea0787bc5fe883501cfc91c20d4ed6ed9207f3ea379ad389f6cae4f8321b22180611214f2baf7b6645808fd5415a9482e3c51f79d51d9da01c9726021c6474742382e30edc151c5a608c8931dfc01a3b801b644642897ce4a64537d21e65e78d6265ca9c4280059e87a8f86ac9814f38ac383fbb8078d0bdacf2b07493a3687fa44b9670039d3e2838faace7479ab77ae0978df4482378aab2646614fe6bc2a5c7b023f08a44a8049956bd56dfa5332e9cfccc38b171bde25032bf4bf3ac05b1584b3e146246f2204c2b58218a338ab13e75a1f2a88cd39da78d1205429f846718a9f1846f3eed09e1ecce78fc34ce05f0451eda86e1c49535e330cc66da8fb0464f94e92028b0782594d1656c4040aabec5bcf8da642b58668d182e65139aaf294a91ca0241cdb2e4e8acd7940fb8fd5acd740a6a899d8e1728ba85e79a40255b50;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h774c12359222f720141b89e854c1821a790ba3094a86d2bfb27b70a9461b6d3c06f9bb98dd6a5fb38067c3a79cd754954051be57ab5adc273daae13f7513bd378d45189b4d0581b354309c57eab5804365a3b5c2ac6d036ab23da8f6c3c76612d72ad4920d026aabbe18ffc5cf8b5e7f6144e839f6ee3a7f6bc4d53868f02ef9ac5b00dd08a66f4e49bbd6c0d5fff2d97b89e027946b6594b20cc5b4a0ecd148422d1ce55887359169b51f0a9d8837496ce8902a46a0be1d5313b27f2fd4e8bef2436f5db885e4e274dca444c4e447ca95a8ca3cd66451cdaac3868d6dab5403ceb21101c462b8376f6f60fa048bcd80f01dcdb04074362a5a28db5cc10f9bf3c053d53f2ea4a9e397a911ac86c75ec2a47d6a3a465efe572253ab57c33e9f9f150922bcb1190937bd26380412fa02e1f6cb2732e824d6404a8bbd342e1e9f4f842dba9e6b9bdd9ef4ba5eb53a1d38e2632afb2b0998d5415e3464dd64b4015666081e3730d9a6a362c17eb83a446223c49cc60f49e650999e697b9dce2a26e71f160f0892c16ed486ede974825553b9141f6586b14d9c699b6da227bd16f5b8e41bdf3a0d11b134fb7a004518437f8d6909c426b30e60e71c422bbe4399315ff9b30137a32c4b1069cc29c260b7952ab1a173e0893f75a7fd3e149ac3343727ed4941113dc5b65c5ab3b96e3b7ce2b18133b6a1caedbf37c55b6c67f660d55beb18dd5f37a91b5f5d9e6d83924a0f0ba0fb1246b5d509658aa0c120b06f4d9cf4334a7d6aaec93436991364d80d96127bf49f0b1ccc0cabd08e4d93ec3534d26cf8ffec5578499daedbfb9d396b397e25bd15294b412b477a933c3dd0fa4fac11d13aae2a87ed7469d3aecb5a23960450d03720f644e67bcb202b2be4599bbf50ffb513007cc6dd919f0034800e9b10009b00492681c4f4791166b1aab5879fc4afa974a95382f1c4062fbec3be6b7f8f68cffd88abcfa5035a601d14a96c3b030e0303c13cba79aec52c7ae0f6c8079e3a74ca9353861031e70b6b66b6d2a285ab8ed241211f7a0ada6d331c9f3a3d4a43baac2ef5a19473a596b9767cd10cd1dec63e450764513403576cdf1957831672b779b079d350ffd01579db50fa49b7e108848a32f261abac8fbd2670b965063e6acc2d557cafc2a7fc121764e5f04dfdcd376bf4a7b8e8b0c8d40032b752caf8e7a8e31a68baae4650ce46effd3ded6c6015d0a36807cf5997aef16d2d6a0196e237fa2f435152d5ecef3ea95e5cdb318d61116030d4ef513a27cebeb95b3174eade1b34c4df6e3f6f7cd7b69e1ec3c69738cbb879362d95c57b93851c13921f0c358ea5399f90e9e417620efc29769cb13b02878a9419b115906e367b48554964ed6677173ac5c881f7af20b315e7693ce7abe843106b796b6205ce4bbd4200be621168f0aca3c8c0cbb77b5dbb031f8add8427b76425f88a765f8b62da1fd721466945b37c950648eec38f107b5e15b90ba7d40246a7fc1aa7f18d5964d9a9d0cc871daedb2131a167ad2b5e71c62e260c90bf81c161e18e2f820d842afa30a1e4a718c2dc3e6c96c7ea424c7ac388937129c55655500bdfd29a69a8d59cdf5d285e77862c528296cde03be3d92f5f7b421ac715eb7e08e6577c47307525eb5229e3ca8f2a00eb02d8882fc14534227b5fda1e30cdc2814ea1aee71aa1d5bcaa74ede382fa9e6e4169111576b55a66134afa002789dfaa334fdae5f12ac72f5105a1821e1dcd12671da45710b9aa5f700054b59d3c9d83979446e5d6ae0612d6e2da509506c9b2378a76aa1e04f364f358569ead0d7a2206758b40caa0e61e751daaffc7ee918c2e9475f392e28227d64ba26be0f2f0f7af6a2a9a520aa40f10da22147c442b821e5592135375a6c29d1bc7a16ad0a6fd0f9d6969b24d4508a3ff13926e37ae590f87a2573e78565c151962a99094e1e9a4ec0b17c8c4b8c4bc0902a3ab73b6925f613778630e3e03c84310fd85989729e145a68547e340bc07e72f5cad7eed8e8dbe0366445c95a621c2c0305fe7b4fcc768f7232eee1fbf4b3633afddbbaf1104f40fc09fcbe256376e866a9cc9427db00fb2ce4d83b2f9fd34f00cc906c00180da8761da443841462661a54f5fa84c20b1f7298b84194907257ac93693cabc343dbb858ddcde8eaa13c613078a287be58bce13ab5511168ca9619465fa5f49f7b94cfa98bfafbe02187e5f8420618c61b3bf4247958c0832675b51476ce6a2e85d933b023a441a3638b8514172a9284b2c1be7b0559db5d50e845e917af0b09be89a0d7758e3606d979fc642d7c06d2a3e0d35d4caf9dd70781354b99d96f2ed4aa0c7a1a42a9d1a09090d4b4406f4fd7a8e927cdbf81dceccb5c9700dfeffc2606bf9849eba1b2b9c9ce0a5650f35e3a5a675219f9491839a8a941d29e2567e2a973f86eb8a7226c899b0db99dd26c103528b027c9dfd48a834a43b36f9e16bebd92c540bd8d99991948ec5cc382de95fd098d61856ffd565073d7cdb994c3f009f489d7ab892fe6fccb43ed372654a702eb97ff8d2d510e8fb66e0d93bcb95a44da244007f0870f5e04603ef24b563d69943f6997f8eb4040dfeaa78b0a58dd9f76daf73c7bd762151dad9edf2ef4b3c0750ff38ef85887b1153762eee711afa7f827ab063e4853d0bcba7ad19a9e559cb0b86137e62b1f14aa5f4c45429cf8a5e16465f2e6c1ecd9520cc763a80c1fe9d42d9abf555a2a92b2aed1043b2c63244056e9758c7b7fad341f43d9fab9fa6d73cd28b78d9f2977d43ff22b453455fe087fc1e470f064c8ba10425839ed5c64246ce2fb299586ab537cc93082dbe4c500488127020fbb9efa05c4dad394352fd1653d89ea753e4a11bb151c0da12c230a9f68a3e9fa1926d95408e5349a60a1415ca8b45b6f5b3be3c4758c067db84aad2849ef07388fe1ce1b4c6b40f9fecd7af553b9bbbf4787e477908a4d241cd07dd0ed850b526dfa2fc2af6287ace191a602b48194f42d8b8b96fefd64eb68c0b856a6d7da1b7c9a099d75e9f05f559ab8911701b7670eec14e785ba87e8c9e5b6fb87f932f7e71865c19d667882e7d3ba13db3a255b95d89be5d0c08a6099cfaab9bb68c2e0743163c991089b0054f33b98cf8b016ea4535fdd193e032b20d5777cbd20d9cfa35b393defb8e48152e6c95e7d965374c19913daf4aeaefe0a6bc868f420f30551416d9ac5271ff47e87117a9f634cbcb7195d4ef2116bd8544c5717a80bfd193c384024b9ee4be48f1483672c52f8dc5088de36ab938a4183e90ce9cd9803654a11a26042c70ba7b2c87bb4fadc708b7652747d5261b37fc736c8a5a0fd542c3cf73445383a5090e6b1f4ba349db99d5ae56595d0175b5507a1ca97f876a0d3c012153ab662e1e263723104150935a45fd7e48738836f433f9ab766925f8a50fee998f5a47817d3c29197df99896d79ead38811b3d0bd377ceab82b7d6c39deb1346463f7cebd7c8d9c13f76f4c6e942fddc381523ca635c82d2544fa293a1862cddf13116f301a2f38295d6c6b926b2e7c1eb17b78b2de702cce9e692d2246f3fe14e20d106760c9445858ea049a72c21f33e948e424c1f9eba681384f6353296a9d7dd0c3c839364e5b0a282146017803b4dc6f594c6b08f441cb738d63a518fdee32cc1b364e482e9f3b3e785e9e0c6a8215ad20a4e471a7881b3d569f25d55e8ed81af645fc48480c5458bb47e928deb165cde4bff2d288bac1939074b997fb89fc150e4134b85778a29a7322f4eefe9d8eddc2312fafc561ef85c9307c784d9b3182cf00cabcf296ee2b10eb8acb2f2462631592e45abc7918a208c1bf566860164a0206fbd178a6c16da24400654f8970bbc0bce473919003a4c67d41155a8d9b78b3e5b862639bcc6aa5d8c54df5533575e5e4807a2803d8c517925009da9d65ff89fd4cfaf676bdaa88beb6b4f531a01eb1702af880861db07bce8b1c479365781e362c4a0df802969a4cb825240f327bef0660514a72e691ddb20be2eb1393d7aefccb95bbbec26e43391f726bc07cf5b0ee3eb8b26f692d425e4fe04191ed7fa1b0cae750284260da67b3ffcb0ff468577cc24a742d09e8758f128ef9992e851eaaac87b5a95548f3077f603eff046d0edb54cc911ed62e3f35bfc1a6559aa0096180638edcb2b2a8690ede9b326638df400106a53df36734f15b77d50b8859da8173cd2117b4da52812559ada4b1dbec75d425c3ba546de2311902d994d57c9cd9d496e7665faf14a5868e050b7efeb44c0b502c5962a4a5c356b00e3cc56c486fd9efd78570f1d3ea2e46e800fca44b9dcd87bd32bdd8f007cb01f9b332583196890b580c33584fc179ed581218305cdab82198ba1a3c0824c2c45d198f4c827827ccfb1d0e635dadee0823569581216bbc4c58f242933278ebfbf9d1a5c5faf35862e7c3a8140bcd9c5f12348efc4c49219f34be5e84cbf60ffca767800110a4e94cbbcd28a001614c2f4f38e0ab9b5d0ce1b8aeb20e366e238120551cc18df61013724e01706d82ab10f7732e9a47d5ef410ea7512711f643ca32f91e77e69447a1b7b4317101f23714736c3589f79c74dca9dff4f92d3580773e042a536908785155ef24f378242e72b88e6c08a81996b9fa04208ec4d074ff4b73fc2fa152bab47ccc140fe127049c0aa00029d4db5bfb8dd1857f8b6a6799ebfbfc521520b98183a3851b0497db6688326c43bb2c6e994c97e532d363d45e4aa95f0fcd6f724eb4ea258dd066828abed40130bf612a83be46cbe7f185d1527181ea973b41fcf50eca4506da07ab0c6fb3a2955454b9b42286ee41baf6433b4899916c6f1b46ffbd77c38f86cdf3bd4c4c7fbcf724f93487fd8cb976fea4325d8b677a02cabc8fe6feb3a37d1f5f13acceba11cb32c319600b98b7700c38c36f73d43ecbf81457c2a15cc74108e04702cb5e93067babf8b810ea881c43433aed4254d3ff8e6f8e669936a3da4f1b9620ea91baf48ee90805cab2dad125d98b3a371a409a9531bdf7e5720b49fb705cb10909afb7bd267d36efa53df59b8f53935a388e8eb1ee19ab9b6d31a03ba323919d6e115f017907bd680c22e2a9fd0e779e2f877b38d4e1477d44498b7e4d270ae3d1a832b5a53c8ab88ac46e5c75679bf8c6c75527e877e6d6c6b3b0dcb5c15087978a760909a66536b59465ef4059783d089c42f5dba06153476b758ed70dbf039adea4c9e6eda4919a2d214c83cb74f32f904fab95c2496467794c7f8b7559ca7d0ea7285fa4865ab397309e1dc3c62b711d43d045e6d4ac823b72374b11f8cdd186ad0f0eddf49f131c8ed4368878812773889dac7ef7b094f4f8ad84a1615de22355d6b7fa135bf535505a235b9ad9e8f90057aee960d971ec950707fa8daae32ecdb9d1eef747c5eb16d646f81a067d1571862e80c2ca59786cc19a303d7855f8a8a4ac266973ff6346aeb1cd2bc2c408ffead236c22dc38ed005ba4ddb8bec599b4317a038091e532525fa11c98cf76af4155526dad64340e2ca24db0df6927abc2bd17b2ed160614000d9a1ad6f59b6fbaf2061e0f998b9ceb703ec39cd88573e3163ff2f35b0a16cd2c14fce11c08db60f780e19b13d70b8691852b10a8cbfa47b795b55ea0b66d1aa19081c030457c015279d2ea47d71df7daec3af8a31ad6aafcfc3a67542ebaa86841a47fd962e6266bb9cda2c5ba97264ecdd7f8ee42a575e6c7a2f8cdcb399b5d07b6c9b4fc1608d8d5881f6de2ed892adf20cc9ae48a7dd72d7af083471b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1199798cc59ae6b7f85c39edda4f30b3432dc0181ade86bf92441bc74597acc926d6d7b829fa492b3d60fcdab2600f044e7ba7ab4de64462826890ea8c6baf5cabbefb8926fe0ca5ad44fc3cae3fe403aebdfe265bebdf10c5989a75e04af44b46af11d36f718365166adfb54c48447fed32cb538df03b80d07cdaaaccbc6c961f41f0b4982d9b919ad93019331b19f11edb0c1ca2db0f1ca0bb6bfe32574ce25b447c7c5a98787957d43c0034058bbc08f4bb3a8e0aef5d700b4d77dc27fd69081b29baf21818b3d3af3d8489b298388c69e5881921e2d7132f3b6387eef858b06bcb231f38ef71f0392c28254f47d3e2f5688049859458fe0781cec8733a91492718bb433090e44420024afa613979d1139bead7842139a513a7c31a839bfe6e028a655e9bd5c49b5edb100f154ab1887510226b8b57a5f7388eaafe649bf197bbcf9d02ae91e8a2427e5ff0c92b814190315a4d3678dfd38136d1affdd0e4e60c2d13677e93497bd9c2a79962edf71925f4b9ffb16ba128c98a8dd25eb21a3ba1060f7829af6c47a451ba316a89d209d61cb1e5b3da69a4076a6e99f3f156befc1accdce711a19b30ae21a7cbea465839b1ac495e4c778546aff90c71f548f1d04b2d1621e2666557dd177d76a55e60c190ec0b567f8e94378dc6f0bb95e65e940701183f695d9d973cbb93cd171465c123ea401dca0253f87a598f10fcb59ad2c89856afac67338322e16ea1e9719671faa319da454f15b6f53c2cd9f1609e465daf2e7fe29b83c3a7fc9a9a1a56674db759b3a7b50d545f76c844d3db70ec20db5d5a6924baa6ca1c837a69707a47773bd124726d5933beb5f226710529e6b3293327772e599736de1278692bc7bddc5c3a2bdc0a5d399ed4cd33cf86e2abf2a69d4d2099176d0e11f0772bf4ecbd609278cdcb5841889a8e6af90a2fe676fe0f4ae9aac778dec6d2e1be4c3517bcbb7809b5098aca8540f4b96ff329f8003864568b165ad0ba1c06a92a5baf3b2527efdeae1d35876e3abfe2a8c206e835784c86f924c202ff7da968507163e25cf857544c5db821676a1e1e0673fbd345ba0b3fca3636575e2b9416e9ef2f1930aa0446795cc5eeaa77a1590fe4d8eb483fc372a14194e613cb164735ea8d1a75e1a2b3c6df1374c1ba9f06521bc97efe1457963cea96adb671e75db36c11af90687732ffc3167d4773e9faf45aa8e14401654b29494676892bdb7eb6b9edab5f6517a3de3386899b726b24a7a73b017c796c2f9fa19d107c2f0499f5a9d547f663f5769a7ab39cf7914a84cd4b43ed90d2c19ec101300b08b9bd4bfefb0672c460b1a090bd28ae07f5a7146b8a602064bcf6d8a667765b78f8a0231437339e17a792b3ac3a3ddae3bd4fef8a2a729b251925da00c730a35594848928e98eba3dab669c95101bbcb022591a7c38ef2cf383e27eab80ef1e621c3d30ba338d5f24e798e1caed58581556a4d05679aa439d040a82040396b27bf76b0e1097209716f79883f55187fcb986dd51b3dc5240087432205034cfa2d715c64cda0c9ff31e635e89ed2c7998714aa54847975408e366ecb0458f5215fc47979dc176e777d3768d2d0eef50dc2c7874eba7adb6daad238dd07a0c37803d5fa3d890b2623ec0ed03c0a8a70bd54e4bfd5ee15db4200e23e68379bebb1766a39b068430d9de52473aa8a171a0cd8eb2ecce97b5dea5d6c3a2c6946ae017d878e21d5171c7c00eff44f9b6786119fc5ef8999f3fe973d3443b59ce131e464865ae3fec8ed1577997734bcfe8aca6846d2d182c85c2df1dee0df92c8b13797e74586c2b99c5a97834130896d8ef6c424e59f05ad09bfc98688994c590554f9c2c1efdf52f222a784ea23bd1d7d6525c5c5e0754410f2021cd970a767ef8f5af78c07b91c089e6fcdd14af1d6ba58b4dfaf863b26c05d24b620a162f2573854c34b27f5c0661b500e9b82a7608c170c17f893ac4b2759d059745feaaf35c5f13ae4b4e8bc9284dc9e431e8801fd374fafcf9812e3066cca958eb9a7d96a035a09ff61a1baa2a30ab85ebf7f58a6b00d2d66aaa2a239331542b2c86e0e67a06cc411be6ad554d6aca323bfb40b1ee7056e14a16aa93e9e3d37ee20c14fe576531e3a31ca6d0200786e83f145d37715e7eac3d79ed4bd5e417570d7807194539c051e22e7efd32c9c68f093e71b8d9d24ff5b719f9b45df72eca92c5b455c1c569177051209b10b6fd0f7524b941cf28e72a6a718e8c578d4cdecd1a8d942bee260c102dbdc543e5ade144b475ebcecde9dc0fe95be09fdc6f0d1c7eac87b794d1f18d0198dc3b3ab104ea2324f802ea32a889cb3486c777acaf2b8443ff30d042f348aa7faf24831c0e1ed46e1bdab751bd39586d2c0f5f3690eb66d0f5ce6b82433b40072cf537ac99e4b2624aeb2523bb8d9dfd6536f63f06c108e8a0aa3fde5ee9bad34568769cf6cefc6bbf35e7e05bdba59509405a1c08aff006e6396a205547d8a8ab19fd0be571c649d6bc745f93e885e3b492124811fe9988a7390f86d24a86ab2ab210cede41b93556ffde37530f684725e74483cf7480c5b890dd4c7a0afb9b9371fbee212037654c9e8a8f9d11932d6cbecab09f5f00cb4206ac84ce63a5ac9e6fdd214268ff0218299d0799fdd3b96c4e77f155807719cd86b287a32ae5d293ed3b3f8cfddaa3b6af9e25bf89bc324a392c8a54e7551c1cde48770ffb2184b2874347e32210855b6fab92b331aa8ba0e92fca6268504f6ab37dded0944972692346bbe85748b6bb7903a56f0abb21b0a16df7a9b5189cc995913a8b33ea13c239aad60e3a86e400593c66bf73bfe1b0d488274a0b93d8139ffaf332d401cb5b6e361046d009ead169f039ab5d176fad11ff583101a0adeaa500e048f8f7902cfaaff8ef8e81bbb974855e98bcab8285558eed7828b1f994d51a670c854cccd0e3314b066dee78d46fcb9be3f8db47d5159f264a07de04225320818702298a5a2ab19a3e4bf0232b53ab6fee7daec17fd380a94bbcce1f78cf08801bd490d11a3fb6f4be533544206a04220df7e3f31de99fc1073ba07ef624e8601d0f6b13537812e0f761c137a6aa6a589bb950ef61b61a51f13efcb0133e073711d309b94fe309e778177da978058cf8a71f1aa43b78bfe905349d949fa9c7fab5f97ef7a29871d7c7a7b6e6212f09af82bdf6a4b452a74e73dfd3175c78c893418b4c6aa8e3ff5d953e42e8658458a613b98e38fac36f4b6895d1cf9af1037b8929b41708c053aba7897ab6fbddaf07644e16cc6ee49a4d15b8b92fb50f65c5c9e92af468c71c28b5f3302e2f5043f70bb781c2169cef66d87b46d01a14cd1f346930063690a1f10eaf6f869c75a535d09ae1d0b377e7b574206c4359ed9d1347fee774124a0aaa367ae649c297ae1c7f41c210e7de95114c691a88fcd5868c39e7330bc7e92b7d5fa93343bca026c60d71d5b3636eb20fb4f0ee9d0c2197ea751483fcf720a85df9caf99f46c497f555e4f6d3a75c6739388b30ba01f3f16dccb9723a16454ef3c93624f522daf316272a083718e0d6511e998ea35d555024bff2c5e535d722ac2ed1c028de04c11398bb50de10ea7dd95431c68c6199eb4dde897cae37b83c7c83a74d939871f753789eb41862947af40b141d8703bbefb12a9335c2d889cc540698573e069296e8d9a7b853628e37feb225a9b0f7ffb69a4a9ee5c0b3ab43bc22d2dafa9097f2e174d3d4d19b504b0dd8e6a79287db1b0819838e9ce27b4b7f9b0422a0868407289810f46b94b46ee5c2e3b9b84a01ebf0191389f884a04d00fc9352d8cd761d2f4b219fbe88dc05e7b533e111db20e747de821da60edc09c7ac512833f80975676f53df50990e741b4932748fd79f9a265e11de662007bbadfd9bd91bb42a138eb38fde93212634d05337a2ea8fe19d275917fa505375faaca64d581efb617f91862f369a9d5debc1c07ee8b638511ec6444b79776940de178ed7d7be2560fd0db834144b966cbf74ab6adb03fe0fe5fda07b237ed900b9d6c3a0bc5cc5c6787abe87c54a9e5665fa2ac65f80d25f354d64829c5251bb8c5f9be6624cbd7e35486074b3398448451ea4e1dafd1743c29e2f92426dd7f2d032bb579d01f5766bf931173cd7bfcb717eaff5c6df798a6a5ce1cc17200c39bb2c6bb2a247b7b36291e7ec1e8f40fff0aeabc72e7a37b85462278f8d9ebb136a760fba3ec5e122e34fda814da26691ac432bbd707e3fd76bbcbb4472823dbf71c9d5469fbe73538df7669e8edd9c7aaf0e21223e7e9dd77b3f36a113efcd8507c335189c2842a9d0f8b02a5b8456245356f3d380839c3c2ec0997b28ba27371fb12bdbe78bc4546caf725e6dbf7d5694f9406685c9eca271f1a7fae59be5660f1723f5542c8be688be455755641aabbac3caf465d2104208101d3e11da1452e27fc4d8eb3e65753353ad3098cdfda5a6fc18c37ec2a173ebd1e57e1481658cd9e0a989f200afd8eff1c0c1a510a6dd30d8c123102ee48619798d8d84f5dfb202965b4c7e3c862793cbf338b66b2b91f2e64b8752e52a839fd5faa853725653fe45fe3c5e4dd037a2eb1ac467336194b9f2b88fb4eaec966086e3e380895462a56cc5f95504811317dd4d7456b775044d8282e465e321f84d4ed3e981858a4e38753eacc9afdeae88b74a7b788b7198a77f4aadff17c2e4f01c0e9a1f9951192705be9b82864cb2eb9251aae0390c19fa3e0589a4766e02f1ec8746fade03638a5a0c3532d9f041c0ba94071182aeff6eeaed59d65f5f5ce5a1a28f59112a9b8cf6eb4ed95c85e9068cabc80ca5337d26a2e78c422261a272a267e47b06b0c27f97c51baeae087c3ac65f722cfcf9e0a55755e11cc6d71db94e1f244aef06c43ef04af8ed6415b706244ea72b16540f01d4599b40d59e03d8dd3aece8aadada262ef5c5cd9a62c431e92ad74b7bd29e16e256a52b6e07e406cbb50ec68e400c2fd7f0feaa993a068b2c46135182e3fc145244ab039f015cee601127b33224df76363950296eabe81e9e30db72dc0dad5ff72f3e1ef9ab28005a77f05de4a44051739e0f4289e2e331e06f425bfb4045d111c940aef70102d13d9ab7db0a70e6c6a0c1893412dbeca8d49e5a8feb62f2a038ec675af9a933a25318366a46844c09550ce2e4e97802b955aecc9b1d8c67febae349972968dfe93c0233634e71f7a88fef77c0aacc39343082dd336cb7f48f9dcb059652160bd3e2d71a27bfb97fdcc8e91d0c4c445520a7767789a0533bf7381651b53481a9f584521bbd02c0614f2aa0794067b746d346c05d0600b9cf34973a8580b0c79e5404e878c908694094849ad800775da885e8129c8f2dc97d482b6b74d9f65b524c86260fac1103c672dcf8f65af834267f6e88a0f6fffeaa3f123d20478f609a83aab4dd2caa27fbbe43ad34c48a4b0c96c58f6dc9487bca28b4ae64fdb6c3c3c59a1151f8a39203e7c60cfff04cba64afeed4bf7bab61224d141abcf51b78aaa5bc1ed5663951b674afca91ec62264ef6443c00ade70e84d661793e5617b57f07520c2323764ebfea7f7587eadfac1ac2ddbcfaf4e7acab3958a4449d4e9e1ace4565588cf8f970d4369061ec8b6665818358a3b5c2b209051d10b2a7146ceaee57e3823708feeb289c0f08a41fcc2536c7ed0cfe72d3295a6363e6ee8b68943cdf63ae0a72ddf94ac3b266922e241c7bea7142064a9a9ef08e4df12ec8f172986eb849db771b5207a8638386dc5de083950b221c3420a7d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h172364bcfc63f05df81ce6aab54e28ede31c6c454617f60fcc14668d2c8e61e00b151f57a8b5c07f129dff93189c166b6b0a707c7c079d612c6d40fed1180d8dd24789f9fe6c62b6791ab0b260ac6110d1f05caa5a81df2b3b60a76e194504214c18331083d37ea0b29a1253b9054f2ebfedf0c7848e0c21dce40bf953c501dd8f4791738e6139ed031f7167ad688acc13cab89a10cf55a7379d9049e7eb8dbc7ba233dc2cf21121909b7ce2a8c867f466aa8bdb6228ed36d78f326be76d1f03038f6caed58a55173fc6c32e4658f5e159b45c21b99eff43f409051151e7f6a181ab53d2270c3741ddf35d193ebbca77fd4d6fbbccac6bdffd5ce630572d67d29d1b8112845d25e7a719fca277ff12153b86d322fb634df625f3b5bc6d8d8daa5104ad01eb126f4568b868041b91390bb2f445b3ce3c7cd06a5b29461e62df93db824df3fb4b5851db5957bfa92d24b900a7c10c66b2b29b08a594a4e42dd4dc547610bf461eb3d4e40270b400cfc6927e21137245c12757218d36b629106f6a5f6ce89a2d56ccecf7f5f00706c927ef2e8f77ec824011d6f8fd66e65ef2208bfc9ba47868657695e87481158f04c65a0891ac772aa35684f161a4dc6dda6472fe74db9e6861ef55952f78bb61c5ed68abfadef86bc0ae60a43507492c66d6be3c0bc896d0d5673e8712066bcce02ceca40df1776d2830b776f0b765ccd39d22aff3130cfdf2ab032b7d93adb0e2cddc0ba9b2faae8f46bc4ed7b418b1d1dfb6d19a42a50e603aff878fa288a84b151ee220aa7498b2e874ef6c0342c477701dfebc7a2f4bc3db98607bf648ac68cf640cb248f38077b4b1d829e13e989343f65ec4f38e3cc2be10afc284306bd0e0fe71d3a62bf2f3c52a96f9bcc0201dc31ea3eaed565f2116a9f6ca3a57a89d99c4df73fc247c4fe288e79d52554d45cb6f58ad10f6965900f17c9ba4547f1ac3d3bfcf6dfcba96d2069a624f8697ba1679cb00ba0b8da1ed2a4da3b6f3ea021de4bfc46a8014fbb85dfb8bd91c176a3f5317ef49ae516f23c1f052d3c620a84d48d5dc23063c419ad1a22f69242a09ca0ef32bc994a3e19ce9a96ee6cdd47f6ffe5719a2c4125f1374080d5db804e4bfae5a9902f0762e84443e0e15336ffd41fa2803adb60ceaf7317263c2b96bed7965774dfa9a6df720c0a2fb62e0dd695983893e74cc9d89a1837a667dd90ac37ad3974bd2ea9bd0c0fcb22971c0dcd17511b488dc2660e4bd4c9552c983ca70096739e7ee7aeb432643c115ec6c5d2b2591f23d07bb1417edeeedfe74436893aeea2174a0837b33e71ab3ef416dc8e0426c8762c60ba6df2a9f14d4315f9f47a522f3dbe149f2e8a03d1792a458302c10ddab10fa4908c8a650b7aae41d51ea76acd49aef70547b746b0b1cc97dcf6d80020e03b8ca2c6a7a7e9c742bc2c38fd801c2aff606da2bb3d9ce0062ee322a4bb07e993caddd0821a702e0fe9bf02f4b4a982159cc78b42337c484b37a0115bfc7088a8311eec5a64febc327de0786b5a3c995c210723d0397c6a1eed269904870a61c9190bdb427b7f100ed126d2619b2805d75fbdafce34203110e36c62c6b468d13beef7e983e720deed16e08fd63043ba223994dc54ecb54dda35fe1ed65b7e07cde88b71ca65ee8a9c3864e00df16a607843fa0ef14f36c5d0b11618196490ae81798fa14350206786e67205a7ef2a3593b16f5f47ddc1a09fb1152335a1e1f504574822e212e0286164578c3c796b53e456b8995da3cd83606ed023992064b965f7646e1bc04a5a80313d8cff6b1821ff8d7064f9b92074c1d7442bbc702e24cb39d273d5d16e11348926cb9a043e09ddb5b74ccb946493e056a7c8e62c405f286b4a9bc9a9782c9e430a18ce44ffa2dd86cdc1ba4223b3bb49f8e95bc61222ed7e34a453f1f5bfc9668d26c92a8f8f80feeb2ea7052adaa166f8b8bbf8247a214a7b70c0e04036173e50eeb727c19477ea74622c68dcdd64161b2cc625f162c4fb928178498705f3edd02a149ecea9e6e54d60307ea6ea699106c8998b3bcb0a9f4fa173baee067840045faa5f47f810408637fae0e8dd4e7b693712607cce509d5ec0fc92f3bc77ce7f7c100fca5389ca934a16cc1fb0d07c743c686102de246298f0c152f439c01a26629f1b0fcfdc60c258a784aa2d8845cde8dc704bb52ce491893ea99abdaae370094245a19d4d4847ea8deca368b5d0a9d0733aea98406ac6ccef3381f23d1f52d801d6fb1c351fb3e9c3d9c2274afc6dff8b46effc6590058fd31f6d89441a79819ba959ce5171a9f3a7427c9ed06a3e618cd104c19f3ba92578889bd365fba1416e3d0e304dea3f2cbf639bc64af3e9b3e8f8d64090479eaa80fc28a3206ab687638412ce3ecdeee4e237ad2eec8a1089d6bacd24db5afd7bb6fe466d6fd2bdf9c5dba947e60574cf0ca5a6a9aff2646d93dd21db7c7dfb0280244c000dbfa0b28d3dded88c424c4bb8dd52912f46163b8dd5f6ebc9435f27820c566509b870fb60d527aa9bcf6bc5ea56c4563d8db09be793beaea64a6282278395dd115ccf2372c1be8e7fdca4bc5dcea37d5a180fede8990d194dac6dadc20e2860a03b4575de25d459b6fb92e57a3b33a08bfeacc645e80d4a2eb5aeb0ef56f49b676e1e656038fa5348c405d8e98288dd146b6940b0f83f11d1a750965a6ff0de5be3ea7a5bf3410b736187fb1f6a47037d85c746e9acf887daab6f1ba313fa595d779a99a7a1ef486a5c002a300d07fab1e5009ab4dfa76472aeb4190961d67b5fb08ee70d324a6dd9da4e8c4330af58047501e68b79e4d3d450fc3cde72d371f018d2e89951b4466404b6f8a30ba3839bc24c6c0dd561cd358d6304e7502cd61c73d082d44861812a9735ea7664a8926207c3c753367dc9c5527456455d8c83315e826a745cd5bf9e6761e30ed6d3120dbeb3c138360369562e17dca1c8153573c0e37486d4dd0f6a88743a898ca41e506609ec493a1104a0bf626f0c3fd84e53a2ef1f8e6886ddddf28e478cad5738b78ed6aaa84bd3b206fa28c7105fec52e32a15bb8845ec2e2dceac54d2ff493f4e3773126402e44d358d18e831368afe9a525458f0f1ec10c4cc6ce9398f4ced65f85119929515e4868f10805231e01c7a53461767c4d006c9941b6922d714e953f38f0dfac66e2f8f28baf0dfacd3ab4474e1ac236f06d144239ab4cb499b961f8e0c2613ec170d941f34fbf8803155b27fb0775249cb2c69a88a5d63e3f2ac5d732639ecc0f7397e63ce1c8fa6031fdd4fa224b287041011a3e0e78307c2c196923c3b4d4df274ebab879e2e0d3cda7b4fb3042c815fbc13c2f5a730daaebc3df3ccda05cd6b4509dbbe1431e5cd792a5fc411d576c62c2894ca5f0c261179588dcc96261649c9d2abca3a5d80f72704b99ec45c63e12894177f7237ffb6ecaec9f9c1f6001f870a72e8a0b209d562ed16786e425c167dd2812716d79faf14865b5361b5d77f36bde35ba2eb41f5ed179e227de85a9c8ae485bc8641095de9543333884e5aae9359777ccd2521ad7a189d06d9c02eb5ecd6e23765e96bc3941078e218072680462e52723baa739da6096e42ce9f2c7e05ae0c486b6a6005221bd108c8354332f1d16ef5242a584c21a0a801a82092d9a3c9521b974a0fe87d64a952359de79285a95dabf3d4fe9bd2b86dda50439e3de9e3f5bf33d50d7e9c4b41ba65716c7310f63f07f948d9eb191ba4d292d9d2777ef01a75100c7a6f7bd17adafeed41c505535151f83c5d3301c3e502571cf7cfc7fed5a66c673a8bef387e5c4b693c2b2688e983fd13ea90430904b6eeeb8d093c3cba2cba1f799b1f2cb655ac226977ae8f4b0404c23ba45820b912bc165c020464c4db1758b35093ccfd03d6b9f624acd3f93866529082adc2f3a9cf2a06f4281d1f59fe4fd222b37dbf2dce181ffc2b7f180425964e6e3beebdf88612b098867aa4cd7823c78e9a37bd6490a20c5e83c4c3a6c0416a9a65643693832694bd7252ac86c18b80521e70948e7c5d90144ac5d57a506d3fa4454eb07ba1216df3bf2a492d6b4c779f43e9b988b6b8e1f79f580094dac21a1801d11300f34942df8e8cb2047d0f695de66ecab963379e0b81473011613d1d7e607622bf5d7eae8d52ec080a7bab3932e186a1ba7bc3c85a635630d50c259e96ebb78ea195043bc1bbaeae7ccd330f7385ddd573ebfeecb94f76b38b5cc0ecbba4d949705a19643add23dfd975e618887658d042471ab357f0e841b063f6980400009f6c01188a0d0bc1342d32578c85e99808c4c354e7335631638b77f794f93260f5cb5f71bd8508a10b8034521b7baf009fe66a7c49dae97c120c95e65fe3c8d071deb2a05f75c027df151d10ead933739d277645892188c26696862fba72b9bd5130e9381a1a98b119afb28d369b0e860ff9f69fb55455c25837a4999361c38e7b0b80638e497f49ca9dd26683a6d7e270f116dcf481be72c28b12c3b8037d5ecec4699bf82ee3d596807583461187e45d3b7e97c3eb239768fbbc5d55efe9af204d94d045427fb8533a8b304228fd8595d73b55da5a238ec490b89342b2844a0c66322b87122bf307b54147f6bec0b671ce2c5488c213e0ad74680cd048cd8af2c9447e43954e3344c3dd357130cad659c65f5e92a467cd38bb5b0e0e22c027eaeab4276189f6f5a44aec2f3907255b552e869a53276a0cd67cf86d405e5a577647a5a728423ba494bc39540d455a6c497cd97f7135912b197be9729ee27acf60834d68b0909cc8cec53b0334e58e1f6edc726c40c7d9859d78ca58267a54223a721dc4c042a2db6f3ccc487b72ed6cd7155158f65f799d61b4ae80131f6c72215630d5a0e46e386c0f94cf2734c0ab9b61b3fc060b691a7e8b8b778c79bc55bcab3c19edf05bd2ff2212dad6068bdfe81d2fa7c90147a52bcc96dea75eac650d7041e7a746d519932801940ea3dba3cb0fe534961d359285fd4ca7197a045dd75bb641e71104113420f7e291a98211cd5ea5ae2019c3b7e46f3ca85d865ac949c60cd0a43f0ab95894888a36aad54cd685f00f01da75f715520dc9530b7687e6b37f2167a4e66ff35d018b8c0550483831188f33dc2d30e734ce1a65503d8cceaf3c7f6f4fe98fa53b038c34ec3778f9e03452637829d2417beaec031aa37cef4dba1cc4fdce81822945910ef028bbf46c9b8e0140faaf7832b599ce5c69289df9ca8db99010f3cdaa99497409bdfefeeca5350b995fd540a02b00260a09e196640682ceeb5b9ac08346f408db07d6cdb5bcb0bb46008715f97e09644353e0bde3cf594d27b69591279d3ce3827c12b051501dca669b971c582a476b613f010d4816414dce60b9d2f981c70f226811ae40f927fc61692f46102963899d524a6b946752de202162326c1823dde92d52bfbdb16a3869e943cc07d5f187fc2e4daafc89a4434cdea98a1c374771c29fe5ff6af770253d86884742988318c80a9b921d38976deaaf5ca16e51f5b4b77ebd82801496660f5bb5729c3523a841b67d208e8f51a3e05bce1ffbd49a6658f6dcb4fb128f0714fb8ec06b134aa81ecc7b8aef483e41e2a547ce8f591b3fa91e2216c86b1fab0da4d4220ec56e1911619d46df35faae0d3b9fd98f4434c5525da092c3d86768e46e64e4adfcb800d4d50befbb7d6830d9e6c8e3d5403396bc15bf0d3fd3ef417ecd5d90438e8cfe9139067d4d89f3227b37860411a47aa681d40cb2237175fe3310fd334397bd63c63d6c4c78f6c6c49;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9cfeacc87ec3a436ececcae060c7e648af4799ad862f6c237ab8a6dd78dfe659759732acbd68ce44dd60a0356a7c9376dd0d0aeead52c0c07953e8ab32a294bf216a321f2301711b7742bbfed1a14e8fe587244b49881f13c73353a20c54afdb834fecbbb566c1a58f3bf4b236e4ec4abfd75161a0c959b36d8fbf6d0b655919bb7e9af4cab0dc3971c81cdc78758f54ef6b833569949cb18f932a5843d886ea42403b449295f133a15384eec6ef5ec39bc49543f1b7a6d0d2b56f081c33b976c46b87f624ecdaaf2430f1973338c8b0dff1278c300f8370984ecff2bd9bdf3e49cc6706aa77753a8f65c3101caa5d92401757de72be757484843a588a50267b8fa7d9601fc07647362bb1db79556005d3d302c0b860328995da01f8f78854f1dc1768c8eeb7f0379734ef36298d4bd7af001681fda392780f8dfdb0265bca9d00193d3d92ba2793c1ca378ad4713615f898713c71acf077ce83d2894844b18b6b675d3f188f2e274c912d4cf323b0842b0cf624f4007707705d23a493a0cdf02eca37242ec3702201f04e7faed671a9502ef175bc1053fb3ec8904bd5e699e59f33c577e9b7f887abb9d39fde63b4f05b3cd4c2fb0ca5609b3fa7212a8866a405ba9b53f1d7d8ea66059833a59910a400a2cab3b4140c90d9241e485b19fa08ba5f91aea4d88dc105e31cc5b9fbdbad79b6dc542f3254ef68bed868880ec71ada10ef2198b885df3b15ba56ef35459961ff9759149f1e3d5a8993b7938ecabc70071b429dc43704bb4d36365b4055a62d392faaedf2f4d1ed5093f23618908b2f617a5f671f3c322ad67cbc632003f42f2f95706889468406c4db22a5fd03448a4095f134558834d26d192f1c6a642b572a21498682047664da1f16d338188250af69785e24fb375b4a76d0814ec6b941a4e7b6d40f6c9048790aaa90c031de5a66631809c7981d6dad558b80bc11787d3075a712b6985cf3c5d5649c003d638fcf6ff414283f6cdf930d4dd9b331d47991aa0b1a78e98fcd696d26a5fe8cd2c03511bdbf348378105557fd1c3effa3da1b714f45c90f772e7b08d6b528834f78d67956a697b288fb8f913e8c0cafc1e63dbfadb3a3e5b10db6729de6e63e618385a40b883f304678709353cfaa134e0d06b570add8e8af045c613db98bcb6e21f6d38aecf8dea8412774349a22355614964e31f83daab3474d57e2341cff46c26f72b4c31878c19e88006677e21bad3ba406159fd326e6cd3a41dcd8f1577de7c2f86e204088237a15700ea9b0401ef2cea4e8ad99ddea78005b04a4364a67df0ca281332761b948f8435d658bee19197a4cb79fa220f82aaa953cc3fac32921b859b6a468f7628c35ccf4e14634211c88321985d7a95092a4a9635cd15b8eb37a884fe07e6c16d3b5669172f664a95980a0b84235bc95c06b2339dea9018658cc0cf4ac5fc74ae3300b54b226d6cd5c5ae079b5877421aa054b9dc02af82e2998683dee30cf4713427dc48aa30ae4aeacbff5a35b8591fc5c656d7718f645ce5852f62dc01dd1cb9b64f91163b9a54d1cc17875c0e3f6284fea0aea49ec3647668468b4b6173bc97ca645339f97fd93ad6c757afdfd207f811b35e8ff9bcb2458395e513f6d80aa8cc9e4182a2b25ed290b0155b93973f48fa1029b78002a66022487e39e4cbd0a04b9e4bf62d2664e191afc3a72d4eff641ea7436f9502df3d8a0c4372f5d544e34073b18f2c1e0e585dc68156d566331d4e2440fef74b11176578f2d4b49e2dfe2341533d8185973e3eaf228fcd7588188a9e6acd4f17e59582ac8f21e05c71810a202a08f3a4cd932f5f6e74984c024a77ddca28a69575f7c3e26896794d84451f2384ca40a8ee00d000ad9b028d52911af1b1bfc344c2929e797bceccde2d660ecf43f2d9c867c8da7cd85ccd6dd55eed28b93cb36c7ddc2e461a09b3b1abf3127cb5304a14af75af1c3907115ac09183fb8279804f512ae84b37a76314d8a62cb9de2a80cc144c64021668c9d379976ed0a1ea746db6bd592a362e0209a0c9c4050c7eea0d8a2a467361db5692e3f5521f5cd950d874cea3fdb5a53337457d1b4bab55f116552ca0530326a0ddfa0f5f69f7c485c9dc556dc0ebddceac8e99e96067ea6d92ee014d5ca773ecc4f5cd7c039fcdadee0f5c7fa416ec047a27c74bf62c85234859852920e4937ccee8fa223f3c1961c69e349ae914084752fd9d2d2d14a24eadcd2f4ac3a6af3b175019a4a680e2d6a86ff40978adfdd10f1f45a9a38ae49d0b13cb1bc17798555d05f6811a82b95f88563f70297c783fd9005d7daa0d35066fb37bdd6c4925144f3d8459a4a48108c6ec8069e8011ac2ec7e0bd31550547dcaaf34946d1888ce636a5cb088a8df26790aa80efc2bd59f32ac42b6727b1f81ee485b8e2d002ced5f80e49f851c45383777ce34e876e70accff1d2c44b45a5a2cb826abab201781d96ff7c60835c92b2eaaf02eee6311fdf85d3272093b737829205d978a4a959e33966e14fa0d8865ff9807a282863fd2b04303f5f87e97f68697c795b6f66caa2a90734b40e32171b5f69c6a67482de26ee74e26a40a4ca12b0640f2ee696f88bf911109f3ab72c09534c1c32bdd414cf3fd64fe10221516041ed535c13ad70073267f13897e3cd029fbe9364bb205293f503f52f9f123ef8750269a7c1c6d8bd3208947db13ecddcbf4a5fdf5e41245fcb35cd699a3325d9efa0b9ec5b49cc7c854da761ffd0e8cff153cb3b2d2461e8da27d31dc20af15133c8633c231b1803dc795ab01bc554d4c6566a6b7d78b8aea77931ee155e65a13f4678b092140956b9efefb38c480b12945b08960063d4f8528b8679fad1c21539516e6b3fc3592cabdd33430fe98486dbddf9142974f306b6ba2fd0a29d474f36d8322002b8b88326c0074f5035bf4a7d1b91e1db08432075e4dfc189261da368689c323e1d2a4f381b81a20f884d56e28374ce4ab7079153a8b596f3b3a64a555347c828092a5eeddb99c6b184947ac64fc809b38abd25562c8b1b9dbbd8254a6fefbe3fb3150abeb7d22a5b25d1be2dc75ba333398842c3cac1b36157219c5a6f8b9b17cfddd14f0b450ccc32293ea613bbbacdf8db0adac839eb34e709577d0b83a65f05910e3ba7d6481161b38b1e4653071e6f16b63b6f4332e07e8c1b0dc9ca76211d098bb641a53f8e355998e931d030606764d982cb3349d713285ca29a4d3c2a369d8d5787665b2eee0132df8c7c550e1a6a2874e43bf7e93ae0cbb3c1615aea78a021a60ba7539dbb30879bf8b596cfc9b8cae32b29ffa0c3927ad65d904f67cc78c2605ec03fd9fdbd73e1c4d0f42d1ab1d2c682cf5c849f8e0bc0ab68a0b8b748488d66c832bb430543f6a3ec2799305810d0656fb290129026bf044042f1a3d35790c1eafa90c66770d9ddc841cc5b5498bd4c0aab92177ee1e511907d386a5fe80264c1a775094eb0780c1855a7e0913846e82b509fbbc8c7bfd7a6915472fb3dfa088e0000648ab8ba1fa619d2e43ce42048239df20606d2bee6ae016c4f5e594383449859793b1d2ac5d7159bd519ecbc5ec1a3dc1d4282b7ada917f234233c942be36c37fc5b81ee12167dc42727bd4df9b37936260b59b1b3d59f35383c81c163e5579d585b066fc19ca42fa0cbdd68ba7f1b3f20f0214c526880976e62583ef986b6d177cd093e529addd3f080657d564124bb6e3cb1190d04a2cdbfa12606a71dff5652da8b07bb990665243b1066675071d0039f6296ec94f60d7dee85f24b4640894437f5bd78c95577e39fcecefa0895cda392165f1077908a6273cc726fa891ef384d39cd838bd402486246b419693012189c02eb3ca9cc1f63046f2caf362f8ef3ea5224243911e5759e166d595523b76246f911df1185fb186f14a0ec4bed7f00eed4ce85ea27282e77c19e893a3d7c5167646f8e946360b7cadb79c507a73b2d659d97c1ecaf817cbd15bce094b9465dce3752b668fb9465ca24d26aefa9556c151784c724e4c684c20f3d0e4ec0034598f4bfc8bfa58f2e1075e3929dc7889fc56010f078075d1e34133dbbed79bbea141b015369df44cc3219fcc2cd7cc0be53c1ac8670d449ad6b2cca85f5bd81784826fc32709a6025b31f11424c73d55e7e757fee8711d15e0d802952d9da53d8cd2d6faf8d4eeb88758ef5ca5ed116be03eb7660762bd9679cc87c0c4b3a48b7179991aaa32fdea0c0830d2c3768a714fc7731acfaccef6b279a55b661c49e7a02b13b4e897dbb0665c87612aa15e9fe97736523da5da314612947ea1cb22bf8bd6bb1e01db69f40b62b333724b64fbe4fe66b1fbbff132740af48c9a123543fcb851b44b4684568280c52187a33389e4945cc640b414cdd749c26f683ecda0f921b5d28e92df62b368c28bf5f84b1436f46cdfe0b4d58355f51151b9ad99635408ae50e3e2fbd4b37302b419b39716491d28c3e0f0246e805595370a0339aa878cf53c6b11068ff40d2e5ac5d980cff7971171ebfcc155a40eca0c50f9bc46b921dfaaf525931a76e66d05fddf0149874daa26b286ff6394101dc3820d4671822f5dcceafd62296ce96fac5d1840bace8a51924748252a93a355ff3023fa731362043f62bfdef88a7f131d24ae6f9d18f288307cdd19c652ca9435f55429abc0b16343a6548d4826614f96ed3f1c10ff161452ab92cc193a9851289fa39fbdbc4525652c74e9655842e150e2a372ecc32faff94d5748c61ae8dafdb8a5ff9ee24d9c11aa55773b0a5246945875e6148779dcc9a928fb2eefb001f65cd971186d05c24236294ca99307977b6497424170efb50b227ebb028c2b76b0e75390514bf4b5fc816d55133b30c26851c2dcb362e37116ed9d24964198da96523bb6d36aba317dbd78a81b081c865da34293dbb1675927a5daab271743a3f36c082318b095af898d3d785315a94146848fe98f0a0a17811471f1266f2c960b9f68e4b57c7cf2bd185a1cd7387c7dc5142dde61755d56e116062ab8d9ed1fa2677841e4d1cb95c9333230d086ba4fc681cf7327e3d7203c73e14075760be9022958a233de3832a63b4a465f77886a2431530bbf3c6ce12c2a6c84d76d9ee783de1084bc777f914a2156194636efd653368eae1205770d9b3beb26d67e24ee70604dffc65634df91ba4d1bee11a675c4d55e5c1ddc09332eb2522dd7bbf6b4014f1050c1fb594698e38aa46a3ee8c96fa353596d36428d6453008934cac12099e9b2022b4eed97dfe31376d19087ec1ca9befde6ea5a2e78b3d9ca6b76f976598a3633b65412b6437ff73e8b2d5077e147428a88f8b417b008b4248eb376ea2ea3513fba4b23b13a193fc155ec36d91431e094ad6acf9a630717173c4807954a3f178e84883bf577904bd27078e31a1511b43d24fe9329d0790a5e36d2d4be9a02bfbdff9abd6dba16705acee9e1ff19469bed4f1aeb00b752c0f419a6c27e78ccdc5cbb25a8f9015deab3516035032ce5744fc15ed7fcff038d4cadca8f2ae3c133d29864f129c98b36fd356b2a818d5254579df68b0803cb70dfd7575f0ce83847b66dd05c3f192b5281952a7aabc9674f1b6c3caf37606f6bf2b08f71b9edb03c0248ca9f4d2486dce460e5be75e336f9c532599d7e6546343a441ac5472b6f7bff54aaa2326589762d89256f6dc76f2edb1c7fb1ef97dca1fee7cbf33e82c47aa384c4bcd6322aa793cb71db7a7dc15c024a59fbee92f20d8bd7d30961c1ad0e34b1ff58d51168d9c479dc9a8b12b1cd73a20cb7ceb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3abc47e9c12c18ba9fc48d67bc7c3f161d43c452cdb58b501cbaaa72f701286ba531010683c70e96a7299be834d624bd3c3c14ab9a1c49f1d6c284e66165c9545fa549608463b79cfa13fcdb950397f9a9cf4374307d60cb095202a2719def285ae48719c260421090d9cd4d47b689f7d4d71f96304272f469f411e0007d589a0ad478db847f8c18d2b5b2ea313ba534aa51b5f0334c1dc8aec3150e4c92c3bc4f79b74020d7c1313bcd895c50b508d558c801e3401d53fb45bc36192025f9eb4bd12f088b5d2260806a478a2fd3a41f52e8b94c774c20f35eedb28c388a15959df0356741ef93fcb1f6b603639fe7b9cd45b2dbd370ddde83223931e489879eb08bedf42e0d9883dad83b7ce55c9c7d8549a3063b7d3fabb39aa85e268c8e52d2dc2bae89f71736b19ab82f638dfd41db0d2476c003f2b8e6a77bb42385425682c23f8b96123cfd10453c22c4966440d787ddbc9904da46daf1cff6ee09c92b985b1517c6490c7ccab27105fdd2e9f773f58ab07a709ca4e9e45b2cfa4583d7f898c9653e85e4ec23c2f3eb298c6fd841f3fe4cd8b427141d696405f52d1cd575e07ea9aa0b4bfaf7badf2a77c45ed722730bcc455b595bcb6f7d7cac2f7758eca94e9cba64379fa9f3bd4710505ac1390672b83a88160e306518727a10e30d66be63360a762862559bca4706f6b34adcb57ee9e97619044e8badff6e90c4ed21950d7d69b0c33b294ecb886b8427b673f38a979c5bf81e1881465f6fb202ff389e3402917c35db57e4b9dbcdf184118faa9a652c7cb4b5c229ca5d3bbcba174984bba69f5684991993bd15662ae7fa2a9a9d98f9e857c5a9ae39ae9904732558b2f6a7cce436e141af0498755993500fa42a3aea42e4195d6f6a94fe0356e16b9a9d7b7339e438cd01d72f54bdce94066322056d139b8d930ef0e25416bf2882ad32819c3c4eb10b6a049a5a3d095fff7375a7406c7451421d7da1bd40985a18ed13d737daadcbfaeaf266f9b409163ea0fd34b928173ddc33bd8a9f29598107a5b78cb0b0510971bdbcec2769c6bf379fa1142da485660cc4e0b93ce94b5ede2e72c0b2ba74a6adbfbb211b42a392b52f3c35a9187749720793dec75fc4f2d5362200a5e2bcd491f81889ac4bbba09a1150ccb6fdf35f85824a676e0e69da34af699df3ce482b1d541d99d98200a580d0942cb5172d46a4c775623a3c4baacc1a79f2d36bdc0aba75ba796a3ac753b4a25b83d96917b78f41ade0c23e29ece6dcd89db2e73d3751a7a112dd0834179de24f9d9627d68d4553e83b31e613f286d677674a91b2c7682beb9427ffb8af9437f41fc94702f2774b4179b2d85fbd1266973c2c523d1f77065ae5b4794caa3d0c1d9b398748ac0b375bf9a4be5d9065adbff081f317faa656e4210d06e8fda8b23c5ed6a92ac38c4c03e940ffb2153bdc0fe6928e5f33ec23dedc8490fa6008c44eefd8ac72ca2b49b371b0e92dcb38f68d4421ac714c6c8a99e330957d02509ebdff57f2452f552bde92a39196dac36ebeca5c5e71162a2ca28986d87e6326006edd377934e49dfd5b46bf41de683f1411acd144a116b97d05fd1be2e38d5362ead591df7aefd2f44547b2ec2a19caa76e035592dfb592aab0f8708ed00621b45be2f601ca3607b85617edc01d33f233a5489c6f05dffd501ca13e02139e6837c9d4eee8437a1ad189d51802eaea26dda20a4421e3d2f9f5bd29bc77c2215c880cf4907101ae2b2a5c9e202235d89da7cc2f67d00d627ff3fcebe991df1ba1a3e32729d2f0a19aebbf1d5b2d0a683d9bb0497e4200d7ba3f7cb61ea1490abd2bd72a1fd7f2a0086c547d38de5d2a9e1a8500da06ac853641ce05db8db6645c37883472e26e45ac0794b3ed7ff601dc267f38c4d26088c09a2348300bf2f91bfda11218ac10262ffe06704b931f63227bf43ab29c88ff078b1b686bc98c326e0569e127ee58e8508fd2885935151053e4f5a14d15b0a44e71f2651dfb1993adb77f90e52674877012e16cbf0e656a83ff7f031d6ad7773b92328d4de712956205bd1b0f4c03c8138aaca032ec3cc453568e3487d8254d183aeb365f00a384f38bd3dde01e4f5bcb1a71c8ba66a16a7cac1b8b6739968d1b1f27da521cb0176c2f48eab6cb28af95725924c9f37f0ca73df4c11b390ab273dc0b0d12546788edd65e5b18d3e08de06a890c7748386a501bf0b31e29ffd8de066ddec285c63e52800b45164614665b0ea04dcb560dff94365847e5560f02d53336b1296e79508872692ff2e2a076dd53f55ab789ee7ea9b3516b10fc0e0f824b3efc44cda60828f4ed1051262991ced61b87216f97999b902e1449b199d43134c8a0b224af084cd7b4f8992d3071bd79f1095894f348e6bbba3892c619c7110c6b5259a3ebd60df425db49ff50be379a5eb6a350995d19b2c8bf12841b58b13561f8fc8e0ee4fb2147d1364db3360f3c514e016a504ee71a2ae034519f8028e88a8ea99274a24ec6de88c1eab5f7842c66c2519562684b56b1122e8b4ac64788fc0fd577f827be8ffbd4e48c82139a42a17899624425fe6bcbc832881497e1e6963affde96d7fe34d62715dd599aeac06797c65fa53c9c8640601f18f8e53376e1567668d9c9af2d537cea18f432cba9ab6b7fc09c6761404e8f12814f27d16fb19c0913bab25963d222f44843272d606ab53f01d1366cb25f0ecce718b1d11e0839d51146b56d6d5c5c348f55ffb3548371029ce816fe8a209beb05ab47dc095daf7dbbf21cfcf918dac88af1fa03c4374d35b38afcdac457b1f181d3a0607ab1651047e352f507b9a7b4e6411ec1ec2eee846292829eb2a7db6e6ce6e983fa98dd0b8b725aab83f27d2510419ea4fbab509f886d7aed349290449e14e26fc55bf3732fc80fa737dfbef153b19bf188a86784f748e4b92350a6d19218f3195d76c483c421dab09c9c19f4ac765c8c2390faa741b112b404608985de4916b7168ed2d2b4396278c5af4b6b9a8279e6fe19ad43082aa5712fc8953f81a20161e0fd56eb89887a29dff1f222f4ad2feb60c6c7d7e5f1a43b0f234cd30265cc208f8f7d2eb209404930947ac231ae05da3ccce5a928c7b75b3f9c17cf591ef9d71761b90308390af05f1951cbdf2b2f46fe9a66755f32ce9890a37a8c75c702852260ca117b866930682593c885481b4a49c66867202aa5c71ae42a6e63b39e3c9ec3964be0d45c7d471c7584002dcafec4cd7a1c777b5c55951977beabab39a5a64c389516b1ec4616c03f12c9ca99e95b241938f34569784be6fe3734f3edcd6d2316ca1e0151d5179afeb946cd01069bc797f1248bbfd711bf7f830999f36312955bdc799a46fdaa9aca755a633d10a3fd9023726f6187c2a14aed74df60f03831e30c0d00f43aeda0cbebd56f338d63fb5150ac624bed7deca97024243977ec11c3eb9927d181328bbffaa102a9b1e3ea5e5c9fc2140bffcaa523e613896f1e7da3cf980ee3a4b9b07c87bd175703466f4c240d6db7159c95ce6f33597af8daede9ca34e18c90daf1fb622bdae776e164d21ec32f05dbb25a15720d18007bcc57343666f74687138be3bd4e9b7b7da8f92b8d10e4bff5600e72e27fa3bb9c629a904fba909ec6980daaa291555733db691313f8e847946975fdb770b06acb62c00b0e7a789fa788a7082e58628caa198124bb502512982cdf2bdc96737a2c9f108603f52cd70ec026e693b1d1cdb21b32a669a6eb0823ae11d2ed67eda13fdee2a4f81d0658a1d8b9bf78f10c406be52a2a73fe712c16d02060b29b58e1b9e8384c6d48e9cefaabd22ba4d55a4774a98f13355f890a578707e68a15494927c3b439dcac72e96620b94a357d838e2028b757289c6240174aec5e6c28f4e1d06b82bc1bf5ddd3521a967478c32a49137a2f44342e8884284036a6980df6115b4a80d556f53203afbb1bf75a48570f13d49720a93e2ed314ea2be5b25b7587910ff0327083be3af025b0191d7b0467f2eaa5477adfc8caf7c69221f21a556dc1768e9496afda77f360d5771c6ae9bfe7f87f9279d30c37d967da91d0d701baf38b614b8b0492881a4439fc742134be49c03e755ae98216149d38a5fa6da7e9485418afbd13b9d91de63f014d17d760b01568ed5599ca7d5fc90124641a4a7942a58f8f53148c39928fe4b3fd11ec2211c149f773e07ed85ecfde1f44ed3f5f3fdabf4ea56bc67bb5024b517d93ff8ebce6e2d86aeb3fc2e0a2eaeed655bc3ef85466f9c1bd4beb5949e7ba1b7217ea017a302bd5b968ef74996f9b5da9f6186a9beceb3a6a8ee83dfe8ee994dbb1ee355c7ed73cde37b0338b0496b8931f7ee7ec5a953b3476576b9538c86d79a052d56947bb70216cac9a1e33f51b21ac86da9ecbc988ffab6ab48b4abe99b9959a83a3a54c15f94cff446091bbe8518e2aeaf5a5f4a165e681d878866750b8bf492fe4fa8fa842b1e8e8d20d0387795ea32619013a97197d77b6b41fadb3f1080d62b661504907df9cd06fe886a1129ae1368c755a818521f320d19f46758dae8ef0833ef8858e79df20d534a41fede6cc3789104cdfb7839c61540d39a39ac8869e772f0e334f4b476f2fa5c0c3962f9f9321207001c17b56009fa4159ad888f73b1069bfb37ee9ab6de414ff22dfa5c857f1703879b0b3fda80cb9e473660f25e34eaf0b498649839a0a7c00bfdb8ea5a3afc3f1a31de8dfd92dd293a0abf6a4096d9879d8e14fce1c454651a21580444c2d37238c9be37902612eccc5269cf2de175418ca9559163859fce40e7bb71b0cba50476ffbf5ddf78e61cec73eca68da8afe212f3706a84886c832b01b8561783e56f2a4189b7451333a1a116ca8585959abd7bfad1195e7b61c14d29ad4148911632e58b09ca1a78c1bc78e095676d28fae532b53bc1de9aa4600128d62a1a25ded35409062be0ab87fb98de3240e36200233824d4640e9c7334ca3863963311b661475ecdd371e0068304a38e345d7acbbd260872c24aa3cd409826b583ac49fc483e9d54d77a7797aeac33c607e7e12f08fa0c7cb86faf6fbe177f65725a0df89a4ffa4b6f5ac9cf3aea50a83c777f89549482dfdba17d44441b701f0a2969870908bd639cc88230d82ff890f0e535639955eb80ee0156cde9e72d9559f32abff7856f4331110094eb2b12ab0179e993994fb316412a10e9425d03d04992b6bbd027562106e81e0026933cca1e05ce0f1434a124f73972f6119b60051169309941f9d0736307691977c9ca7e1437c2c3765bd1246f8745e33a39d6dc842124535c3efda375339e1fa4d9f5d9d00eb8974181ab53e2b9065e7fbb8ee64c97c43be013b295fe33738fbd47f9620779e06c843058c1e6dc0850c2409061c49b6a861162016aa5665e4b6ad5edfea7f9bf3e7c5320ef91d37332f34bbf9cfc43a34db0e0e48c98199fdc0bda6936bb6cabee151ec164f051edf314f3eb500bfc40711042a60b75b13623fdad05488e4f2b99b249700bfa3c4a80e1df6b1d39aa2a5e8fed827c2cbac5a004182b70d2eb1c6793837b8ffba4acc7f9f5d21103a3ad6bb1cbfb900255b1cc015f1738e28f199a7270b01372095fc9fdb2353fd725a4e75eaeda1a86c12286ad42b7bf7399b545b7b89239c747cad8ddf5a6ea4ac8506c173d2f27e3f8a148fc1ce439092f99597e675d52407961a028b32142073a185d917396ff7618fbe1d29046b37d6561729afe817396577a7bc7bbf9095ab1d8537653cfa289ca40c122ddfa4848acdad9b8153ff83e8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3ee8e92a854185a79cf37cfcda30ebe93ddbeece46aabdfddfd6b0c14e9008c6cb976221e45e94faf9feddd7847085eb29e5139d0d3a35db2438d9fbfb18cab5bd8b9b09ec5dda3fa884367da8a89603bb073ba6263d13d7244477fcb00e5860cb6c6ee37b9131d77ee70e3a964188cb4fa6fc8916d5dd883fc3136eb50ffc844308d30a0e5ad25646a71c24e1b52380c93326fd4ade6c3853b93692c92f3d8586783a04d58a2bf731b5afec71f94395359a7809287b1222a242f2f7b5f00b4d6c48f0aeaba65844ccbaad626f5f5f74c349660723756b00ce81cb9565c4edca2ef70c48270dfb492d0b6a477ef69a0ef34c6a19a22c5519ff9846e1cb7b7d0560d0cee95b44757cf005e4cf71355b7c9a3e10654114bdb1c6036e9222698276ae8330dd075e444315b266744e330efd88ceac327a9abcf2d9d7c93881fd44641e97609c4df7f6914d26cc960b01d3658f9d9649b2189d707782d9743b4e3bddcd7df816f6c2dda37fb8861b689356235c2395e47cb3c50acc21a35a4db253832877a35a09960a04af6464ecf899069597cef3855013307c3c70319184c2d3c69091a3c65d5173a0f6e89e532bd00071cc10c18817d912968e69900024e7a6edfa4eed8c708a58968d9bbaa7b8e96f6e9a316852827fa24f0926b2b1d9386d7b6846a971c6bada2224feda32d272c951f82834895bc722bbf895ea012a2f9a40018d5fa8d9b73b2ba41a46286be731854a4523453278296c164301a049b3ae4da072294c1fc0bf7c0610e2d5bd6d7e2799d145120bbd00fda9693d05c7a2de15c2fb7474c77c3a1cc4fdb2cbc104514c8647beddf4c522430d8387b01fa14cf0d390061081666c2bd947c0f5c4e930e302436a93c8956b74b5eab6d372db95ffd8a48fd5c877fbb12406b3f802a2a6fd0b5daadf88ae468cbf31779cb185a2d322b1b9bb662aa0dab35ac5fe0bcf1f62d475a904ac60d8b83eab99cdcf62d30afdeef7442d639e4ce83f225dbf9ae08edf8499b1330a5c541e40de7693e4257ea0a85d16d6f837e8601fe51d45a168076612a750dd44df282ae0ca94a224af3ae3d135fe4af0fd078e08e4411f377101abadabd15adfd37271617b13196c29f9689d0b305eccf43fd8fe920fefa61d7fbe972d4550abf6c28b2212b43630d508a10be239e946cc7f0ad1ad1d8d1f9d9196563810bfa5a30c960fe81f962df7d81daccf74d0300e5a8f48baf08e68cfa2fddb9531c6403a654817f2b5fda5ea7e198d8a86df24c39c2a247797313f37dafa5af657599519d9126127d58cbbb5988f8b7df25f983d4381e436c45680a3e25a82cb768aa7219bcee0091e99e52fad832289f606d85ab3217cd4bfc4ef29b314d62bbae6c4de30493b830d8ced9b7e6fca05cc8627b9564b1093a0e5ad9fd5df11bfd01481fd2013ee95a44170279627004685009083871d3907a1b4a0c303bb76e4df30611fe6e95ebe5da076fbaf1ab2fd696d4d5395e795f50dac4f6f793dc531e560da856e85945cc182bcecaba5d832465ecb6c92ca332f6e75adfc3702442cbda94033dca31f51f2024fa9fd2bcf5a371c9c021cbd43937fb7ace1ce08e9e6f62ddf59a01db5997232e39bb7ae0c28b57a43d0708cb39383429a343c17e19fc4172f35131417a727fb480b4cc9fdd0515f83a915e5008988d031e43255c045e618357cef0578729928b05667dcc21433edcc447b2b9fe6847b55e0c2b95b0f2f17b1042e53d1418dc910e6c3cfd38b1ece2ea6acc7069ed932f6644f3e065902e30fbed46086b0eb97c10d068e587d4bffb763021094034e55c864afd7784b8d0883273571ea71f2b206fb48a9f4ec2e8c6c52f7fa541e02602bdd52516421cf48a2c67422cd9724e469d2bc685879f0ee9b48c1afcd54414e6a5784c63ae63738f36aefb67a8e1a3879c69450def539c1b8d4b1e5d58d99d9fd3c453176bea4c7715b15b546c088534539813d6b723a337b95e9d8d4b929fcfef6e872a22fb34501b2d3efdd6aff83b4401d4af9e893ad6a1e5cadf59a233848f0694424efbf52e4ff8a8ec3b886a5a024e87d0b500d43ed15af18668f0468d92bccf0e73ffefbb195cb82677d7d9e5eeaac0470caa93ef5bfb21d54f68e31d40154141c0e9db4655aef904405152cf8638eb71cb0e771fbe5acf2a90c63e4a2501f6bcf8dfe4f6dcf19c534f05f127454ee141866aa2c8eb21cef2de262ba43241b3bfcb59d5a3193706e850dfbdcb8b5d887de8de475e52e7d24ab494f7f4a130b957dd040a4e870fbf38b0c56f715c0a8abd5823cf5f5d53850a4b2914697367b78d3bf3ee104b5548b7c9098e01927c72981deb29fdc17c2441c7bb2f1eace16b312c6ccc73b55d01cc82d1e82d816d35e16c0f1de77d0405fcb395ccaefe9fb13d03bf3e08c9e12b20cdc552580892caac749b023b9b3cf3e176ce33d9c5a2223a2a3faa9ed47f952c616f859b7335118c22b76ce3286cec934ee29b28783784e08278f5bddb7108e4cb2740fc0053c4b2faab77ae5317e04f4d69c8cefb906d2ba641da69bc99af44a9bf28fbf2c8a386de921964535447c4ee234ee293159e7bc72d25fa3d05a4a494b03a22c17fcc4f9e3431578cce88f7b6414f8c7a8c44ecf082a11039a8fca087bdd2f5523287a118869daa43b33b56192dc6ef95126516cfc4e64d6df5a95d87690f8afa249aed1dd5dd3ddd406d0196864f9c14966b0372ca9386f64285bfecb198557025bccebf540c437023cb1dd037bbcb39bcb224fe396c49e487703df7cda18afc52201026ac66505bb5a9b4c9c376956ee368a95599d2a3f4afaa9feab8f48623f11add1c2221c009f51d94971a3391d467e914d3254a5921bcb18631a35a4988f43017e8a6d96825c458eb4a51104b011b159a1743d16dcc28cfcbac0c8ee0eb92306a5422de6cc5efe5e3917f8b3ae81a9c0501c5f294b297d1ed763ba6128a5a375dc5cfa4acb0a9e14d48caa84429fd339229d59aa84a16b550556ceac3ec15c341e6c0157372e80b46b04d04a0006565aee98321d3e1ca4cc3f2d037a277d069b52b1f0eec57efc891f82739a8f0656240934a9ef64d75f811dffdd2305875d4df10769112650c79e40cc7239293bc21d3f1dbd958f57fe6af5e73633fa86a17eff3542f629df2c838419d87d8dd633fdd378259b68086b136507c6ecb5dd33c6bfa7fbc6a903147f4d32a9a3e0cb5be323cb6160d55fc45686829d36a45e6e1c405b8b91229d7cf2e6e566abbc357bf0c70eddbec6aba6f48b69f5c652ab56cd6187330accb7b9b2c3c1700ee6fec4b1d00336ea5c235d4ae25fa711f5eb0ae822a1cb3e14b2437ceeb4743e9250651c33e55792063b0c6aee66d1c83b56cc9f15dc87e1d2e938ab4f2d5e7ac3687ca7aa3be5708e75300ed88fcae537dd7dac99636b5fa483068a723efc934822f0fbbca14a76154d6159b5cf12d55b4bf52560a573fc9a0192aec41feffdf3b844332e546ca9c6371ceec7ad9ec66b0a11f240d6fcb6c4fd49872c9609d1bad0726a465e8d226942399fd504d95e49581f82f118588edd7802c302be71f2b74fde01ab143ca366ac2a379d2c53d1986db35f76c880223da6354d4c238768e3627c17b86f226ef1e5598bdb4b79a9163e5a8040ae4d7588ae7710dd1f2ccc444bd7d45400f60998e68ec661bb49caa60a6f99edb0ecbe1ae06005115d8a14ea6bae25d349613e6103ff5e80d0ff8d8d0f90959987f69966026aae34a4923714f781b25a228e1146e64d69643effd07da2ccc5508dd72306a4d3cfe6dad591b7e09a6bc8e541bcb6bca3f01e3d2f57403163ca393f11f66debad316df010a47888874e644ed19301288fb312c13f17c0416da21ca9b6e337fae101e3595ec6ec47d25f7f31f91254c7c91305331b32f759bab0cd67a543a7ba0ef84732effd14b2438773f0f3a3408ac85a997e56dc6c4cd567dd815c6cb73e17f15e8e7dea413250f6da370fe68aa9c46d345e725f5e08334dfdee5f4b28cf8fbfd3afef90fb6a0ae5fa281acd12f0ac5e48189a03c648d6005dbde1ee19acd5e82c2bfc404e28ecbfc623b480ac5f680bed473908cd5e54aecf8864e470e776067d393ae65b42d10fd30b6ae129c031af47e91dbcdd80b4b54ae1dad7e7dd5c5cf0618fe4220632cf2c2e77ce4d5b4f70739aae5d093ff61fef2702b4c8fd2878282ea3722c002d4456a9c076ed778e739713584baf2652a765eff16518daae145481fd08b28064ed7ebc73ec306be103f182906d282d8e3a92b8d028fa787b4ea4aeaf1c335bd32df4484620d6a723f10b72106670c37dea362a85fdcd5ec6b3c95fb2485726e8dd0abe5ed1e165543d493955d48b781a60fc7f6e514744748ea63b13f50368b416877cc2c23b6ceaf695cea5e524b0ccd153cb84143c72f8403d7e134ebd18597c01f90541265a844e3d452b4dd9fccfbe097af5350567fae7ad06efa1f71db0c64dde67712bb58c7d216d264a0f794f9fc26c673f3c9f6845fc55d480595cfe6111337b493f319bc52bc4b5126c43de7f8c6248706f14973650d0d74da7c0c25920441e36c57483e347e05c3801924d52e54fcc392c73e25e0d2d500441b4ae18021262bb3fbd6222f561b609674576a904fbc53224898b83b6afffdb639b8072a215691e1cab2e48dae4e1ab924d8b8f80a198a95066118919407800c92b53c83d52c8ca04193dd0e49b573620000451fad3c8387d5d869955e5f8482a230f8fc42ef0a284265c1207d07fd8ccc383fcacf7f4a1ce5324f93ff5248cdf0c7f049352a9f474c2accaad979a7092f623bec317936851338b9d25abef550a92136923735725b69cdf0e81e60ec5d7667157d56f5f8c700c42abebb947dd1049218431c8c714f7658fdf8c79e0726017d474b8363b1aa160adf764ec7a588d2fdc507860ccd8587f4a6ffe64afc960917faf3acdd38a902f9d48a75f21db6fec42abe66263a09e9e42ff3d7c32eaf3e5eb975042419f989704aa75fa81f48abc0b9a6c7034ffa9bb15c3843d21580c78372ee013097bceb6ddd9da5faf509cb76d5baa4ecc51f8d524bd008aec99286e318a595f7c5cf78a3de8c392205bd9d93666d3c97e72e24adee48b4a5760f6146bc9d6390ceb4d26e8c0aa9d40a075e2b793389a76856d4085117de49cf9eec822c7e9ae862af22d616369c13904cc435f8d3cbe1099989a312c2a13b16d05e0c16335597e0b39870e0889e1932062d7de2a6e0b922b4f85290f4f30c8a4382a655c69e9550720783dafe83c061b3a6457868fd3579861fe167448ad04b82199ca3b4c8c5b710da2184b0d8d4df4b2f620908446a0781d0d180981b2a41fa2d84d26d8c58ae5f8976a8ce9628fd7c50363f54fe1117bdb3687d95588ea6989fd8f95e67f94972f675ff5ca32f1631b3b9b619c9dfbfbe9260fe8aa62d9c0477f58f520612578ed61802056530a8c6cb8748e141d217ce7bcf0f11abd4be2796e65242066ada3fab5e82b4853c1cfba5a4f60d8cfc640f2b92bcb5c7ba4ad8d1651afc33ceaea84989a5fc272aa1262661a23fc191f8e9a9e463dc06afd77cbd5fd5207519fc4c58c90677a12fe175c4a5c1d6f25038e2392d8ac210c642adf8945173822dd85b9d8fe3885d59b268a1f64a2a50f4dae6b2bcd97201ce9db1c61d05a9f4adbcfc45aabe50311511e577e486b01f101227b55d233886d3990441e2a75ca25514e343916d1face255cb37f7f177129ef7a62524e015c5abe45f16971;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h98e084aaa54d4ef5ab235a09fa01ab84278aef04ec3afac27adccf1a893a215f441cc8f8d90756dde8925f41edec3385719fdef103cdebe72edf5943b11b3c498d4242c8a2154a66ccd9cf35d6e55f809f5b8ef6bdeba89b88645f52c99e2b888888cd6ac7f8c7b05db8c32a451a48e7395b4054f406d1753d03f95f8aaa31e300c7adea1a1388787df60dd4b065fe3ad568ed61ed759fa1562806170cde7cba2dd040fa72c463c6b43334a7ac1fdbd98820f88fabb2206c3e569961796f9c178a26dcdd68ebe2abe256878696372c764510742d454949f2a1c62d50d6064d1348a7ff5c04c6614e21b732b9c1ee8ae1ae719c2098ae0f318dae81fa148e045e16605e2f60ac0f8030fd5b74fc56efce54dd0bd91f96f24e2f94120da0c7f0d05c815fa69b1faff177c21ad83ab10e90b4c3a19c174e23830bf718f75d2420070f76954d7a484d7cf943ef6a7a50929836589a1c4db9d6a62cf22503160617cf7de1226adfcdd22d776466af9823379d1c61a3bb0574461ccaab807d5b4046abb1664e757b5a5c3a0a4c82b28c07bd849df80024224f790e931fcba804e0bfd1e42c8625d9b2fa05afe6738154bc194f5b5aa1dcda11e607b15dc2f0585ff4981a5295f1787296f6ba165397b3a813cf9788cacf905665258189e9d45457fd988e6fb5f83b9d0443d87928ab7e35d386b34c0d5ffcb953d6cbb37d60f3a48e6a0f6910700789b078e235d8af1a1a9a0ea02d6677a2034120469753868af19f985f2bb5d60beef262dedeff3ed3ef0da843eb1c1c9a6d80624af7ea11aa2c2806161399fa0a90ab6c516605045c9ec7176bc9f8d3dd268cfaf98a363873c4773fd9579270b62c578689f8b07272e107d64cd5db2ab46455087b01d52b1a2d5e0ea01f1b18335c271f0a3df6ffdc61baf1ac2c4363fd350575f87a693986ffb9717762fe7953b94dcadd13a83056901e210d253b01bec846d0ef9c7030e3731f891e8cee75a9e2573662d26bf5653ce3b434a595e616afd04f9572a0a1b5e0f2311c93a9bf7a17a87c2ad044b9561badd54c677f54453e0e20d529adad4dab3df1d97c5e3ff5ed95cd67376f11771df4eee87a6f7eaa378f09344967face653c7b2ef46b35dc4d2de681bada27e7e0fd34d5c89ed9dd10b3d665f6a2eaf13d14e09e65fd8322958096c57d3fd0479d28b032dec65d565909aec2adbf53e113235b32eee923192f0093aa17b0b7488db24c89162c9bf0b1599194925a581d418b850e26893b546dfbf6aaf7eb7c204af0649232cd9e5f4a8a1324b9b1b2d042af0243db98d294b412746ee000970839271f8dbb88d86feec2d9df3f21432fb170341f41372121dd73cb2df7766040a20a5aac67a43670c1d6e5da8132ab9334a1d042665d2cdad368a766148c008c9f096bd9faa0271f8e026833683eb165e189f66e01fdbc1a786754fd90a9451b839587dd90b0e207e8577a0d4d9cf91319f8f9d855f24e739bdbf0074f649f3d47da19e79a4a0a3e09e026afa14a4f43a3c6a91597054931b985196862fd3f854838f91938d942d49bf5aa7a70b5fead4a0192d21009528e27f86f02d75416ba6ab0efbfc47af5ee407074603fb077a31e0721f06be9127f2c227e15c763680688118e292e629f3975494070e96fe93b86736dcad3feb1751ae7d4258b772f872f09440d334de86ed0b5a4f1786b6fd65d0333eccb788fc53f770ffa4ff67879de20840140cad45e6e1a4ffcac1f1ab674cf9dddf7a5dfc5bfbf5d53a7b68f89ce3d02e5be6cc86e4a1d7d3f3fe4b494bc0b7e6c3f8cface24d67d11e2d84ac5ae50f6042894b9ac7c032d435e4e9457c9316dc0272144cd147ae4918f98a66a7935947de715530f3f7cf9738d4987d68b23edca1768fdd764e19828dd79f2cb90ea78f8aa9627b2a391d92ac8dce84a92017b364946f99d7b221df84d92118893d80e87b2bf6022718a06eca0d28ac5729fa68559cccf1d157d6d1086e91a9025ca08430dd35a5fa82ebea6e50d24c4b37d71d809d46e963bfcc5b34dec9adf6b133a2e703bb1ff4dbad178c74ed5fb565199cd5dce16254cee1a28d47adec2dd9250ac4b5ecea915a589ca917d9d3df85cc1858d0bbd72f7d5f5025dd4e4f8995a7497e025d6de15e432267a16d329b31ed95bb89664611b2c48241da9067095ff6d1c5153c7e1c4c5d7f8a0f0b1e0ecf3293c780ba60cc7b2985d4ff337b4a9213965d9fe2eda3454fa9232d2b733373fc5e6dbd395f18ef932e23b2312a0ed0e94b49bdafa2800bb7933675ba847ef42c259449f01fcdb42f8fb38790b5a06c42dabaabc87e9218987ba827d380c7f8c127b284d0e1b4685cedf4309dc82ac3e52397e02413ac381f8c9b892791348c12d098cf168a4faa5bd54b13e027790209a7fff500fa934843bd5f1193873943dfbdae1fbae54f85a8bff8748371ed9448f95adea9654dbd8baf080b4b0a98bb3c2c733c996bbe5ac3a8158b2783016336863c0e58d290bc9ec8074e89addeed31079bd93dfce9455a83acb262db90f4055c2f5d2f71067e128d03b258e58283caf46481cf80160198028f9a3f82e7640e966170e7c08e28e64b5919210cbf304241a90640b5ca79266cc1f356be90c15d83d7be5bd9f006ab47a35f6cc60a51f1768162ac3687889012bafc5e3d754e0afef7d08c6859a537f28733ff6898a643aed1c169ff3c88b4ada0b35a21d020761cd24f1eb1ac89f787d657be9c5e8e3d1e0ca221b5648eafa516760a2e5d91aabc14223358c0a135df2ceba684afecea5c6d11ed2f9ed5884fe203951a5e365c8453e93fe46ad908a82eb5ac2f24f00f637587bb2d6ebcf582f652082c21daf62c956b9e93d116727584d3dac9c11d7bb38b919067d2e7898537869045814389b2c132f89d19e78ad49ec43b652bf42be833cbf856c222370d97c7d3b8d7efd665217cf052527783d25d074136ae78df8ea9104848fb036a1c8636640b65ab2dae91c3a66d60e15950d191d6a021c4a04e226ab720500ba01cca352a50f6390706f18c689b8deaea606e6d38c2716a1bc943769a22101ba9ab012f2caead1fc4ba44401a1347f17e4eed3410c78fe3832f544eaad1d5260816da2c751ec8bba2ec91e8b1abd913a275d78272eb06654ab5cdb09f2c83d512c844fadff14baf8dd703b94593778308e2639d0e821c45b1ae29ae2823a549e6676026c29295fa116fdd36177d591253e31407c34a7ed479e78c91294a62f5c7fa693c9dc4b0ce9967932a337f82dc4fabfffdd540a3f7d1bc2541aea3e2c6899710fb685e1c0ad9f6dd3a535225aa8260a12d12c84561446a80087ea9606b1517974fe505e145db17d3016afe1756bdd4c69601b746fd6afd48f3eaca1155aa03696847564e0a37bca1b640437234646918715516d21953ad658f6e369407a4b3d3e7a087faa8c0f6a053b0644e7a133445af17e38cf6113a74a9a95df44994126d7ae19fcfa16dab7923d7ea978701a96e08b1a2d445e18254cc7a9c5e7ebf8d3bf94cc3b0366ba18391ecd3c1251ffdaea3c4762710bc122d0d7725fa8cff6d9071b370d233bd4a3c9feb910381e1f9a498d24ec0945c5f8cd2d2a01a1dcd7bb49a324fb91bc8dfeec988188a55f8a72f80d7927dce0ecddb6644331b3e473839a3d724f8a4568170259d1d58428d8e47d5b4ee6179f6f2908623738134c4576888fb08d610843c1a2d226db1af7c3a0553f847929e1c6239169c1cd9f54f879b1c51fd9b78ef2b74690082d483754e6e0186e1b77b22340b9250775879acdf763616b748bc8e20c94bbc96105e64e6456f0777a1d9b158f49d1b6289ed8471bf0c1b90226092e4b5a9be1f1412299a1a686a1a6e9c61e46fe144120527ab896436b807cc4bb7478e4c7651233b878c4b1d4f5fb4714d0c15f2d739c594de74ebd57a6ff51434558e2b463827db199fb73e017a0f39bfac9a8092c9441764de701d8bad78537673d61a81e9577ec471a6f4ecb26fcae792f0b92b100b4e21f95073a1c535e90a103871189d56f5b8ff97a8cdfe3a76d98af6f5ee42324a8fc74e15eb49ff261f726477ba3546d92060fc22fa8090c6118a69a05b2cbc8366e5385c5faf053bf1f0b936c9310e7f0e6d0bc3f292508e7b00a52205ad75e358357885f0fe7b4519b06b0ce1a1d21ef237b19ff4aed502a474db070ae0b8b913d00926276ef9c341819e686a8dbcf9e29380c09f2af33fb1bf60d39966179d833800fc1292facae2832beb024b115729501d0132f487e84750d9a511d670bea4673159fb8bff321bbda7c39ef40052dd89475c0c211830341f0e3941047633dfa5797a276de4dce2e4a2cbac3981ed530548b5358ace83bc73a2a59cc2b54b2224be0b9be31971fb04647fba78236dd54a0a63ab35a6006252c170d2031e0cdd4c8c2c4511a0859e45bfeebffa7016e5dea1a6953eb463427daf932c7564e0f86d688174cda646019f9509a445bc4eaee14cf56b2b3fc289ffc06db36b7e9918a6a9dcb320bc7671deac233d887a1620fe15ae25dffdc74184c1ac22ef13266db772ae24faae6cfabd501e484ef82f4911612372ba708dd7158b894ece1995bcffde3f496cffb09c0d7ac93f54bcd35a45bd097ede19e718bbfe004f28c96305b03e83a78cc9e745e6a056a1bfd6bf51ecbec7588521ce6d2256a4c47cc9f36a0f8c91ebc2aa4e63d2304c19795bde78ba7178a263361c8324c2fc54156d35d1efc9e06f78f11c7ae7252261ce47b996ecc7f318b2d67621122f6327217a3df1b846663673da7bb86a9db20a1c2645102a2f1fe07f4fc888c049183779f93fa0205c1d4ba397c3d907a41608a34440a849f786cb6d667025e4493e81bb0a5c669892a163fff15be66c9ba365b5ee72991be1149bdb7ab5774c026e01d21823c4b9069dac4d031158f82d6a3928a20193d2c7ce5d18d08156ba032654e69cd0db6d29ceb9b488f72ebca3be1cff2683f1e6cedcab31ed829289d357c2ac8fb688a2f90bf4391bf8902125424020277353ea05b11a782b02115215cdd5a51e8da7605e495dfbba46228be58c9d4809160372067733ce4b9cec9b6bcd79a05a8b8ea98c2e4b7e30148b6f05d2e1d140ed2c7fcc0a3c9023a063097c54c920ee7660cb0efadea6096242e80f620801defd83e157be39d3056106d6a284aaec337f4ac98410652dd69e51199933604778ce11b52a74a42a210837591252a98ff2f9731ef9742c9613b9bc185acd5a7e9fe1f0df0633283a2c143360a253e60fee76ac532a2b5b2727b3da3d75d8244ac1bda577cf3e58392d28c21f8328716cc5494150d2a94002e74b5f2cffc65f1658d9bddaa021a5eadc9caf050390d77991ff7cad0ef13dcea6e472a404d42652c86a42ebebc5afa33062b45fc5ff628b4cea198b1abb60c2158ff8949316ef58707e601d25282f9b143c6047ff78a6e497651fed7a96bf77713951693390037a7be20d12163744fcbf2d7e5042e3fbe2b5cef4320ae9bfe6c2a8903e4c1d7f4135c88c9c434842861c39765d41d9200858299923bcba86253e1079647b6a83d7470c667e02684195780e919f324280f5bacbbbc4a6b53d70871164d38b3c5aa2560aa6147134e1a7557256f88d3d7a0f2757ae6453ad98ad2db700ece7fb3898b128ee967cf4b04131daa0a80a4023b10cdccb76c295e5952de10518798dd2489c30871481c71fa07db605d30ae9edf735b4096e5334d2ec49bc48572ae2f23ef80d81538cf8365f98a80c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf28ab984143030eb3fcc98a686cecedbbde21015c9db814f1dd9b873e4610840e2b64c9c58b3a241b55381ff2073ffe10bed1e00ad0220093caa068546fe2480789ba24f77263efe8140a85ab6c5a6637cff3949067c24afbc0e081357367517c08550b869e04c875f1b488510bfb753029e90e25026adadeaef99de98c65238f06128addd743afc3d69bce8629714c948077d5d389749a01c8e84ad42c3b3afd21d73e92a5f0330b64c7b0e24b0c19e0d7339f20f8a12c1848e8b73ae27ef2497db681caf918e26b39bd6578af2da04bb04e491aaa087a184bf553c73661c07213a937da42f9ec5782e833968873484c3848307f246bdedddf78c6fbf19acd1dc8687fd233e8b22baa8c97c6b021d2b29afa162c89023ace5beccbb2d6ba3625bf612d2bc562fdf4aa0deda5d48ca773f6fb694b274fadb4f71b3d0d3e2cbf18597215d8d00bfe7d9631a624f75c48883d159065b2b4642d4c2062b06142892df3f79b5439b2c3f09329a0e9e36f9d89d01288d78fe630329381edd6aa96a87300e905e2fa25144f70fe182bd45daf9651256e20c4560841c79de59b1e4040fb1ac24425a83139433784823fc62cc327f5348cf82375d592594f17503fe55ee20f11e0b367b9023724709b5e626fe12c8b035e0a8a14a6f232c41b8b26fa6b89e07c130ac39dd12d2638cb4af188eaf4d064f3d26aa8d64471becf531ab88ca2180d45e9d27e1a41d9c0d4c63df188bb3021f808e7de77090452369faff7df535640a100b00d06e8a01a39033f3cd988bc83ed4732780ea344cac652dbe11f480fe41a1b2811d01fbb5e86c027c5ad9499951f9da2e6aede0a0981228468550337c20a506fd67819cc3b42a14ec0924828bdb7fadb5cb109ff0721db0adf483a3f037e755004dbc2fcd09a02ced05992db27e15996e484254abe573ea7610c9e92551388a6ea34ebcbda0c3ce1db2b48ee74527c82703fd7576260c22d76957d02d9dbfe9f8f29fc1eae408f02f4eebc581f89f33306093e18c206c3e496e02dbe7878803a6fe3f12eda9cf923eee7c3ac908033886c6053669c10a0a26d690bbb7e1b2b9ae6c593acf0ae28faba2dfb225294af3f7a72291c15a1451972f745de6008c674cd89051f2a404c359503101312b010b4b9cf5a53ffaca04ad0880dc821fe1ad163b39d3ae30b16cea3df31020cbc188defa30fea3fc1ee4d9e4fe22645c7d7367b0fa5add18c0cb5133fb37d3940bfe5d85e0114e6140b28d0327c7a44dc8595e09872118dfb9091becb293ba88e688620432ee372a865b04438d0ed39201298096b50f74bc91c121ccadc685ba1c5e677053491a1d1b5a03f3a177b36527280d31dc6cbcad7fe21ebd5b4d8ab0dbeee9cb1ec037c2f23d544f2598dc90eb1eaa8d0e55cc7d65c5edee36c1fc9ceedc28da4126fb308c7341c4026aa22eefae6ad695f421bb2fb90b48dad154b165b7d614ce9306fdc60e4253fb2bb4894160f3c23f31ec5de75e8105e679b17f5e63fae6fe65dfae7fb442922af1cabc5d19df67d50e355f0e73b27f48a493253ed76ffbb0cd0c033d163965a80ed968e062720825d8c18e2834e5c95f2f2d612b03fa8840faa78ad8130f5884309cdc7b3c3ab3189ba94961283d74d424c249cd3be7cae3a5e00e25369668b1e9ade1d186d560c31317957a986d896871a0c9671d6200c5267bee8f189d693baf213aa6bf7a15413ed17d54cad1d1925bcb66063b840ce38ca5496cecbb25a67ee60f61a7a0136df08290a2a5f21bdd7038389db3700c3986a2cd83febadc6ed9e1f6023379a474b6c054e338bdae0c0264af0f8e438569b61e02aac043c098ae0cb68238bf87dbee76cab26ff342032135d32698ebe1b028f534603d39d9a6f66fa5ac398cfb1ee660dd14973a6a01b2096fb599ebaac960c9461319c5af007b0448523d9169c5f44f55375b89bc4744586282820d64fe3a8c73e3883fb45a08eba59229a5116ea9aed40bb2f921535df9bb816e09a79c8f3f34f80c5ffa9d094c214ef704c087fe16af19dcfd5d048e9ade2fb471e8490452e960ff63f0ee0e0fd3596c9fb419ce2b509a505dea07d330c03ca824d78e7570fc5d3ce00ca60524a6e4778ce3c6e827176d60ecf6625fc0097e4fd90c57b10986ed2e0082c56ec89371d85680e628ef97e90c670a2aba4a0b4a895b496418c8d75e139750f2251da42a9095cea04f235125a9ab47a51dec9053c2424a1aa907bcea4802d13c58b20c6c68ec3de3dc94ac0504499792b65bf054a0a8484b6ed48c275f15ccb419d770df5431d693e68823a75fc07382d6450bb1e4a2c8f68f7669703b5c6db05f94ac17421cf0f65857af56a1880ddc84f8a8f0dd0b59e7dc268a288df01c5434ad3aa4fcb04c08ea863b5f4ae8e633ee4347d27a7b0e1bf2eab01236c430278ddf7667e168a20fdffe0db293b47980c82d7f938c0897564184043478dbd77d37811b1aa971e7f79dd4494e65966ab0ce1a7b7721c1c31c2ffe0820b7b53b0b50e5db2518aec4f7d66beff9e730d60be93c0d567e2e8e0cb28cfb204c85374f51abcf12eb23828b239c33a3a71d6489d7b6ec6bbdf7209e9f4335e4b767ef785c70bc7358900e93027343bd2f690a73ece75e239745e69620cc98b2031ac8a84952e14862aa575a345c9efff772981a7fb466ba5cd6cf09d0c998f35ef02dcc1e837bf054abf040f45b7dd030caa610499c998de40874159c752c1ea886a7717e4a5dab7456e07f396cf26a3ca493f9e3c72bc5dc7c9f19de8a22e53c217e1214a322b98487103a9598b375597445e016d67c07580ac06621be299e981142b24298ac5a2edbf66955e005d8dee5d5dc771ee753fc52909f81801ad8dacdafd2ea12d94b766ba9ae14c5b7020b11b81d87f6e56291a9d567f6f159952d5c10c19c4d2c21df8e63c69293c356d7efac7f2a267d50360e06beb61a03860c6857de0e2d242061b6d025e768d3becf43ebd802ad30b3d7f0f55bf000a3a09d52e44f357934d155041bd06f143f9b41fb5afdfd8707b284114acb518b6ce6de7215ba45d47be19b1c648d7618b798247bf6a7f792508b80337a3fc0fadd3bbf616e43e8b17556c6b6475525e5a84ff3402fee4a5249f47b1d20adab56ecd09412c469287a62379e25ae0141ad55adc038853fdd9d71282b1587591762f9b5c40123c73415a1c67922032aa7748af9a93394e7d3698a0bd5dfda5bb5daa5e72b080f1dd7a4591af695e00959c4d4581815049695fd3bb33edb4afef43b3d06ef0afd5284c2f5f4ec06f0f1eccf111091a9a7aad9615072544ccc3de715b3a8c7abc44cf77838383cd66134da01e313b5e3ff23cb50abe6469fda62c5ae95e07bb30a31492951eed3a4d0a3230488e7396f1aa30b6dab3c53cdada18a8342cbcafc68cbae1ea539e7d50c411c63e45abd8eb1c5d947605bff7e4010ae4b6d0dcabbc101aef13f55bfe2ffbc7701c8b0d754c971ad0ef5cfd5c89bc847cf8470335009703a9b56f932b395d3ad0534870d9b15b6cc7cfe0709c2955157d87a4c067fc0b6e4bff51d9c4e334387b3702dd8a31f9ce7b73f7b94c9524097bcab220c0d227ab0f0c4b283cb18bdb9487508a9c787efc5ba9d242f7de03669a8c373d602f9bae9a0c7a79fec28f84f874dfc4b3c9060549f6d601940d005e5f1f7a14a685fc034810d83b6f331ae914e069654cbbb4fcf28710a6b66a04258bdf029a787c8230d9ba05fabd162ced0a471dcb967b5f0e6cd132a5ee1725cdfdc4e39eef82da3f829b5ba14d2b6804c58230872ee59c5027957a129a0693c0dcad3ed508d181b2b1f9a1a81b083f5d0e6b2822ef3f5fe3fa48d284e697e000dbe21c50f567fc88ba9b4ca6fa2947076118dfb51bb11d5c09ef550b656854365bd0af38a1b2cbfaf39c1c5aa1bd658e9a11d921e841b141504c08376953b835dff652c13e3d8c4e9865255c6a6555833c566505749c2354ecac393296de0f5e34e416b4fc7d2d5f3bf2568438021bd261617f8029f513cd0ae6f35e39c9a07bc3b24e1afeb4a94ccb7e3d88af46f4ca990fdfc763e2ac03be76350f4a9ccdec1b95b5dc8fc4393a6e74e8697e5d09649a97b0585f032084907ba87745f8d5ff7c1474b109a4f577d184bc0ee2c78375576ffbbabb42d057a99c09cfd0cb266cfa37467ab48a2fa999ba576509e5e9673f5052e67ff24ad544752cefbfea105ebcd6c609cc6b484802985bcb0dff15d204aed841eb558b8e615046158fdd8435166026775b3d69b4c658d44b49307bd62225a2978b0cb1fd46fb6fa9c5910955d638c5df7baebe18aa7790b091056481f4cd1cf0322014b81bb9cf8558232dfe333dd8666b33eea630a5923ab086ba72eeff65a2a7a772f44d47a49a2889f95bbdede82429177e7c2e0eaf087cc1231b8f6383352243c55d350a12ff020d13141f19b1d6ea1cf46956b12b3632ef395368bd90061edf1be6a1afd6fadac1b79aaf51d39304b21696777f3091163ff7e3526d63fc0d1fc3bcc4e77789a3b012fae32cd27746e570e61720822bc335f4b119f5e5a4fab69d49f46127d43a94b3ba27fcb38bd78f88f92b14bd505f8249696d92e0ceda3462c0a2669bbd7b66f6d622b65c60a31bc74c1ebcb7856184eee87cd32ecf1d72951441c577a63ee5b5b46c494fcc0b310e61f325c0428d4033a26e0f4011157e8c37767f9a2432c95706c5e6ce2e7f7a50d9c2a5fbd39147c60ae5ede7740b2f40d2e7d69db32cc6bbf543b9d419e7be2d3ce382b1c92d3b3570d6be12634da1c680512caf388a25b2affaf886942e0b1dc33aa554cd5e97fa53a3182afed6fd2f1af4cf08a72f9baf83a72218f8471d24a3d00f34bad44527f57cb85dab2c2a89f06cddd51152697c5ca4d0d226af5459a7f78e8aaa94b6087fed333bf083a2d5edd6eedfff8f9de0f9a3506a54a05cfca59aff933ad038d206906da77dde447b908bd95b926efcbf34577136892cf0158ef1c793b2e4f6226e3d2b7f619cb6db0db33946f21c0f4450548fa002c885d948b1202e4aced5d7442c8451815687c83971cd3e9e47b835c77271dd66b0cd8b66ac204f951574be1125640bbd996b374bdc76b015748d4d92bb1a6047caacba1e764c1cbeb4785dd64dade53621526c1c11d86176ab084dd0e59e4db577dc8b043bb35223c86dbb7b27ddd79d8b81d2a0aac70c7e4d5dd15f0542d7765d7e9b9fb2c28c50a46c60c83d45b789f9d2bb884f13c35d0362da5577cb2738c132f20305c5a3a00ff47a507323407dc500bffadc84e11733ec29f5ead3d04649225232003c20bc461744ad8c88e7e931412cce8a0893ddd67b6e0b64234ecd3a4f005903c72b56703464af3e69a1e7a3c680247720e08fda2625066771540467f2a01fab609da312dad78d193f1a1145056f4f76b6ea87154595292e2e11205e48a9beb469922cb3934de7f2108b38f5a0440c7cb897cf9a8f4a11859b5fdc4b0a349dbdd157237d753a5a910500f83bf7c22191f6e61f202a59cf1edb2299c805c8945302c8713b6258974e38f945e4bcf5e2691bb43378df009f614294e59af71fbfaa65ab133d90cddb7dfe05338eb67e11aedd9fd82d582b1fbc5810081679772a99447e1ced329d876d933d267626aad35e6d7545e94d10120245f86f0af92f22b9fb21546682f322cb75fe7b1921099da59f13366ff50fc8cffc270fd1ed5d5aa29a80a51211fe646a5a9b00375ad447a520a3ed53cfa66b0456fe56f469270;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h425b2e269c9ca9a9e0938cb78e3b3028814838767b1fb4f6453f9cdc6681b02bcd57e6188bd5e360ee0945710de840af3ec72f8f03c7a76203d8d38c66d25be48faef8143540590c6f0c63a141bb3c09a4dec25421c8ae64b913e1525061717fc8a62e17cc06475ced83ccb1b588de8bf6b4af5469a1a2ab9b41847a02184af78d738eae3beff916308ab23edeaebea1610006dd28144d4e3e43efd87f6246045d2f444f66ff804023d04e470a819fd82330baf332ed0eaf6543df1bb83aae6d28e4087163c7554f0bd4b9aec5a9d982b204fda592086177f00489b9078fa1386ace3bf643935e5e6c2f290d2df06be70dfccf2a384c6fb23868a2862b210c5c04ee74ca84747d461538e9084a025c2d13974df427317b1fe73c5891544b63ea19209c0be4e5c0720d4f7345a8aa25e57868c0158475825e4bcf4f73cdc1e40ef34074ac371b4f10586c717b7c353e5733dd61fb02d5c866153c2e22c979c46ae9d16c2016406289a1b20ec7a4c1041d9a4bbff87333684fbc05f0024970789a40161abba97067d1b001ea076ad94569f9bc61f3edadac478ced63d717d2a929a01e92153a2e98e54d7227f8de96d6a3e74040ca8db91f7342c5f6fea1e8506e1d147439d0d6035838351fe4db0a4fdd571f7afafaf40d016271b6af94f5b8a177464a14c6b59e1d3b0ae00dc78c737a10e520978879248710373c0402b5934015e02ffff5236a185165e958587ade7a7b88538c16234b671833bd9460b64381ae77ce39eb190b8be4ae114f243a703b861130e9cc177ddf9c236f6bef21a1ab2f27c497417623c57d6de75d89d7c27b62f525e600ffdfbaa1802d4c1f134b80807212c16c98f9c8ed5373ffc6cf42dd0577b751e59d3fe9b3b94bcc88f44b723de644ca28f4c159919f75af2eb31c315eacb77983f07d5635b34986111d5fbc06873a22028ef9083a4d74f760b35902b5d8f56dc492cd7d4313d49a79c7ec95e5ea1c7c03d580338d86d683e29dfe849a0a934bcba35b7ec0d99900821eb6232383d7e5825e0bfab637cd99fb9c8d9fc0b00cc4dd9afdac4fc6f462becb6ef58094e9f3a4d498b606f3caa4027d135849d33fbc97163c9dc867ed1b16af47865615c50b614575267e97d946b83797bb3c83a17cb8e87304b73217b318c393ce0166485b81664074bfbc67ce402f7d79545ecda97f6f0e5572981507a0b7165d25cfb77f3fd5349698c77a901b239a54eb544d872ab8b887f06d893e4dcb61126a1c1467f61b83269ab433a15e2946c47c1c5ebd1ef870f981780cd95b72ea49177be079544cbecc88b3e555daece5191a6213151b4daed5e1952a744363bf0993b558ae17897df99d638224cc6f2a767cfef25da513d9cbac40b7a2446ffe1a5791cbf0cae1314ab2ae4360b813e074a716850fe550cecbc9ea9524a1d056861daf9638f015d39f1696b8feedda0938c975809879911ab11184d89d2ccd8d3e1066831cca12482747dc0f062daef046e0bb0f17d2f275b53a34b1b8cb856476084fd3060dcdd37a053ee859d2f69780873e5e9ce061d90eec82dce55e4a2df402862fb29a36a5c0e9462df2b6bc3e2f5b4fc6d8ebe0ca6391987a24e8844f3ba42c4d0f2621b903fd0c6b4950c97abd72d19dc0270f7bc84875d3609c3a2fb91897ae0b23d089dc7777fbc1efea8426ac68ab114b8c7623139db898d5f0f470b34906f9562f260270deb7542be2028e180d5e8eea00f915053e97dccdfc882df2571c69f577c2e50a4d72323c8288e36f8eccfea8a7d46cd81f4c0e80a75073682f526f798ff5b669fb2c1a918d65e76e83c203335cc0e6acef19a8b39b7768b7f8e47e5516f1e0f6e3933d612e8cb9f768c3d8cb97e16475674935c82541084c86298ccb22516349bc913f758b531fd848b2397be3d56d9948a9f6fe33e3f2b4b2c079744e92c22f198ed25ad3b6995f71a8cc55e02e6fc7d64ad9d25058ccba8a27152ce08aad45474a09cc8c2cfd8930f619ab9f8425951e4745f205019b5b499eb61ce22602ca8133f8b0894525313e3378c728f513f463eb4879bbc0dcbca450e85f52a2bf5a3f376bf7edf0790322f0af36457e2a3cc415f43ceeffbf05cbb7f87cdd81b7b4410697e7d22b5c3875c6e710816edd3d1886bca09b97bdad7df43b9d62b26d667c8f3d8b39f1dcdfbe409794856191ecb44df7c976c0d52017f811a80d7b720badb7b4e2c5277a8cf795172b09297620fdcac527404c3d02ef7f77428092a9e9e50fd4b1d77aba8cd0d1689ac5d4ed1cbde926f795fa82f8e53945a1d5d185647527e221b58dc84c36ef75801d243a7a9c8ca1cc7bedc3411af57304da4cd2ca35ec08b39e39bb15be90945e21c59c54b1229005c39c2274f7b5a958d38f5e9392ff7cee95429eda0e4ff06c7afabdc1634765e0ca87dc724203a80cd7a7fa6f991a2b5c5a1840dea11a65c100b3120d5bca5c8432748c7f251f4ebb8cc40be523f6b2f49337d9a2c3ae2fb837265ba4c3fd7676a5cb4f3cffdfa024ae74ab07ca2fd358f94377c0e058ba02e7e5a2532ccfe30fc47b3feffeb17e7905ebf7246374a0400557cc3bb7cc321a912148972f42f20142b9a8cce608ffb04d71c0fade750f90bd6e81778705d4fff7cf18bb247a1f82ffef06f4a5a9152eae78a0c799e9b1a3ff37a1946d233950205917dd72bd6c9e1e3ebab6aad5f7aba3b2730d24bb2caa2e12191ea7e4769da4a9ceb7d26723fdcd18cb595a51de6ab3eefb4c3cc5ee497e755db29e5c5c3ff59834622e3320c1e65b0d3f770e505593f8e918b23058037fe026f050a7d22ebd6f0e03bb3aa306b4ae7904bbf69863c3363af0db6b98be6aa0b4831c75ab1c27dd654e52a3aec2a0db7052a526324b136b994e43d5fdc18b41a073ea8fbffd5f86dc6cf1d27926b3c87c5b7b098af4ad82f124e66aacde6b47280b48903f699927bf9f8a271fad1c7d70a57a6d143ec44a0a2076c91331965bdea4944522b2ba0731838a2aa1f36ed4ddb1767d9cccac87c7b73d98b93369db1b2d1416651c04867107c79fa88bf2ba6fbc3be38702895eeb36f6061934e98bbc50f06df2d14dba48f68398ce5667ee221a6a754cc9f53207e8fdadd65339fe7552c2f89cfefe37e8d83dcbbe883cdadeea72488a64940e275d9e3d31de3c1d2f2d5aec7e0d3b04f2da111f433a8c8866d0011494ce71a6111857740a6eebaa3f2217f15456a3c8acae467804997d5d22923623ccbad9546b05c4fd5d32877e334e6c79de245ef4ac5d73b06d039b8cfd5dab7f7adfdda5a899a48514eaf7239617c68f4ac1e23eb2ffd920f5504aa15ba6c859bb768e8e7e42c61a81d3eaa61f4b2b6e0024511918a3f1446b495ff48db9459e15993e4ff25fc51c8d8549c609bb5e672b15358018f9e656f7b2279cf1e8d458791d64788b36e095b4b2b82568b6d72fbee4e514056357efe4d4bd3c28c6bc53e8d440c387142a72518298d0958e460ffe4e7abb907e00fc52587540d75866706fd82bd0920eaeddefda9a07d57209d3ac33a4c87356c2b044c1e0ac86f714b4dc5366812b220dd22a6ce1a4fe7b66b97420f947d31646a3cd0a0a57a4132a7f8ef394853a2d4e4bce03002012fefd47a5654a609e3e050bfe591b8be4e497a93d26e4c1286f193b814cc2032426ddca9c74f90661ff383993bef0e0d6a353029aa7f85c70e8c898f03e2b9f9c22e70832273e2d37955dc303f02a845d847605b09de810071b1ebb601fb957831244ea82f05e1099e85d21de9a0dd46a8952e790a91727efce0cf4e8bb9778653c8183cfdecbaa5ec88d55ed2c20a690146d3151c1166d74d966e2d19fb995614d65781872d2b4958593d4421d5930835d65c5027762a941b05eda91adbdc033a6a9645cbec6e67101df41b14f6a39cc196045e30d7dcbc15c8780444878ac1daf11d90335bba848ce4e629dff74c6f6212eace290446cce53d47362f6488130776eed9b295e73f23fe49ace195f8c5e34df6d3a36c2146ed7eb8296628ecbf8ffe55f1fa1db11ded6bba4faac57056904b1704ca1ec3d2d9f6235451075ed091935ea3023b7c871345de88c828fdd6c4497d8c3159c9a137eb6ac4cd8be0330e8918f5f6c18c9ec62a76e274272228d89483df8a88d2ecc996cf32f541c338c2c241ed92c99a0fe3a2386af50b82ad2e12eb1165319277e8e5768e6e6fc2171c18cc63d0d1a91580c75934752e61737eb24fccba7354e448ca4dff94341310f536560f5a27e44ff31baf8be1d56b603ad6ec7b6739f4ca7acedacdd5ae6e8265f2c65e9dd993c5696836b855f5fc271c1737e9c2db4ac035dee22fe81f62bd4b8647c18ff53a0876267171bbc5f26d2479e55c0ed9fdef6835bf4c1892f5845a91940a307fc3dc528ff9de1036668b6a593c9594c6a70dd4e3da8223f8b026bd158261aee86b1bfd4ce887386f2980cc40c1f3f263b5b1c80630686a6e09b7eb5333a61511bf9df0c36fcb916cd9303f8f5b239372e72aa0a6df2d5999c2b3e9265595625dc28fbece10aae27851cae36dbb39f5d75b701fe688d7244fa6554efd3652d3d5fa3a4fb33895da2dcd9a5148b04e8a2ae12be56b3e554ec9afb3d84068288210ea48963da538744920b619ba6ffdea4dde7b20a1426a9267edaf99c62d221e35dcc9449aab32da7767773a11062b2b15a8abd3eb6067298be0c41c7d7dbef212c86d172d80692e764d10610ca4fd48a09bb6f75065cead60946efdb55ba9bd51875341f7b0e651420d24b61e5650f2cea3b1b04144ce54ed39151eff73145b3ae57a452720ff2af9b4734038a63d088ca731e970ed4fc0255d9416ad2752a9538b2d1196b9fa572f4917d91380c1ddbe0cdd0b7350ebcd28f610860f1d876560acbdb9ce0918da9da60ee159696d3aa97b71ccec63b3688f979d7f478e29c882ee4a8a026bd3a4dcd48e7605f79bf30beaafa3992e750486fb9cb40e8ffb839b5460c6a342a704d07ea68dc58b3b5e440e25e1a83afb272f52c2433f834deced317e08ff8fb1dfff38d04e0c61e89a092f2755ef8d55584d5c822a56695295fcbcde3abe8396ec3f4c09d0033c450290b91c8a0016e5a785ff1a0f5cdb976ba5878ad5f97b036098929e68b13e54cbe594db186821f135a66f7d323ab0249d76b11b71be4818a3539247e21b1afea556313e316e993ee07b6acb1001a3030050fc3fd027879b61b7b65e338cc48179c2056ec87cda4ad98353e2a6ca42f8dbe499b7be3eb4cacc365d790713a704dab6f2847d17de6435144727818b86bbdeb188b69044186fae652b569adb6d75091395d84fcb956e49f87fbd695c3fab42ed2c663e7e6c92952ac2ada9827bf146bf2cf4f412e8adb6d51ffd8af03f0f40df59c9ef43517b91532e547bc75ee0afdaf9eb4f9aaf822366c204a18bde11d8c1fff5233d24102cf3292749380f9d7274050dbe385af827e3bb74e37ace54901b4738ba974c396aa46cde5e8983d85cce32fc50b22223e971d1d5cb4e6388252fed5262b5c2f34dc4ca4aef7816ae9fa07f1ae2296559a60bf85e2243ac988675912de2c0993374fb7a1b0676f9ba7c20d82721e076c81b815f36989df64a868ac75ecf282426140fa5ab6de5f984a725d6003f13391232e1f03af7d4a7e314aebafcb9778baf329694f03fb0560a418b069110f8a12810012bddaefd9c612ccdb028f28016883d23cd4ca29a551705ddb04f931cfa45958a337e10f2d797bbbb837110a0364f4373a198;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd82b02a91e523b4499c0cb389518f2c10eae444357a6df7e96e5e429bbb97cda854efa2a025dc84ca38a284f35f87e3cdc46f3db364474946fc94348e7cd9442cd68a09b2a23265e78090c3647a7bfb2f3d19d2e4887a0b7fb56e0fd86306ee7db864fe8c23cd132e22d5aed00f30bc3cc20016be43dd0461bf4e1ebf914eed5475d692d891f35ed6e134362b008660db968c93f549034efe0bdd59106784ae1629634a63456327a3357d8eb37ad66edc4b0810bf04e4d7f04813959462adf29ecb619306c605e43d8f107cafcac330e067ccbf8deb78a9ed3a132403741b7c65d88e4f25724c4efc46bf14d3d3c64ac3e423c806f9039f33c33eda1d5b070d2e23ca3c7dacd5d6eca95995bccc968f4aedeff97625143561fa7867de41f7a89a263f8f64227f32626f6e9887af9b7e21432257e6d6b657c7e11079d62b8a653363d77bee1f6bc3e6a61c46cac888040e8888dc96ceddfaced3f7241bb605b599790a3a2dbc04c8bc89a87401cb275473caaf8a003024d0c04b0b77d90eae1c3ecd9f0a7382f62932ce23d42b2b3c48ea0e879b02d4ae1ed65cab47b74854c6dd18b950310d301f383fe5c9467ec0a3142e1fe72a152612f591c865cfc89891fb3eeb3548ed74b7921f62a9d906d114d011d5345d761ca38a10e952fd3e756b9862c06ce30e960b4584c500236723727adb6a926f86707483d3ac896c1e3f5e8656b81fc9d71e49cd0325ffc98b42002059e9c40c44e322612708590d21620b81bf2202a832ec54875c2293138ad7796efdc562c4d77f9a969e04cddc26c319b5ef7a9934e4af7f3a4310e441507630954591194bb8404c64673ffec2868e8bac0f396684e3283370dd6ada6114ad5e8cc34070d7b37c2e802b02603e0bae1c1fc631a2840474c1786afcefd41e45c1dce69be47d641151f95926baae3d763729d8c1c41b541559daa03e221ba543da1bfcdf563694f99c3dd43b71a902ad1a9b86f16597c368184ef508ff93948a72257b534735d35d1674a463a15e910359d0e00244c191a16acc087626e1bfdea14fc395108588d06bfc328c75c2573999c1cfdb4bdf83881a2fe444d65c01185388cf430e557941d4a24c9ad3172a647e8b42d25d808c95964ea523575a99da645cb30f3c606cd13432b22bff4a3e9ad23e3b294197b1a7da3f0087ecd06fcb38bee112eaa57d33cc176adb45bfa30c169d02f89e7e6b0f497db3750b1dab2dc6b4d07b36c87c72dcd30444d27c3c1e0009d0e7224be02ba2182fc67e033d174d758f2ce8d345c60b75dba478ba9e20c32b5399203d9e35cd87588c388dc7b5aaeb11cb1d48dd3b4e22f5f0ecf8af36e17a6b4be68d18017ea404823c5578a23cbb7efef92bd3c732ff53f2b79ca95ec052b5cf3d97784052e09dcb61add8c70b39f70edecd73736e85fb2633fed8d8b61d2bcaeabee4d798122891835bba357ccb86962e4afc8f5501545a62ebd484df7e8e951dd5a80fc5a6263470c6d48521ed01b20da6b3306d2106435a0b9ccebe3de95a8b2641231a2d79adcabf99e28608e45bbbf7ec64760447bc1c28f70f955f601e4fdc514fa2f7862da9f7d0be50448273e2818f07cd1f847bea00e751182e9baf71bb6d695f7a187bf1dbdd0583c4898cf4a1b50cbcd9e40772cc892b982d8edc9ac6049fd60605f0b7ecee70096bf5f69f27cb66477eb5bb510d427c237bb73df9f5966c3f23bf1b3f4a8fba4aabb24adb51fb1f2013ba6e80a1db785a09b162eba77bdc85695879dea561b0a0c4bfea6caebc7560301c5aa64e89ee2b94dd1a4a872e6c7b94ce5103620484c1d00fcf10ee649f7edf418cf89fb9d4c1d314c89402eb3f6bb76ee7276066c297dd70a81fa5f3f6a22bdcb27e0fefc162477424c3fa656f4f4d98f4da1cc29b6d314ff8ef38be5626bef0379921c94249958525400a37dcd787ca2d87b89dd1352f4306a1a0676156dc1aaac844aee4bb75e1b964592897546850244c2eabfd666af318c27c05f0398e192688cf0eddef8b3df09982750d61a169effbb468c9aafbde0e69b2cb926e3f9557f2a51693288ff2cdcca5d1e89cf8da0dd76945f579bfa685a74ead93924ca43dac490405ae82ff1df270d21b4a45bd462234a4a7235dca2ada39c06686dfb2d289f5bc3316c0c0b72a8b3d5cab6dcf4255f10f19368468f9f14aa2a41e48c47cbacd4d6b038e92aa56aedd4cc647a7643f4e1b40dcc8b07a3f3d1ae5702563e6912995e894dd1a66628a03c23eecc795eb1e235f9158839e1fda7bd7f723c4edcc495382f36a9217d02a20b32addc5f21cb748b25fb61168cc63a73b7eeaa37c87bc1e4491247c1a6c40beae9cf78033bbe54ad347e4748bca8a1b0e1dfc0c0b0a379af7586f988900866dee2469f42d42bd6708cddfed9b23374ac80bb21e058009e2aca39dad29b78b35365e891ef0ddb0e9f5fe0c868bd69a19cc741ba61bcc76c3c2a1de13d80e6fdcef5d4672d34c9462d1009a4a641a61390e70a393bd0fcddf37190846f059715caa4da2e7d60d07d0b5625914d095575db9f2f55540e4b198f18eb76c02901eab7e0f91bd2241869fe73cfdef97a2e8fa923062091afdb0b58e721d32f33ef8f874b9682a3f64fdded0b40b56bd672ce3641ea46c39fdc12fcaa42ddd8e67e22e5ba06f930725d8b077f186e5993842e0fcef13e49700614403411446b4c13abc2e5d0dd6b0e79b5b22664efd1f8fc72be2a058500bf0b758abf15c75f558f8e21d0ddc543c6cef855803cea1d91768e1d8dd0467d6880b2bda00a82830b9bfda633dd3848c1371ae46b1578b8e24399f0aee479cad94cd6df19b235d1953294addb0f4c3abd12c9f81fd187b5bbbffa9c92a67fe331da833e6aab02c561dfb16caa333a8111c043e6591c65417f50e2c92ecbfde6b339344d9ce5977db5f4b7887842d7741e47cb12951ae8ccd94581a3ae05c1e6817588ff3440b578aa80398273e10e82423c9303522144157f4bcca39500fbe042db65501bf18e06cfcb94be27ff5a3079ac827b51440b477282a16abf29834df13681453e7ceee312212f14966b4e4ac556909d0a4fa17a7a6e7986441c433b808286e9e156479d8d289de1f3e65d948e12321c706963e2208c3717b4de5dd12b1472bd7c8dd2fe850c3061fed09765b62de3573de39d0b9673e5566d548a2b1dcf126d2dcfd6d87ab96809f211971587eaa4334e8170cc36b76fa0188937557da7048e676528ff5331e204e350db8b6fd4551cba41300fd46384a582f909eea92b5571bd8e45481d94f26a3e91904cf8890d79412172b3c39eea4f99e4315fee559a0b7670e5e96bef9b6ad1bcf65dd96e91d7f140cbeff87efd7704e03c6720eaebffff00da6e698094ecee2cd1de52e26572104845876c4bfa07024dab209049f7e4dbe1fedc5682f85982d3664b1cea3273d8ab73d91bc393c5c9a03242b9d0815e6c77383c9860ba5e76aa8ad687d5cf4f733b2de2af1e2af61b9c83b2bb91335776c6e5a510ab1735ec1d90b42bfaabaa4bae99e374df369a08d578debe980d6444597d6d9e592c299efda9d3ffd3c64ca3424d950ee5e3159d37ffaa02b477fdbe2fb023caf72b99a5dc939dbd3d43f2948900ea0f8b9833c8c22cabff269afc020d1ad33b3c21c609f7a1bafeb72c7c8dce3c19430ee857701d71b91f6096159fab52ecf21322b344a5e14cf921e805f100f7fe8126f33e724772ec5e6d58f174b1628f1fd63889be62f15cb229cd4eebbc19fa429bf30f25efe84a9fceb99d3fc195380db78c9c52e8e8c0995047b1b923d446b78d6f8a2175a1f2c4df0fe3a1c642e16937ef49f4a68e62c42f0e77a9118984fd372f14d59a34ca0924954a9ec01be8390a8f8bee3f890c4e361fce3a7ebb9db7cc901d6cd89352e69b175e61461b9bc7f2630fc51dc82ee53f1773e3c5e012a4dda65e63e0194270ba23dea3ae5689c34ea74ce6e1ae7fd20f7cff3460a0ff596eaa6443655f8587f5d4acada08967f4c5171c45fc02a1cad5a8fb0705003087be24af611bd6ae29d5f729b877ee3f29ddc8b743a6b0ca3068916d7129da9322ef8e4bfa3c11c51b6005ba72f2951d3d38d927d4d72f1265741f083bf2d2309525fb79bdb849609134cd7b16a19431e30cf6448bf4c2f8de37c3db0818c1a4d813ba28d49d90ca9e078c010cd3d669b9b98ef4e77f8d05beeb39637bd6372c8dfce62f2d720306317742f57070053a62187a14557b4f8afded1f821828edff4ed8b70652456de566ba71d79dc1751f4615effa806756c2a6341e417b91c96650b3017139068604a62ffaf066eb4b6c7bd654fa868a3c910b1cb6bbc04953c31189c04f78b97a982359bf02b2b421202c282af891d3127202d272f2a3056d934bfbad8742b952e6e9b0c155349db7b6da1d5ea444cab8ff3e0cde7ef63fe89a0deae12310775bef9234df514ac1c523b9b6b490d1267c8b8a63b70c4cd7c053c2b6d071084a274c5259e13c726970f3bf5ad4bb40cf1baed0246f78ae935ece3660e6d31470131eb74c00d2af1e3cd1ee6735e2011105abe7c22c72cc4772b1fb7d06421b5789db320bab735c7205f2f6d066eccf2633084c9c95b10715d02a5b12f49f1351bae7c54c923eb639f5b7c3cbc1da868728e1e88c848c415103b025878dc7dbf08442e370849e11d1c3d3fa59a176799c9d848cb78195338f3366d473767408b22e5eaecbb3d85d39c049cb7a55feefc9b4a6b4c3a50da540e987b812a4d4119b48c75e4f594e2ed26e3d49c168eef1a5a05134fced846d8155b8364c678b3d80af668014aef09cd42ef7164fe25586183c1b509846e881f360bb8b4a064a304caead57b2909d89db3f951c20f2ac0f4a57c4c7e925e523c3c1d1422587aa02ebd82c41fb4811082b06901a8cbf48566ddcea07b2403634fd9ca0b3f15543113721bad83f58e65fb30cd07892cd96c61f1dfd22203e88b8a3a1b6c48a23c682240a9d935074c41f3fade422ee4f4fb3550ad8b110b536872d29d4c5be8f3cd054018824083afab35a8868a39f147497b756d26d546038b8cabaadbc044973d43e9e60dfb287851a4516f9fc5cc6390110b53286165f2179d00ca837ad11ce504000d582d83a5af4a5379e9070e8aadab23251f20533076ce6084c8af65998045eb156373ef6852720964e291a7b5a47cd7c36dbd9d4b9ac0863e9617377413a5ecbda9e209350ea0205f0742478a40869bc329af0ba921705991b559abfd7541226e7bbe20b8db3ba3078ced920e2afc841c004bd1a5b4aa64565131d65084d34e4e27f8cca2ed271af2909aa5e73b46b1e860f3419215f60151f733438f1b08ccbffece5b80da4f9f22555ce59a569c563cbd06cd535877995c9e74f842b8f3fad8db4bd35f2fd4f5f9e9f477d1403425ace98984f59cee611b202d768f58f3e95365678712a4ef94be52fbf85439b349ec2761e575c27f6bb584f2a2a863f5e8463787f9d1d585f27aaf970ad09f5676f2a8d791818a1f5fb71eadc9672e35a94ea808851cfa9c1ca8acbdb8d2c7a1cebc8e2ee9ab0e69da46fec39b920b8692950461144d24d5cdc9d75afc77999988ffa62816e28ab3a7aa6aebbf95bd8c3d9078c88837ab3d2daf802a0ede8b14e5d20e2174d7af978a74cbce00e0947219bc7e0abf4be0c87a77b99b3c8721c69cc0667a8af96de595ec96c31b7b4af7f540bdfcb9dd350655dee42142548d943aec2cd9a0c1154464c6fce5e53cff7e8b19e47ee22a8ef21;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1d523855a8470c43a79d8921bc4a955b1e5465296bf0a3b99fded71d74d45cd166f54781facf2aa2600f025503ca08e7f7214d6abaebc2d687204d58511384b222d3f7aa80ecbdfa1621b8cbccf0ef5bfe533a497415a7635280344063a4d12188fecb8b5b7ae66b0a9baafe933a449b6271ea2db59cee8edde9201d4d7ed31b0cad46a40d7b7164af743e495fcf973947061db228ffb82aabe3eebc948903f4c46f1f5d99e0b853ac9abbd01f48b8e97e481a5cf2e6bc700f892491d81c51a57424bc12d2ee5ae9834bb1769ddddf73c6991d33cbfa57f5766c3808d703448c39f5d15d159d6a89d52c6bfc8ec943e4b0266fe49d43acbe907469da42eeb53cefeea23d7cb0fe3a4bfc5df1d4533498abd2bda5716299efa830087433f6a1fc8a9043c3d9a309224c5d2f3946feff46676e1928e64aa1721cda5d58e587ee0f4ac118791be2386be45756c58cbfb88fb084a8929a0e7929d5ec66e499195a777e7279be3b51a0207cdbd33bd9ced4deea33909e8954a8bf04539a43c1497f3495454066508728def4f7ba55a69fd144da3d9672bcfa4fc266bfb78f5ac559f9c50dff6634918d84cd0892f4a20f432212f42f5f2230cb42e7c19f470b6bf15ac8eb625293d75bd8c0924181b229d757fd58584df2a3ab0502814a8a7dbfd17bf08fef2918433c59562a219e5e3dad7c04ea82dae73ce29daaad16fda75e786c35ffb6f2235e494e85d905d7dd9653e8082b9e0705ae5e0aa5adb4815a96fa50b2c9f11cb554a59daeea1b53d8cff3bce3d9af42116e9209e065617af375a153b6f4b256d6b89f1f1b5eabb163c7960424653d9063b186d753e61403efb29e6f5198c73f683fbd044d07da73c547bd4daa39e9941fc4ee7c690275372ed8c2b52ef1ed93ce42015dd1fc5fadfee9ac1f26a757ce3c74673000b3a1512e1a1df3c0a4368c8e7893a4b865a227b9338daea4c86b3eda09ee144b5eaafeb8ba9dd0f0904ac3259bfb55d055786dcd815e5be697a9b7d1cfab32ec0c2a86b998fc01578c6fa3368b54e4968c64cc501298096ed16378fd37182da7cc3795b6ffc1e9ecc95872981cc8cde5000d30dd09b6c5e38e6a49e7d8c3faddbafffb73d305a1fdf114fd90bb12c51cf448cde12c56bfc8307599469be158d857493b771cf21ca5dfd8d47e49e44143b4dfe0c6da4105a270eec1306963bfa4e2927db53d00a626a4f512a217a7c83b73d627b47ba3ef32a2fe4a04a1a0772b3bd9c401cfbf4e3fe32a8d219b029ddf4d9dcdb32a4b3f5b12a548a9ada61dd5552043256b7ccaa3495d53757e2eefcff06292601cdc527cda1f7a38e05ef738def0fd8ac2ccb23d92cdb409c39e14b4a77f3c469de7b0973890a002d66939ff30af278ebea051cd9b8fc6109e3e2be50e8799f0ae08cf2477489d613fe7951ac25203ba7c4176a318d049bbd78d3735c2adccc1a4ad316b499eec38e4dae9f91b18d14866e8c323dea3c8f728ac314e781b2c7fa7756c29340b7bba1467489fced0e56bfb83d45a6be6079614c49aa9fc5cc51bcae29b888240f0ef5417567dba98ea0ff644ff721c090514af2342512b23e10aa2b2cb93be6db8705de75ca6a004d94c64846eb6d4c334dae348a20fe6831c4e9eaa5d2c9fe2513c7967025319cc79f49d915f099434b574c03b0f53dd3b0d37522c9ad3dbffcec551694609d92372aedb20b443a2f088f4ee16e36268b7e8fcdcd256b03fc9b614d370dfe25d25a65aa1d25189e49267fafdf2022f4b8d8bd8e93727fc67e7e00d207a7648f6b0ad2a83f3dde4fadd08b6dbd2a261aa54da1cd3e43b6ac7f343aba2c448a9e5d15c37762dc97940feba69288860df878fd27a207b64551f744897475ea4a4e0868275a0715300e16c89fbbce698eda6e065011e97779fbb390a07b21470811a58f798878e420af8c99498291d0ecec0848ce3ec283cca93fb49881acaf55d21b867b250814bfa211aad354475899751cd9c995a9d413fc2df6745c5c1b44a8cc77f4f24c1f7983c5777239b0c6a476588c60cbd7df803db9ce8f134388f3257557b5f156feffa3c9dd172e1c9283d43930656aa0dbee2a6a8a48f353a50f1b3ee070e622b5c5287f4784e0b8653eccdaee556e175fbff0876745e01c7940207a72d39125d959012281aa216b7b4899a78b6f05858e33bb184b79671b0a879f258444c04c2bd22c05e73e3c2dd5073341925ae285ac92b0a370572a573877b8df84f6953e4cba2eff4160440835afc0646704d9462e2691b95b6a447363472b697aec98be7e2408b42b4bcebdc0a8961672fd1ba00198d1701f810e24ce5e8ce7997567eaac0015ce37767311ecf25490ad097e85daafc267a9189b278fb46d388199d1faab6826851f2e29f776244908d225a65b77c9b2d244871792849a87b2297dfac2158e59203996364e8498a0a8a718a4c6d12710fcf7d55cb0e05ebf7df39b1ef1a47f4752f7d2920e52dca74ba541ae451cf52984c73456e30d681eeecc9cc6b238b53eefa206a6cc22b5e25d65e4b239335b03a36eb93e3f0ba485379aae978794aa312d9d4097293e6d8b31e00e72d4d53b14a723b2e7f37fbdafcdee2ea11800e8f2b65a7d7f3aac6a65a8762bfe05178219542186e99ff29c055a726d8175b9a7d789367b222fa3e5acab5d650d7b5e45d673bc2641bd29b12ee5a65c8f1afb514c183d16e7714b20be2992827723fc454fe8f18676e48eaf4ab5661a5c7cd647cd995f4c5addc2cc846fb0ea3893e6df81e514722b6630f6d6940383569630fc37085dc0168a6f8ca99042bb9bfbfb1e5e02cde43db1d71c32521b1d1b9e6060e2f8c11737501a00e14e4e715ac3972369c0fd137078d1c8f9bead3aa8516a603ff974495113ec5e371dd1e01edb614336c57bf731f742158fcc2e2d2f9b03fd68e935d1a2c99a47cc1798d48d69b219dbabbb9d76b9a6178a7d77ec79600e434421874af7d8782f1f41b9b2d1dbe34344609d71799d7a28cc68cf74f6b0967b951b1e004e2bfd6cba63418dedd12318f63f71ad2d11a217aa9749aa42f310155f2f7317538080e19113b1b336a4f53ca3ec7d08484f8c12be926cc4b2558a6d9d929d4844d28f48e01e1f53a355ba60ccceafd09b771fab9947baf451d08d6a03aa164a190b7a290ccaee61a0046905b964237d75a4fe2dd661514d16de1db4b6e7472680c8ced84e8bb322b10605605068b4ebb2830df37c9a78a75a4aec79149abfb9265b825ffa32df11e51c31c4f7c9389196b01cd541bf6ca42696d0cdb24d869ecdb32c0526f417135959a19524fb004bdf2f7a390aafd0cda569722ff8500a68d02aa5daeaf1b308e56ccefe20e7261af2c0aeddc2eb787206254763212a6ffbf4b31ba4fb2af052637ebfe0d716a78037df7ddcb0239299c4b6ce960b119ed1ea034e66fda78f0452b04137cc8e5c62fb2ac0d24230cf2ba03281cb708f1608db2eb8ae80a53544d07032b932c4506d53f806560c5cfd48ae063d138f1ff017054f5f4b062ca34498177aadc800dbbfc0fe3362356a340700fc1505155867d38f5e19dc364e5f5a4d3b4f5eb3dbca46cf70a546c5c9ec228f7f23c04467bce9fd2a67929981b7e254da6943cada3b4d6978b6e34c592876cb5f18dab0c9a3b2a4e2797c231d8d2094360e03e6a1b56d8d97e7c95141cb50cd1e11b76e692232fc6aaeb29f6fc552e29cfd82a5c12c383bbd3021296386d7e06d5071996c2cdfc6455fdc3776a155633ccc5eccde809b6c4aafb516b4d79f08ac447f5dea6f20a7eb8c29bea59fa3a3ccaa1c7d7ba758d3fbda82d218614a408340507be751c09cbb18a3e5436dba39f1bd313d4252b00823e1b91916f324a7b09f52b5e7a9649db2dc05ba0749d6d72c40ea6e8cf67d236ff82c82e2fee33ef463b8587bb041e87944bbd60aab112ea62d917b0746d871a702bb445a6bb8ba426aa67f585a918c68947ff5123f67814d4106be1759040d26fe2d03ecbcc272b1fa7d83330849bf69c09c25b6affd0091acf337409e4a6114190a3739e63152531392cae4b227f8604f077e6d875f90b561122371a2027a318ef597f03a9dfb7297fc444ba5c2cfa9e2a6b0509764260c6aba1eeee17c19e0de70c51b91f36f3db0c9c34ad1e4ea862596d8c16a848f7f44c4c70a9128e6eeb46d5d2efa585ac8c63d52611128ba7f8a6d860c521808ec75d688d174c558816ff72ed1c5d1d549ce02cc040be3e0d874bd662e5a8c4c81ed57d9cdad49fc814ac4b6b709c3805b1723918f5eae006fbd60312ba151014222a669c7bbf062808fe7220c7b9e5774da3bae780d210da7552d7a216558f61b1d09bbd5a38e701b896d35e857d946a3a3d0797e59fb5a95e35401794f7348967b49afc9d8aa3fce9e17d476bf757baa9c89d22a7775d3d0802b508fcead96a117eee42ac4c657ac9e406c03f8a8a3e2fc2c67d53e415b1d3cda2d18b3badd141d33cb1df496769ed8e82e7be2654ab187824a6b1af9a0f3aabdba0a18b91d95ec0aba88157842fd561d0f70a1dedea1414c421deedc78e9087d931809ff56ec2efd9349d5ff0dd8ceec5be5dd4c1a575dbef473ff45e35cad1a25d515181f945c847c604abf1a801d92eb6b118ed794f960954028561e88c3555e14391902aa4c78a8135a6ba3d8bf35c34b1dce94164951c975c6d9ae5f44d2e2ab1f67a687c4b3a8cb429ab67c18a5fe77d38763d039436173ab5465991fb055f25c2bfd67b006d7d67c568f0b748c24944d4a1b9e9ff995c1c6b03c3c75b18cfb6b63ee9768a07bffab1fd179e1da71f49ac44448aa28a77c33cc134e0d8f30f0f41db42e2ce9f77cb8a31cd5c01b0c53cceb28104000e3536bfc9a0a64f0fa0e1212f68a82b595e8faf7afc4b054f71ab7a6a0cd161a97414735c8c3e2c41eefe0f838511f33842476618c14a1b172237a905538ffb69f208379142add89cf958997ae2756f906c8abe336d4bfab057690dd96c9e28af308ea9d7bce34eb86e2ed5f80c0344e0718886cbbb4214c5d42e28824a211459a6a5080f452fb8eccc230243ecaa19a3ec945ba4b4064da1f5083c4879393b2e2bbba7733f0023944085bc63b5c1df812009a8bca1d15acb3d8537383c55d3ddc3649f3fb63f79e9724312779dd69b9fa9582e7dc9634198ce912bfea180208499bc7767fdd87dde577ea7d9677baae487b2deaf768b7cff2a8683a3e811dc048d268d5f73bc224b11d718e4cdc73b940c492fe336476007e4eefaff3b8cfe3015a4e89709bc5a28cb16fab943dc37ee67fefe070edd70c4739b580c8b775c9114fb5256ae0c18820a64624b694ce0de95d7a122732f999fe861aabb0f0441bb4f5a89489646ff12ad2575d56a5ee7b855512bb89c36dfade30c253ac115e1666642c079c56401ea49a968174a90886f084ca8996042f5e487d565294a92b0cce1daaf8dcabbb2b2e562c7866b758e98ccb206219d1f52cd36ed53ea5dd24c29f8127119cf82cd0cab8a8f9e549f05ea26a7c27c02eec67924a2f272c0b32a2ce0b31d90c904a1b79b1385080533400835179560cea947e713fab5ecc083f93b994202150c6cb067e2d3db66b801fa267d8c53f067271f71299d912ad9c67098b6cd55bd503a7d7f5f019085ad8fe2cd46a2e8cf09f887bcd57e885ce0e6b613afed721a422ee16858530886a37b26ae17493b2d7caf71b323b71c7816bad68d55c28f3cc2cf26f3fdd33296be767267c8d5c7507ac3058c0742f58f6fb215;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h192d0e8fa4d135502c8b7d5b4ac23e44b246e3f2fee23ef572913c6f67c939ef025e64a4d00f961aaf518aa49e3cd53c7c076e09b183c802f9ffabc0c42a6946adf81ded5fe6fba74522179d7e46b6030f7c649781bc935c1d266916c727ca64ded09ab7714b14a4004b13fdac9ca440382e923796d7484a9ee79c03791b714e85aa0d19d2b870daa385a3ad53e531c213d43fe9aa5070ffd7d31de9005802a2a05b62add049c97f445e372aaa37da7fc8b099fb349fce16369e5b1db1a3a44d8041e9ee320dd7a731fe1e8472a5653c0fff404a593d53931012a01abff144a161b7f6ff41d8aceafc657218d1e9f0e6fbf14b07f00d03094f40c99eb7a01154b51c461600af68444fd3e321a0d26e6bfc09e54cd5f27be2b779b6a85cbdd597cd1897761be76ff196a7324fcf31be96067762831895db8f9c11fb603e0a810ade91b84f56fca0438065e48e78bb3bd051d373ee5379790c51b618c822de1025da1a3a89a31a1cd58c001d0124a8194643720fde64ae5c999d5e894dc4a6769115dc6d478c7058b948047865c283c2849e7d09c836066d039981cec0388f02a57f969dba922001ece7247fbf10b80aac325df20f85eec608dcd06bfc8d2139113efa015aaee3abd853e0b1f10579adbc9315e2e8f7d863b69ec79ab3862cad0ef11540afa6febf6eaffb38125045b5580439bd2f860b7c8840cfe8d7a3186398c53e2d60aeb9b4b4dc270e8e63019920d7f1add8c75894c17f81916d8aceb64de1e210fad5c1e03dbe113352ed5e321f261c590ec7bd6a23a69f9cdaad381ae4f962e7c189de9874f093cc1326acf3162d338c89c7443ad0b6cec76e17930d6fbc4d0804ccc2486fcdc1129887d9a7f6e72909e8045eb9736388fd5cae007e9c5a9662f3bf66e9465a5f46bd622a4a2b09639cd9ca651c489ee2a427ebf998f1419d27811d1a9cc167b0e3365af66384262a61b3bb700f0cca1c6168cef87e72e2b99148c146b53f9b675c3cb149d7951d082490c42caeb84c053b705da3770024033801301f635e3f95b02c29808f2dca8111a1722b89348abae5b668e92f8c6d4e7f80a99818fcade9c44a76696652f0b38def7cf6e7cff339a3c225a81dea3660b47fa3a725a30e7da9eba8e0516b16a58437e3c6dc4ca6b99f666fcc8cb44a20b4320d1e67514e66c4afbfb1eb09c89b3fb068b7bc5e07e140c528cdbf4c26c04785bca73b2e78fda8d4f08bf4cd9c7c40b755b8b9fcc7da4f3e2e9e36fbe5353aa29b9b34c0d4b983ab80359cb0625e3fd1409a4c82d5693cb469390273d7e339f7cb4cfb2ede6d2ad6e72411289f932070c0a3cdd0d4515a4cc56f03051407612fdc090c2bf540e7ac11718c6fe85e5f6e9b75c2542f57170650e418ddace950f28006a0fa21b605a0a371e43fe5f97ef60c8a5ec347bfd6bbfee587b3c2420a3761bc5d9b572049ed78c640089140d250e289ddbf84a355dbedf67b49f152703197d4c758acffeb22cb82893e963e5b44efc39fae14cd2ae1efd453956d53e6731c466f41c263e960cb65ca0195953d973cd7533d2e8930c3357b74e7bf2209d9c84c622ba8f59e82d40310ab0e6f677c3a9efd714bdd07f5798a6f18211f849e00c48d5d74ccf13ca767a0fac1be27edffc19d4a6d843ddd71cbce7c1db81f6915d82c3455482a04cc1beb1066067b46e883faf7e190178936e5eebe879efab704ead9a9f2136abdb2286fd0efadae71b074d158b58b030448a936cbe2f35a7cd698ef4117a11db9039b4ae1adde9d0d144b060f96e1958c68c9588548a5b6c445994d78279dd621a7964c9c317c2c094b57152f32bd5ccdb89cc2b1d5507e38d5969723088eb4cda5075d6aa27a1f944fd6060c4dbd35baa5109d95cc5f24a21d0a8539d3fecd7ca2d8ef6bea1ae7d3a7ab54c77e27ef87ea2565f69485f644b1940a14cf327dee4ecd95801babf5ab7d283a611ebf7ad70fcd39495f84787355d4b59cfc1ea79e18d2a8e3ca97ad5d24339b239f47e6a1e48dcbd244c95da9e470d387f89f3bfc630d99621fd120ed0ea02dc5da6293dfec9b07383fb9eecf3839045546dfde3c708cb38619a646b7b062df2be20aa753a76808dbd611fa547e38341e07a9ef2690307c8567e865ba0acc51500c7bc3bd886b5bd0efe02da27b9df152dea272e8ed056dc5cce74133c2d2b82c82cd319add6bb1adcbd387cef5e4d84fef810d11fc2252ae95e975e7c778ac30b595951542ae3b28dc98419aa28e16efb32633679a8e7bb7c854f098899170e2ad457634feb77f99d3a17e1a53f193637f8bdd83e0259ccf1c2f13c47af3b05251b68b313f1fa8cb57ea873db4e569fc6c8e0394c7e0307396794a646e0244a336903ae078b1d70ed91d234ddea631e8506caae0447f19e56aad0acf486b1b6d366936ec1a0e1d5dcf21605acdc67554ae8b4a01b71f7ff67cbb47f3537efdbd300ef0e91fc104cc0a1cc1a110ec9c7fdb0a36f5257e5cef2676ce3c8651ce1b0544c756853bfad2e26c3c30692455a628f5147e6027e08d6c1a9dffaf35d79f08010c993678af9dc3a03564112d1eec2d24aca66047c28060dfde32618798014b9a4b8c10a9e6c88adb2a7819c405cf25372198fbace05032ba38b5a7f8e4d58923d9aea72b316010ffb45dc869f1754669348cde5fcedcb133aef45cc35bc0306a44c7e9ae7297e047a3a7cd8acd653a0cc0fcc163d64d808298d8c6852599657286e1b5f0a9bc2a9637519f13599a6fadf7750a34d1e8cb36fe153f6b541d955769392a5cee7f3ade08be1da01555d2441531fb8aa4d396ecab393e8b728c69ade91aececb1d8c3f1e5bb085d10b75836d2b1868ef2a65b73d593de65465291a53fc4e96b1cd05c21cce4dd3e8ea1fd2dcba9d8164d269d2cab87ea22df962432775fb4351d4f4f87fee9f6426bd7b19f07ba31673f30628c6999dd66f3c62ade8c0d45c838082568e39f2979b25c6f377c7a8caa56afa9753d69444032f1c7cb1dca626171c0316e12cfc0e72cc085ea43fe813398cd34441d7e1c3529964692b083e2e81aaeb974aee091054eb9e1d9c91048f4b859db4b321d4fc65c5fe612a2d5531646d5072758cd4a7bdd9f73c5557e7b1b7a417986a417d7bdfee6bc271414d8697fbc13c3a252b51e07b9c2dce2a26c3c4e8b4be2681e5ef62915e057f125206c21e3d74d804b92d1a45795f323f35637652081ea7fa8b22436898f8055e7cd5356ef268c8cc197ecff65b906adfe992983feb7f7801ae31f44e47b76324fb37f9d722a5433c10b2755f90186ac0a10bb751b6f54a4ee926d5efc0c97968e1e3e55d7471b19206e30162ce684d9348368278ba2a0704af433e076c03ad3fa11586f6f4b3a9aa885b0059c662a0e9d9e0b0273025f59d7cb845e1ed00530c0aab0ccc262ef9898aff2f2a42977a11d89596567ec584967d2d25ca4110925d78b36b11d2e1f2a9dcd9f0a1aeb6a75e378d946cf98e6a2e4178ea5301d6782c8c2c9a1c1bf3c7b8b5d397866bd2c7ffe0ae5f605f6046584f199dc8bc32c1a6b8715097231814e7aa1ac19fa06f632f9d9d2e2d8efa210e2a2cbe71fa232feff26c0b7e3a214fad89324db625397bf67dbeb2a305235fe7b7c7562557ea0f07b126227d98c6ec7e7353ff8c130842fc625e07395b472db2d42dda6aaaddae4aded01f6463f7678a742ac1d88d2273c8bc0df8df5a71e0fdbc9b8741d56c3b96386f4416448bdb7631bf9e1b9e146c5834bacc59682592d28a27ddcd9750ce7f9012a408724735cb03423807c7e586aff4f646f406b35f744a77c8080571f488289426e3147063924bbb66350436729e525d5626439d73ad3225e84d3130b96a42c62deefbf7dda9799ba6931bff9eeaabf631c4ba8abfd8ade236361eb7648939e70fdd0751c41d9026a7cebd51620b9015efa7676eb89dcb92054a6a5b3a98fde50fc6470d03ef816e7c78f54cbf990fb8d20066c5217b1b11bc2436edb3aa29a1aa21753a29a2905be6357e5af215ac2e2ba53921e5eab26188e1c508e3dcca25cfb84696dbd2fea8c7b9fc55f375a6453dd96ad25f586f87c49d3752f011a8617bd6ddb0d1b8d407abc81d24fd4afc7066cd2ebe67ae73c73817a7926606f5ec93cc0f67636f7558785a8845313df6dd41843afd8f3af0875c77a3fbfa920c1aaffcb95691de837b740f161d6720432331a3be6d5a796f7fa04652bdfeef8ed02c522ade9abadb845d1413e9c1e876efffc06e85f618e15d4dfd817238603658a8b37acf6fc07737b21bb8583f27e1de8cd54e0024748a47b755206cc3fe22503be2b3caac00228156f9f07c3c03bff24d1522f2fd369d7861d6843347c50802726a71529f36772f4732a1cc2a9f7b08857735ca012c650e48b2ff10844fa87e3d5ced6402e2861091b26a6c226a0975267389a1419405a039140f94c8ebccac9a52197f9a94b49438f2b194f554086f17f5a776fb8105c658c4ce6499cc406191a621b0589146ce9cbef7fc893a5a34c0d9e5a8f7da0f664eb56ae4a85121f3c0c52871244695da9f537aabc8f8d87a5a07288edb65b59234873637ac35d5b74846d4a86c8e07d25ec6feeaa2a33aef4bbfeacff084e0aa3f9328a278d7fb374b4f48f0e339fc39ff56074355f548ce0342a2d25ce174b039a9bd7ab38a3cc85d137dbe004ef26a34692657781d141bea7ba26057138d7977e9678e73ca937ac3b60efb13ea0cf58e11ea271bede0beb4a13a755c0a72ab9a8f3e478e4a1559b0831ddc945cc7e7dbaa38cbe04f5c499fa2d1acfff71d404da93f81d93a3180331bd1ad982d4a30dbb99e6d2d1231f13bfa92d70b0a2d10c0f0ed56e0bcccab756067b6032bcbea653070044b63a8e0c8ba4867980dabc824bcacfdff18142af162c8c5f878217d15d9da49a784939aa6003371d52e8ccd89290fa2623637a4515f5fa15cc9dc8c63b0bd53936c7bbf768ef0904b9801b4b599b402a80ccccc90d327797d39df480b38749dd4f922da0ff3dc67ec5a32ac779fd95d715e627d4d5d9fc944392baa7b584414c2e802194de541f83deff4d4801d083d8b8efc57dcbf6dafde351e592a09f926a5a96a894477e47407ba4e8ff8be7ccb0c30fa2693d6e7b80bda0771c9ee5339f92078832ad8ca97d64a90295f940b3ecefcf59802a3df40396e30816df051e8212f8e75097ae171320720b49468d59f1af1c3e2a60337be9a2b4b5797dfd65a0a52dcaaf09aea8d5bc167fd102d9fb12538fbb415b5205f51cece2529f818594b4b701d0213a9f88e3b157220b43006655a88d3a375ca374c8fee3bb70bf1321d019d741f04fc7ea76872a1bd740d5ac85cbda6c024dce9750d62827f155bff1e002091e571fcc858e97353bdd0b830b4ed8a3061d2299daadded92c700e24c67deba2a28be1691dba2d4fa7f8a185ec629bc5aedd6959a9a53f457a9b1a15abd58354fbc2caf912d4447a81b36c3827fd828719978ae81c2a9a563966fa236eae423f93e1dc5c86d945389562a51ebb43895d8ec63f6a5c11d78b2b06204c2e311f768d5532998c60f4e7e0682526a5bb3e5a20c97b8e59dcf7f9586a35aba86348baf979e2a0500fbebb329a9db95533eb7e956ae785597764d62ee1feb3d5bf7605ef1fa689e0266af12b172e15c049f6170b2f077c9fe4af3c9405858cfc5c9c4f9d0ad299b9f7eb906347a38a0d7b9e4b04e95479bab6b86e491557a83949606d1f729b31d735a0ed41cde0e0819fde8b1c4555;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h787a38aa08b2b447ea07d46b37f7b312cbb8cb6d9d5d050c3537769f0497e468f020439b6ac3d7d28ba2cf5ab04b71924a55c33f4712c20d8fb9a9400ba9b4b3c5a13435323491fdf0df802546c476581140ea7392cac35a64fa1828e461066b6f91edd8c26070443fd7f2c23c98f6d5b17f36da77afa50b951a11bd4325a817499932d1a9c9f70468fe33bb27e36b174c9ce5979d9db2c47ba194bea1ca5c0e06285c3480e3ebbb22de59a5520039eaf204710aadaec27d423b3396f785069033c14d9af47cf1ae373b6a810b0a2120fcf0e9f6e834dad251cb2bbe5196f79cf345652b35f023aa3e34824fef194338cd7a31633c3730b0294a24b64281a803fa19869f95d1a9d870ef15da2d56915a57c3fea1bb829d35924c3a16fb2f21a2ddb07f21849d86db7203c09334bedfec8d61c17447f5654b77eb312d82a59b1f93189f143814bed96959d7fb82028c4266887cd2f6c0ce7d14d4cf4e353bc560434b2cca573836a45d69300e8e4a064ca00441a5fa33e550dc61791640b7c5246c586210967d6be881ee23eec9899733abeb6e09e0ffd29a26a6a0f8722bf9354fff09683445ac7838c8199f4032baf60c973875221c94d5a7f81c4ca1a5f2e71cdcea6b1fc45431eeac7b6a8f1bdf9f163024b21d2a10c3240643cc50a054894f19b94d9b1e7358748163ca172c7aace69c0e1b26d88a91d131990831d325883a9b73a18f6b8e888e847efe7d09a25d316e298373b74dd74dabb7f2f4d4b656c2e5d06b1565201cc2072980399c13b792f51573a75565799a93b2d384f46a3b24defd92dc729de460c25eca73ebf9788309f3b20087d987076b908b66d9d27b63ffcb41b7dd0ec57c8cac1e62f9166ca8354f9186f91f138c208ce06fa79f03189fc275d9e730a89118321d24d4dc10de1d45404aacca56ff0b0b5876016220b22cbdc6df8a9c282881129fa2220c73d6fbef769f7bcc36535ec3897eadda1240829bc199c814ac310e1a89d20a41ee95fdc37b281e9c41d5176014eacc4c4da8430d311d2032c939dadd16b0757f1b2cb4bcf565ec5c0ead402fa69f108dd261188f6aaa68c502dd5455ab55269f218a3fe673e884dac278e5fdbd19ec8f6969f232d0ff89d60b0562b906899439b1e202b99fb6bb72b9b550169a4910a99e60b34ef046a1e30a646a5549410919c4a4c870a3935d6b9cad39b08767c4be76f3f81153a1515cd23a0df01db411f4c4c955fb8008221f77ccbf3385c2f5853a3d7c165603bfaff83c74d9292ba2730ced9a168a91f6d6ffd73b617cff2766dd11fd571b85d1e5a6a9a8f3fc97fe64b62caa89f642fc7917d07b7683db7ef32a9eac505343823f6fae70253e5bc58aa2073c05496c80708b1daa5bbe9a7558c7ad75bfe4029b77f2295bfa5c46df52d7a7860ecebec5b88167f667ca316cc6f6dc543b64ef8d1fd5ca0af1b7e8cd3e7c809b734dfadec79c098d3d6922dfe82e13473e9c94d62fef10d9726167dcb3ff68898697b8838938f8d66e0aa3b91b6dadf4d30fd08104e65cc3a01f55fd53e6ae8bacc0f5a894050ea9c6aa67d5da803d414f08cd93a490355d3a82f09b08aa3f6f24241885a002a407c29f599ad6301f2a131a3d0f8606e315b081f081c8cc3d5dd94d02ec3a902a797389d7f08d796c42ed6d24344246e97b438e8819d713858b6d6117c320c5664325ee9e7ef77addd5adf8f522559a64760b94a3dadeb204c1f8988d295e846d5226510b1cba5b094cb40e8798cbae7a9927f8e1d603f4fe33002a55e5c46ad6be8c7017e7ad97812c8549ce670860dfb6f6e1d82532e8a10d2ea3e26a35f5ea99ccb9dc7d11b34741cce4f2789955f69c9d6d630a9c9f2772909b9b14445123fc9218a776768707447eb1245a4251623cbdbaee80aceecc89f4a9cbb3ef93fa7975e5ab76c1de7af93a73a0f5262b882b07d11faac53048d1e4bc7c0cca0fc1c16be7fcf93bb9a193257c3e74f74b0e01e0e1297f74aebd7de8edb8c66f93746f605d801c65b8bb3f899aa6b6ed8d156c7bc67a9ce9e63bcfa6d46658b3bd3945e51c302341aaf004cb6bf4ef439fe7db6264c2d0c4b2b55b780724e7ada350f87a841ef01338be472923538f09f56d704668baac5e4b2bbb6d63227bc5a616b81efe6e1c9f7200f8641905319100ed673643000bdc469248c7499a4dc7197a0ba346a2acb8ea4f1d69adeef9099160fce15e0af338a1d4d7a423440d60e2d3ba7a0f272c4727a08f33995b4fec0fe7fb918fe7bf8cea8f37b5de727ea44296469e8e5048c2cef04b2c1afd8710df7b9f88ee8f9e6a8696cc445e3711b93043ac7e9c4441345a87bdc9d90ccfdc7f76a3796df4f939e2307e4b9ea1ef120ffa18bc7685a40e70ac90c288b8d437c82688e1a20bd29102fb8b8aed880899ca50e808b21a9c37d333938e308447b6819847e662790eed3c94065a91d06456a99edbfabe2c4a83961b4cf5d7befd412ddef9631e074f11d037ab2c41f99b886383e349da76556ac025a4cb02b36b8307549a52f2ab9ab8f7cab939a59954a945260f061314ee224fa7e311a1aafe80c27f7aa2d40209cf5831b4941d3d54ac64e08cc5d0cea8e757b602451da26738975d7a37abf33326db9f883db0b82f941a085bfb35823d70605351a8fc6766663b28593e96a53034b6e4f717aac59b946b408dd1b04ecc967b00c57192f2d340510ca7bab24a06a79f2ff54c1ebcc6870d1dbaff2c0b20ac6ba576ba9289fd9b507e64a0b02c18498cb9b9ea72bc77bc055439bd7a38b51ab2f9db72c461b8fcd98e56983873a11390296704b647a0bba65eee336bb5bb72cff6c540e6812f736dd2ae7a75bc91a0611745ddcf6fc0bc358692ae5c1a5726bb7e239a4d5eefeb4c0d9259fa6e8dc5bc5a0625661e54e98210f2cd7d125082d5b1f56f8bc19705d1358bd121b10d2a18f6395b873e469ab5dd6a81f0995144aa073532b91f00c66b58a52b1c3559217ce8bc6d5069a36c06c402b8c78f65833aa23fc88a1163c6aa1c78032316d72f7b4df18ad1ec39daeb5a4d9a570f9ef1f0737572915a197ea1c087a0b1eefea4572aaa16051b7772e74a52fd3cfb4c444d2b4f412f735f119d288a4032f7472085ed4d9298d0d1817a506c593b0acaf7c359b8f8e6af8412c07bfe0d3ed7d6cab1efb74891d233b824f3aa18450d4a4e4e6267a2058af103cc7fc392ddbbaa87236037afba49072795e2738c7c90344c915bc6bce43931ca7fa6811a0d6827050b713947efc6903e4cb49dc2aeb47e13bea7b536b1dd4406e359f0551356877b794c8c9e2ef9af11f67ca700b4e480a1948881d0f499186b9062ec85baac3270bf0a42f6af8c8362c0d3b04af2a2c2eb39e9abea730be405f750361382f97b807362d4b8c94657c6c2668d34f1f95eb71cb7e143ec22f9e2d1761fe5b6f17c2d08635d3ad98e52b86ebff7259373f7a589c23f634203420987fe482e7cf96877f789d759aabc3457cba0a982a533b4e24df59309ebeafa6aef09926c4cc73a00f3cafe6bc1715e0144e8d418023661c9bee83f7ce19f1056e396a88290586b86b7d77eaf2ff174b48dd5ba5c0a8fd71be9b553ec398737b73e4e70dc67e110822488de151454a4bb2cdcfd504ccc4262bb4e8dccd765212d555299dbaf31cce730cc434b32ca0539898217dfc12ed0bac5b63da83437cf872c6408c349ada9cdaa78cfab6e9944ccdb8a4feed616783be1c1c2ac9daa36af0b0fbf4bd710a5932a38e44cf15c2aea37f7d77f49cb192d3315dba2c3aa6396d86121378c009010dbac09698d166a0e787a38fd44a43de2f072a6bf7a68d22c77aaca0f61600f77d52d96b4bf056f6f98d66d544611138fbd00ad6454149fcba0a173f6eddbd122ce67883ab237fa6ce3a2a7bf49966b07ab2383a41e54b3c5e184b4a64431822073f1ab5b9dc4f15ba48159c9282cc2029d72fafed713f4e428e7c43a6ca96179803b4c1572e33acb298565b3b9c20545a08df9b1744ebf3ca0e96d83d8a59960f224f34d9311ba9c804dd6ba7f70abe77661229a668642c6e5d799ba69aa92359bd9d84854caa6b11cccaa48c021e1ffecbe5075c83b105db619c79c58f50f9c444b93e6019907c9391388c015fd8ad9c7f0e6bc3d3a258f747b44318630f642d554615083a1cb99d799cbf5144ec61292632dcd6471ceca2d60aea14a4074cdeaea1d9d78886b78acd369b8e04a7d8460265c3c57504c54e9d4116cb68b46019ec84c56deb9e1349abafc5cd142d34f8158a40dfefed1736110bc9387f763ce9258d1a3395fecf24e131eb5efcb8e10a5651cac068d7b879e416b3eabfa10227fc962ff6348a8aa368c7c147fb299309bbfa1fe85e44a44189263ee8fe5bf12bdd2eb683c4ff1afa74b7692afa89d6b183b82ade7a9b8f7df1e4eb7d039a62af7099154cb03603cb2202f44897adf1817e59694ddf091d78b6e5ed5a3744c76c9e07ce9a8d6e38faf7a736e1f97a9dbb08af041b4ebe096446bb8169a54b1cf0e1ef14120e68ea77d08f2d340ec39c49d2b67a91274f2429598b1cedd85a9964e200591871bf6681b7f06b2f5dad3e1547ec1d6820f6838ce16d7ef173860db40c1118ac9ff28512b591da570f3887345fd02660d5921e077b4e07b018e83a8763797f5e26a45182dbbf593bc37cd65b58dfe6808e11d65136ebf38b34b3242f5ec6eeb17f0c46e942e2e2d579904f71d5f9b772e2e45e2b4bcc7acf5a0c2b6236359b6fe96b8eb53da7d01b88d764e7e36355db556b7e4f6843ebd66b843c0b264a5d79fc16186470c36b2a3fca3bc5490dc3f7310adb176918fe71794674bc92f9bdb9f531dc17302daa9a5fbc48eaeaa5b7b3f12595e71890898a2796d3c9a4dd2dc61daaa42c6a50666f5d2ee86aff7fdae6a8a560b1a27777f3bd1c071adfdf7e15bce58e432e9038dbedbaccc2680e7d58007c33d70b9b03ce4e85f0906d3d762afc8c2fce84cc57f42c65c8398183e3a90b6404f9c608664d981671a0d67cf642646029383fbc104ac2a368d0b8934f71fc3a588b9558a1871015491c01b93969400fc6de1cc2d03dc4d2914705c4101d72a8c5990f9c45b8ac6f0779f8ad9e4698558e684feaaa129c9368f411086b0f73a3411aa550e4798aa945192d98e9cd956edcc6fa49022a8ac1a8ad8ac2c330e4d1f3aaf20dfd7dbb7eb6a13d738d8cd4f33b96648247a3bec4816ce0b9454bf37abc4375256e893ce864a3765e769ef6422f6743cca34632b564361077287163a78e77a0683ae2ae868f3eabacb8b8dccb40bce7b19f6a8a23dd448c7bc2dc2b14217ae4f130c568ae8a0c79eccb914e1ca7ccb209669dc665df9d6977e3ddfbbce85fbacb623c47c56f5f82f110b7dd974d0c29e2dc62f23924bbf6dd3b39041e25ac38a5247c4871527ebfca9f0ff06593d120f10e598054478cbb7257f8bd761fd546398ce1382cf0c9bbb9b2ac72d52f78e273d2e09a4c17417f8798b71148bd5b1232e312866021bb5604b3c7c95b52f965d3ba97cdf5ace5e324f54da6021d99aebac5040802c522dc98b9b8fe6a60c8c9b0da4041872653cdf625afd63e25e1c0ecd0f837cdc89158f6ec9dd5c08746aea5297821dd76d4bf67a4e5934ddfaf144441875cfbd2c6309ee0fb1926d7d64679543ff573c8f2ffb4c7bc53998a034e814df4253f08a23e3f0fc61ca65483e14e04e75da5812998c5c407632132ccaa7b79a4812e049d4ee76dbc00ec48ed1995ca7dfc59867e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4cfbca500a5db326bd70abdaa729ef729215d54f185600a4c305b9bcb39b245345ffe3ee51e9f09105b7a764eb9438523adfcce461e259c83a304fdb16d01117792f59bb1e2d09cf5c6541fbd8de58f7300056b8c4dca868c82374dba2ddc93bca16559f5b6f584ab50aedb2caa818423665b642a70fd9b6ac14be723d998399a81a7c8459e3f6d9aee41e5b669fddab59cea894beb3a3acee8144583855b2017796f02a7aa8217810361cd06965b5eeefe9a9fab171fe51b16a263b26ad0815939965cc0938e6b78df44a41eabb5bdb6917d3ab0dae65ea0d69b528abf3327be739945bf9bb7a3ebab04347cd28262fc17e10d6fdce46385ddaa8c94714f71c316d7cb1a7c27798d439f26e54a08328bf4855c9f6253d1d0bed2e5f93dab837053ba6d972188f367ec9bc78642e9edf3af61bf7a86b2353bcdb5cc3abf7c0ebef97a817846e17ee8b644a09eec9d8f8cbfcc4013013d2b927f99f4c41664ca970f48dc6716f1e98d7139f42a5bc85b572d615a1ee682f644725bce22c9a956fa814aeffafcc626e437a97de471832f5ea98777292dc180850ef80be318576defaa6bc3b38965ce8f5f277ad1ebd3512679e24e227fe790576e8d04d558d6c9dae28ca959609152a6213c0b49ddf7a7ef9e87c4d430e1821ec13f7ff79e9e2c31d20e87e88aef88a7e34a9293f3d2362043fdcef8c6f7eeb2d14dde5441419a2739361d908d5158342b02822cab968acc3c9709ea3c57ff4bfc58403c7a5f8900354f20864e23094c5a95c5f3fbad6ca565d045198ed843c71f69d62009d6bc53894fe756b3a0f648143069c682545db441c6632101a434cd0a0e047be2e283a92d7f853650e97eb37c746a3080d6c22ac5b8f85a3130e8dd70fed78312802f7dc0fdca9b83ca38f27cc8551cd876f37e56df5b8a85832c8571a8012910f1ee339a94b38a5b0ea11aad801a7f81ef8c7ac9ea9614ce7f52e989e2c28dbcb13308a217ace78be36817898b69b0312addb20741d889fda342b7d648d1afabb8fcce1c173c067b82e46311f5397f351687b3d0f0d921a7c9ce22aebdade23434ed88899b818a59a770fae14d673e05f21fc2619cce908c345aa8c4e5eb61d678ece60223bee0204ef456043b47d6bd1f51590501caa21efc54e967997429ba2cae1897393ad8789f0d15b97d486c113e9e7efa6357798f3f0596ba92813690b5df967624e655e16af92e12ee916220a4412938810803301de213dd5082f3fabdceee8ee55fdbafee3b567df77092c0cdda6681c29992f9ce4b2a759b1127875e2a58faa1c01579bb94648be38074a107bb91a5fa7851e22c2ad997a61e0237df9dfc03d960f69b8d66d545bdac8f2626011b1c2b19c060f323d3688997c3f1dad5705a35f11e0ddc27adfa7a9cf3878416c147c45e57ef00764a56a965d2872eb66ac36006d425046f371d1c61d971a61b6f60553d67f5f9e5808233e3eb636d2c880d07b4f591aa50526d3ce54e6fa6b70babbccde5975ce8250deabd13349f915eb4bf3bada5c7986c1e6910843935dad8780bd5472a9f7a8d0161bffd4c5266c7515a6a3134e9622da1c2d32bf11c908532427809fc7499a8980372fc5005387b77bc19f9ae7cb70b8f5a90870216aba51199dc336ea0712f7896cde89371f52c6fb0549ae56e79644874e22175a5d3824c6b7e228ba50d13f48ddc5b484b9bf012d4e7fb10f3fcc02ba6e0a3a6a85d111cc368021a2a138a27d23b797f50d60a5de22bfba70828d3a65b939c4fad8f326f7e4006b6e34a75d73c38e1c5b4127438945fc499b2b4965ae2b3e71831ad442dd004272f2cd39f2dccb792aa4829b6666f6a65f5aa38b594c8f85a4d5b27055577b3143612d0dfe622364b4c04c12c218923147d097ecb5e6e38a57b7764d9c5d01d8c73d72a8a9370e45b2207c89755024a10017aa1473a3869b9dffeae793b8e7cd18eb7e2ca968bd9a89dbba2b9cf3649274bdc98dd0e6ab59a567e320fcca0d7dbada8c4c48edaf2a201bef06b13ffa434cec503edaa108c5afa06cfe0ee83a524b8a2f021239114c7a90059df2c134ab5d5f7e44f2e795ba65fb7f2c8295093593112cc140c3d08c62f4bae44d869eb9de4b21134053eed8cc70e4617ccf8aa39d07b64d3dffd02169e06b355250bbd44b1d68b2374f02db9f79c84179fe6a69bc0c8ea1be8245352adb00e5608a6f69915600cb6f36d8c4fd9e4af575f5d8e1f3621349de57cad4d977f133814fbe802f022c8f8a47792f1f8df97ea3d8a3ed181a8569ff88af6fe2e1af2547a4b852dfa2ef0b148a5384e2bcb67cce7bc3e80b04feeef159eba518454d784255ba803ab2595db86d85aa9117f5d0127e1741fbf4082d90ff7f5998cbb43f94170f453410ae9c9728762b8e15016e60e1e80c38aed2b6f3cf34c9f7efea9966f082b40b43d08107ad398a1969777556a654ad0ed2aff7519fef3d18f61f562495c29e84347565739471d0deb513d984751547b4098dc5f4d1489edf951e3910fe445f6a80a65e63c752d376598e097717803da1a16c5288487e822c003c44f4b780fd4d0691136ad08429d00baa1a4823d922680f7cb36e0a6b7007c2326f5900838fe4b6451a3c0cab13f8f3d7941c3a26b8bafb6da376315148c25d133a8e13ea63de8d5a017ca6ae89d8f0d99257e15c08b6a7498ef13a2c150e9204b6d38e1600743005578d3665203ff6de955c21b25ad4b5e436a1cccf85357ae0cbfb2d0f459377f08b6419ab4e5bc9dd190b73729b54a2c3343418a0e0da4f6fe4e4eeed6680e270582ff37aefbe78c5d7b22007141ed0c6b58a64b663d82cf7d67e31db2af7120df039bffaba5fb587981cb30cba5d8662a556a3ba9f193c0bbce0452b23f413c4576a4f4d6116232294e0095938591bb1c5eeae335ab919efbc5e5920109ef1aadbe22d4c151c2ca73026028170f2efb01e8aa50b1dabd29b4fb9d4c94ab812541dcfd9c0ebd822aa337de9fbba0e76e5471aafea78027459626f21a17e2e99309dea26aa7d00901df5d66e67866742fcdff6037413fab503bc35a95867d6b33c9afd6d7609243f7bdc4ef08e0797b311b72f670b4ddcf64f1e078c48a1edf92e6e03846c87af3f717ed108d48867fe9f64ba9bf26c54a9b482a25b42ac384564b083f3a0e9bc5a8ba284aae2ee19b8f1c6e148a7a42cb4f59b129519fc86c06e416feeb6539818de5057321399318d83bf350fea092d4035a4d4f7357c0b1a31839685dcce8eb79d1abab6e1560a8a781c7ffc5bfa12042df942568570fafebe0bce85f17457556c707477d4092eba742a1da3cf8281f236d8e451820d5b241cadf1560f51345764233256dec38417b54d7ff6100d512d2e7acf4b99c82d54c64026c8ac5f07ad8af029ef1f50d8d01145d0e0240c5d27d875452286839a5359bc8d8df86c574f68a3aea80d0201672ac0a464d850768f8344b1ab2c1b5a2eed4202d00380be9e27c2209aedf0f086af02141582f0c1c30774a4fae5732c7a8fb83ee8cb425b311d3b9e960f11af635a71fb4101f9c464cdd3b9f4dc8fb846c04981b340ec6a51cc212e6c176901054a68f89b715dcf16fc370a74ee5f3cfc9d874dc3fd4c8747f9818ef98f732097eb19a7291f0cc6a00978d8fcc168035efb1564f83af38519d69661b33fc7f899a8874bd62d58af52fcb1b43ca1717078fed76457d3e036b22c692cfa3d5ac1ad929c67cb7d09d0caa8a254c66fe73a32ef1a02519225b801c11cca4386497838e46fcc9e5a2b6f92e022639c217d7a52437a7d27ea444c3795eaa71613183ae844bc459c2582f62b112ba2965f978daea46ba05e02432f15a6cb2b864967b2df99489cbe0cf7aed07f04fed89afe28583a95cface68061ea96f31cadeffee922bb15c2e9753e517b132d44bdcbfa73a03c10890aca457e52af2fbcf33bd53c21d6ef3c6ad76d98c14d5102520a989b9d25e7904b96d6cc956c62dc0f6c6807a057ae59679078fb899f1c0afcc5d19cf1d4c8e855a116147959c61875064f21792056101144bd17214bd54d89aaa1d363fbc1f7e68e91cf3f5a03119240f6d206adb0902f0b5822d30b886e2a4bd87ef592a6aa0ab700f77a26111db609e44f198c8abb98aaef7fe12107432edf05b168aae7b5305ecf0e3576f2391effe81562228cdfee306f4f779f92c53e80ca8d5e6fa157178a1f17b7d4849a62402411b761fb38336282993a6bd5656148b964c55d58615f45f0c57a749565def1f760f1bad2a6dab48de6e47abde4445999adc6dbdb3701768df1a33104de757ba5766fc502c4c2b6e18cc90d36c12472bcaa5c3e05426027d6f56e9c90fa2b39ae55997aba05b0698595674a7c2c6966f8c838bfa1b8bcd443d1ca265c054b9a40d11bbbdaa3b97916c8dfe8cf76a77c8513e45e78f01b7112f969033a1550cb7e1b004dc649dfc8a4ddf9f5ed0fa90cba717095dd71326a4e629abaf6e7d76befe70c23c21bd7e19f0c447635389a1bde26768cb8a642c0b402c06f3281df363a0d2b55193f0700494a3d7b493bcd5b4ffc89035dae1d75be0cd828c783994b2521c075c8161284e51265dbdceee9f0462624ded6ebdcb66c6c05b4d6fa755c3aa0252d73866a84e419e28de3bc8ee042c64d43e11560f27ca4f04d16d111422d92c8ec292df0a83ec38c08cdfc3acf73a959b50525b4351edc3469668371a273daceea917d40c04ccea5fe28d14fe5c976d70792196f2dbd62309971f02f1888f59beaaf812c5395c470733cc967022fccdca6bfa8aeecd3c572e269a7868deb261bcd38e01d3edf97f1159b7e1a5a13269d6b05fdaa477524f725a6dd0a7c96cb644c4a2fe6b15833843bb16d469228d2300d19593affd4148bb8a0c0951d166980f38b34261be820f25b8178c5404b2ea17eaacc1c2455fbd459a42152c7a3a06a5db10d7fde71394a91516db42f95c17d37292a28ac14625abe01f205dd8316d9b5f7459602fecd84e1d3ad24ce5297befe96910a9101b21bd9889d70bc58e9e804655921cf614996f5277ca7bc203aebdd49013d8029ed770b1dd754ca9d17e593f7189d41b6d21513316fdea92a49903f07fe1db4e343adb40da1fc0bcdfe1fff3e09cdba0a242d46307cac16dea6bedac367b826e9378e669c4fbb20208dcc2357f8a4acaae8e7db209789bc179d344193ad90935134c718f2f20ee4912bdb506bf8eb912f6ed1342bec771e02b0202566a4b27e1c8beb9f704554d418e69da99286bcdb6e3404b8b242b28726ac67c6d5cf9d295bea6e5051e4c95dc3eb32029621baf529ebc43cea67f3c055e2303e90936b6b89d864353471d80d6ad83529b158258e20c899d3bbafc5f2cc834bb45b13a1e364cbe565e0f949999f7b4148f8a695584a9f42a8d64efc40862b12a3727d99b54bbc1f66f5341a8b7adc0299732382b9207b03be0707987a7db9862ebe14d28290ea1792aac3ca135ccef618a4399efe825421763a438aff50d3e325c592d8235d2c0e8eec24159fa959d24cbfd33f4df7488a07e29c10c1b4e11db18623e88c9098fb53b5f6c82a53607c85535760fca2eb773215a1f39f77304abd84d68f27f495174095f3fc80d2da1167c5466cae721c272a9c20e1c6fe0ccb8948d35e1056b77b53953e9c41296adc4bc9ea5e4f81bd2fbbaa70f2fc866ce4411b2c2ce4a711f4c38cbf5a5ce25f156d7d1e7395c02da5bca76795d375267e834a03f5073334f6131ee7ba45c4745feecaa33cbd62025e69cc;
        #1
        $finish();
    end
endmodule
