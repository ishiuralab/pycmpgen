module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8024a0ab7bf8f61ec80952cb766b88717a1825b8ece3879ea934142aa9496a7026fb2a274c6d89a1f24b1db66ae2a1d7f2c49f7e25dc683cbc5ed93dd10f0687a9201f6f0aa74e32451d26686c11288dbd3102cce0c4cb02619c57ba40815674ad77bf2b633d009087fb0b979251b3102a0aef855b645220970d9fcfd59dc73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0569667654859ce4e4f0a595bf3da6ca7886273263aaf58f7ab2016f3137c73f0a97cf624133729446d8dee2b8bfbefef1c8857707f1d8717db38f4c9cabf98c7e052f31adba90ee8abbf852eb6b2962999b8de8578f73f001d0e9a71d25c94e36fb87e5d7c8e967ac5072909af93fa9f3b9bb7312a44b2f2973942d2d24b73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habb663e15ae48f4db98df3a5a25301ab838e660ea10478f309e726ee78634d0c5c39eaff5af69974d28933ca69e4289ccfdffee579360ff53fd561ba67b92d1a3782f54d0641f337cc65acec0ade7d7cd50f631d177903a5904478bf77d2d35f173214b0dee4017ebff5ca49208eab83df7c223e98422428a295afa9cb577333;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8882d3b98e0ac1da0f536ebfe7634ce79b3cd5e3985a46d5785a191812d6a215b0cf2891d16750f78830c7f15c6f24f251530b99749d1ab12a6603a38f3ff18c48a448159077596fcbe7bcb71ac737a31b81eecb61f7ed7a63656d359314189ab07b8f5d23615bb814a8b1bab0bade7b3abe0d311640e3c41a2e50427352a653;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4e1ef7b85c08cb00777d8a005dff7b3347ef517aa6ec6453e3cf4bba44dc30d7c41f0801d8ed7318d35501f435b01f3f024f0dc7e1dcabaa6b2754292853756b2d1723270e2fed8e8a041b27d96b7034c310e3db746974434658483a5c6053fecfdc7bb3d97639bc572b52d4a832382a6cc955608c6dae51d5f5003865a97c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3dbbb9961ab22bfd2a0f825c091c88ca0b59998c7aabe687454ff19ab96f1d5b8818451b52c46dabdd1588ef5367b63217094df627e665e3363603ede7dc3ddebc68fe618f6c4a0ce76c3943628d1cbac7a484cb27b6340e4dec5abfbc1f0bb1f2d4a3aa9dda5891fadb9a8643273c94b33987c3fbf3ba3d199bbaf3b139f7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9ad2715e9b5c73ef5c771de9128e999232dbb699da0bf6d27feb053da81047c93521de88ddb90f3873ecbc84761a166dde707184e862d03efffda4262274a426c5e7a90e970c7156ce5d7d7eb04ed10b09e3066a92c807dda755d09bbaf7f9ca8a3b60c77181d33ff9d3db6bc1f37508756a93aae8c240f6093a36842176238;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h710097f08f8c8064b81576fd3ba440c993d7a0efec4e8eb31701d316de9d8c0bcf79a3b8579bd6a34a258dfdd4916ce620dcfb78b2bee49dd840ecb0802005f89a4ed38372621498d0c3eee47f5639362125f3b4fc1bad83cac2461aaabe1a349f063d2d049add926f36ebe6628db5db7447db6825b3cb4e2fcba8d5648dea1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b6a3f7ca41ba5b6a677838b20183390a6ecc6cdac555fe156318c1aa75beb14144c6d7cd7184498d9d382d5c0ead51424a1d22dd5da61fcc86e8be56b9a2af42ed90af2897e6712bb5cab6d0924d2642196f6531df6187d5076f31b41fd4257ff82b213b12577a518df00e5afbd5e1a8b3430d08ad6e138ff880a15c9bbdaf1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h550dbcc8d8dca375edd1db1c0a44eedb5bfd8fc022df0a49719e183b43e4fc645e3e3a97da143b6f785024c0556b8f97cf779dc8d67bc26ba904333469e0fcf290a9d90f58ca7ce5284ca5bfc66696f5aca74d138e784191b73ab887c620162ed6a953ba60dbc5e2bc1ee0aafd9193176a8e6bedd6f02bb6a0b717c15a5068e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0838989c74f40a9ffb71b823a8935ecd9cdf47a2c0dadca4c5f62c37b4c47f29fb21737511912441063213063e10ecfc497e164890957512414454b826235d556d10e7a2e3d27716a671e383680c36c50f6b0686b0e7c56555f449407f31742d662ee703087cdd461743bb048ff3ad4d5a733de4326d0d90df5ced391d60585;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37dcea7cdbc9743646b4f4365b2047b2d64d7e4b7cff321af84b06eecc4a46d341e31b464827311a48c3f43424333c5cb4219450e731aa2cb26885d62a469f8d54a402e47e31aefd3b0aee09979b80d1888f4f597bb1781a5954c953582f1d7ea60cde220c68af0a756e10037b1a81dde008a7f43aabaed4e8dbdd2b69474390;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeb33b52e261acb253406bfd6476976f52602f41910a7244d849b2d7f03aeabeca92d8f4b9357647042dcb04247bfeb63153b259c7bd4339b45be09997a8b4c64027b6714499686e1bf9b99e152468a92dfa7113713b6e7ba0cf674ce80152365676c63adb3152fd31ab3d1817d7bf69e6df5552b2c9f0757f5f98b51af41c5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b9cbef2334a8fd100b823af8972031db78134679ca37eedab196de6c6cedce6112271f0d734215cf0a08eac1effeb1798eec799da9848c476c44f93886790f0db07d16330f604d86088e748380ba3cdf8e07bd4d19facdd3629a62a97f699837205fca2d29d82739768d0b94f67d44cf218de31e474dd98c25bd9bf3b7bc654;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57c7eaa15e38e9db9c711fa6224416d83b946cccf084195629cb252248c2b1cee5dba4ea6dd77a220fa793319b9e3d9eb5056f5a806e0e49beaa6472e7fa16b98becb7cc97fd5e518e7e59e4b3a12af57fa2f4094eb7ed32e8fab4df0c0ce369b06f0a82b09d873fb6277164bf767c1d888f16379ad8ca8134d70719b8a5a484;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74f702714189358db8599392011e01370ecac0905ed1ab0b26057c68a6bba1b08f3d02cf7abea4271aa3d5acad49031192950b706bb151ae00185f9f65abc0fe07c4f478d40f97ff294b8e3517b8166a47e087c349587dc84fa3038553d4953294c7f01131cfcfa2548d63c9b7da7292b0d0c61adf13bedefe5dbfe5ca578639;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23c93655ecd852f0c07adee3376c4d4d1c346741142ef7d74b0f8cf509376445130a4aef7a5f5f5c811d26abc3e6eeddbd0a77f12eee4f7821ca543c3bba9be4a05f7a3fc53d2193e14a1b3e690d401154820d232eddfaddf61053cdd5946af4545bc86cd28d7feeb841e2bfb7441cd02747c7394fca87d50452b683871826ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95bd3c97ff7e72c82e38a5e5b82087fa960a944f0fc590f15394a7187c25c41192192ec5851c4a52964b6910969b7c25d26045dab8cf7f09c10ac5355fd5273c28e9e3ff2ba6c95bf579ff65c6d438edc7033da358451af4aff9d9b77ad76d82b5f21d67bb1b7e7e8ea09adddc4d97e0e43ded5a5557e0db0684715ea798b186;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfffd005b1f58833438a0af24ae2c9106cf1e7e8d5ba302e551adfc5acd3f554dce9d7bb5b58b8f6f378c8bf841af6274d421702a710e103bd559a2d7a885df061476cbc4fb631a4f45ddae99d8fb05f0181697d939c32638b5847947dd85a5634b095ef132cebdacd7af5c40d475a12a8cffcad6052c7ea5f7b4d6e94d95a71f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7de2d2afb13b656dc17cfc7669b863310c81722bed144daebe4d8f67a6576ff5fe62e7a528b576b240a251a733619b5cbc1b0e806831f2ef6ad7cfe80404b16c8a65e9632a701835080d2805a79724009d4f0d6f8ae1b7c08e896e182aabe9c42590093ddfcd6ded96d96f2f9d3a3fef3140631e3c720b88957d166b88751d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23789958c9aa188b4acfe62b02340e04df7d972dd4e8dd4aa9f8fd2585a83df0b47ca0e39a4394b4894b6d18a1e95abb2a9412b06d3fc516766312ed1d7b640a73e25906cb83950dd2ec9130510177e16f5b3354ded86dacc0381f1006032067c69e1da6c18040defde6b4c506632c1b126a210893930b3d335e6953e14e9f5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf912c8ae0d58d652fd0bbe3cdc707c68b3e974df029a7cc5e9adeabe3fb0bf70f8cc4eba8fc373d446166f9259165cc4cc2c35e56bd8f2621f6544863536f215951c592cf890641e74c40aa825754272936de430ebc752bcf97da33d55974a5b7cc57438207732f2c231efad7edbca5e1cd6f7938ecdceb1e2ac1c213dd82330;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33c7d85536bf1561c6601cf090d451a77121cc38a43d49be1403749c242e7e7bc9b71234a5c0fe30f7b29a24fc5ebf1dea901f60d31c8707e2ef6eef472a13b66987326f38c6a5c6036fab0eecb437782bbaff1a9f6c07ef90ffb46a9b6ddc00c4a195f98bf83970bfdad646f73d5b94f659c6750fd7c66d8efa1907b69fe690;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a3dc5aa22d6d89d08157316a63a142d73a02808b3520ff40274dd5b8eca20bea28f7c0b7e958df5dc8f9940333352356685116f7183ec4870c8cd6a4bd49d5531d8563aeab1634c88ecde8861cfd169ffc421913978139c68281243116f6a4c02575dd63e67c2199f1b66393d8cd4d88857947508a2ce23648f3e5836919e02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cdd29abb6bfb8a1e082d430c866af6eed4879654d2f9baf70c25b66de0f47daaf22da9e1230fd1a8ffc45b1782dda7fd4b11b235880e40c159acd91991ec05fcf74e3c9e10c6c6b7ed17647fb1736bc41af4c387af2dd6cb8d4181f3cf36f89c229e9bf94e57071fff5a8cceb0e7ed9827a36729db5e805f1a12a4f57870b7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc3a534dc6059c9d5939c294e7b3f7e79a696e8ae10f34e4bc4491f877ad3d99cfdfba960857467562535fb07e6b580f47bd3d20b81e5e20d28ce9d67eed85a1dcb49561d7a17aece889d213181eebe4c895cfa65bcc704f2bb24684400aa9e94f40c3c42d9b2b13ded8d9abeb2837a8cbeb1434e9748a6c7e814d3dbc1ed2d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30f09b5be781ec5ac5c85d12354b1c45286d51108c8c75c1bf2938a959dd693c3e6f58f15436517fb317a118f4614de60b56549a5d87fcc518edbeaa453b896e4234d09de6e237f521a2561d296c7ab6629e595a4a8de1f4ccd6a124b9a417d70ea2fb4dc7c58d00e658d75d1dda0160b7f19e086041132cae9d826741f6b5c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5ee7418eac4c14e5a44e45b18865741391f5fe58cf71d185fd3a4cc6d0c7e57fc11f50b014265314e6022c5a24aed573dd2cf5a63e9d7b4d9745af003ca2b8e284d47bdeb9811373d7661599a28739f937e15a46a743d9dcb27478bdb24a6b46e135b2b8efe67e31e38cfd5978a2090ad58b8fe1414e89353aa3e79d7949855;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d868a9305b7dd91945318df2b06c727fb45fde394ca154672fbe341c5d58a2f498f4031f1fa59827a1cc40ea44ab613ac7f5183d3901f8ccbcf87d512fb9302d097067ceed8cc617606b7a6214b138101f8e56ad1244d84c7f6f6c00ff4e3ff2c01c6da88e7c58bc44923a80843e286af66a10065637cf6eed7b31e2d22a01d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c36c9524aae5ac5849a07f44f5a07baac5ccfa734a5fbea97b60a0cd1aa7401788f1f8f49de6b163c252386ed2afa20c862ab64a7f4a8bcc66886ad31a77f90805271110959951a89dfac0f86a058c02e770a16be90a7e576fad45a03674acfb2683e8d067d65d6090cec22418308e1b5deb1ac13ae0f76eecf41db186b7605;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31d02f1f04dbb3a9b8a4f0668b865ba39702a7123a31ffa981d403ba272c2b9ea4666d748298d4a588da5d3b7cdf829bdd08941c8c26acb7127fadf8ab6fefea331fe9751b826c556568c85e6cd5703bc3a2b21af93dad33271fe1487a330c4f4a97523260ac244f8f4cb212e9f6282f0eea07ef7eee3def5a3d986d4309a69b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d94fed8ad6fde53f61912eee46b04cd1f2ed5a2aefb421f138a30293d6e41e52c323f070974bef0331d3912cbae1c7e64f71c720794b93110a131508df2da088246efea32e1d7c426085541ab9c47c244601f6772aa3f8dae2ef335b05a97c86218eaa29e75f578bdf8dc273513aac4397fc8adddc983492039e78bcd442793;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3621c318baef158cef2dc8bb02b25735470a88c0bb51feadc3bfb7dbb44d021b75d0106c3d7630750eec4ee25ef26ec9b45231781473977215a5803cb89aa911fd7ece4bbcc723ccd2f52852b3b24f8d0a4eca1176231ae7d0ef075abe255a983c3fd6b01e28aca5076d3f4c568c7c1f88446fdbbdc594b51794764c4175f4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h242b7b59a81f84a8ff55cae775c5e62bac731168d54e10132d63e30a0f5b927c7b713784cbdadd6db05294ee6c8f9a76b54446de5892092e13560d38cc4cff3b289cc38e2d451b7bc6e480c4672648d3cdd16912596b63ea66c6dff086fe46924b69895aa4c61c20c41a7f6cfdbe82092e0a656b49dba6bd384957665fcfe717;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1160525464483bfe404e582c21ba82fe63dd60f60c3e244a5d721ae678a74136daee9e38af3d25c76c84cd4983c877f2d7a7772782f8d26607183039e87d0ea6b03c72af527094e709b5116689b79788485905d15c14bef567d53cd8dc94ea04fb57fd983daaaa83832d5e1b96123b9a52947c7144d469b9a1b65f7895f5d244;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1de67bdc81656b3cbaadf0ba7d7feea0b79ad9253669f9c2e5e3ec936cb5a5aa1f28251024caa2cd1afc6244dbb6980101ac2dbf37b4969721f548ab89c08c1f932ad57a757f567b871e9b5a03770c61dd6c92cf3bde57894a0a1bdebe9fbfd1b72dc4714efe9e9d16cb06401663c6279395dc318a6366cfd29022620fb79ac7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h809164010a9ad67ed4b49fb8ab265e1463ef0cd80f3e1786da20177ee1535fc27b9a896d09f58d2dd076ddcac50b9aeba101ed7b7c6a6a6221b07d8cee7070690a6301ab904d93842ba1ece963d6e9a522b995534d8f54a9d1f5d0f7f48332fb966d20204d0f916c2d6bb293653e0e160a0f5d60a1d41c67024e1d7ba195220;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd8490bad5178ec5a0dbffe59bc92740712f645779cedeeb7264803bb65e2fdbb35f1475c6c1bef86a16614ad4432f0f6ccd3e62723fd62ca7ca160e54854947bbc07cfc349c689ffbe45959736653a0c229c3acd417bb5c07bd3b99841fe8e08d437fee90863993bea584f4d0caf2a4b3e624b6b2314325b3290e3fa77b3aea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cfac5b844d149def9e9df13c3e3081e90319c7cf601c2f626e09708f30da410d3511915dae3603eddb8267f85422506549fc28bb38e09f86de0a1fd192129d702ce83b0e61349524e70519b26d3751ee2a5f94af37744045ebf49aa12325cce229eb1c90f24e294acc2f858c76107266ce09374a1cf9cca2592213848e3b079;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fb2f2b3e7e7845206313cb8158d555299fd60d212b2451f416d90520c098230cb148ddf59f93c9b6a4c9a75e597faa095d0b893ac6dd65720e1106b6735b342a48e08ce5904adf6b95a17537480cc23b60670707e16a71359f3c320dbe8cc129f6fbf48a6aaa5b6a17e9aacfc2cb37df207ec1141ee6a3d1672c1707ba7aad5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb385e08c25e5b1bf252cf87f9191ae85e234f2232628bbcce7eab0ce564fad499eedff07e668bd99687813d21a42f5ff6fed382f257a099e7c6fef5bf7205548e32419b785f3c180a0916fe2e29eea19b71c34db4a759a76d3feaf94a85f916945b34afa00a41ace657603e5a3e678bf2bfdf3ca5c44d8d8ee945d1183622eae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he44529920b47a6a17e4ff9b445f50d81b7c44b8c3afc2b11d6c8f4ef5c6aa5a91b13d5e16aa7a483811a66c940143bdbbc37860661d76d947e0ed33246f60c011a7edb747ab17f443efe0f5736ded4d2c265206d9c65ac05bc9c8e515feda2380db4ee0f57fca4c4a36d284167be328683850c61eb08702397db8511c7649c40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e75a4c8d4a1ecceb08d4f10f2c55f1949ab35f8b22d6d64fe14d06f609a535b18aeb6f95fd7e4dd3af30eb701e34ccfcb6a66b5e21636cdb43ec6070e94eec4604346ea985719cddcb3e4983165edbe5b9ca8150e424830f108b85d7a86ac96ee2759778c2f31bd32a60d9aca15c9fbd11ad811918341d1db4e6cb9d66cacc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fe59c6056873603fd5d2c1327fba13432b4828b33825fd417a887d3d87fa7d491871c2b51b97cf1b3af52f297781d581ce7ea5447d0747ff9d09ad1202f6cfef7469e7a079abeb18be8c5c9be3d6e04cd05499f5a6633935b3f7136619c08c0491e6717a76687d8e47c347a79cc1ce71ca7c6ce60d387a1688223b4a1c2ccf4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5c1d026ba1045737147d1365eb0cd16e84576dcda50a7e547c0e2eec8f933385b58aa26b1032f1a1e49de96d8dac48edf1d48df669592e02dfcf3596058529c11a28f2f1c39564d6c2757c83e52f73804c99843b2186324450c6635c85913a723eb8ce325fd0094d98a4bc91b32127d50eb7d0c96c44b83a050f2a201051eb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57b84dcce33ab1d01bc459db95a96596176a445f3170f92ea223dd0f0990d1a6fad900761cf600318e3e6fd594274f7151c0d2c20f962d7db81da25badab719d9cb82ee8fb9ad98fbc67d2be4f28cba0252876908f235f9a702a3fa31de03e792c3ee936e7032d6f004eea10f8fc2211ec2326e93d183d055e03900924829380;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6230bce9a40f606d0ef319cf12e100b8f6390c7a7ac662b1a30f2fad7482f9275d4410e224722c188c1ae4231e8ef7a2ec5e07794fb09eb7ab50579854973c4fe8a997e5b99dc50d3363e0b6999d89d0d55b983cc866df748efb3a730e7422b0b4d9d5a2d0111e9ad482c952870598c809e5ff23833d46e80ac5f6050a04a74c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f715333ebe16c7418aa09008573416f4f9490c6c0bf73ea2fe043e17ee73f27339a8d0f7a270c0029c3f3bfb4f1da252538d4e97171f7e8be0a15de367f67864ca3d8b92240c35374265c4d6dd78acac46d349594c4c63d816a2b867093b88ac66f208bb94bb38ac101bc6e93d313d3ae96b2c0250d1bfb945a7ff704844ea1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61289b515389cae47c66b513d97abd7ea14fc0286e09cdb5a1618f5fb1281aa975da3dfc7633c8b18437618bb7c0e999b692f0ccaa41be6e362e6de11cbb881058678fe9a5cf9aeee039779fe8de1247f1c44a7912c4de672efd1cae50f862275ba43f8bd3a58827fc0a1d861c1a4ecd0932d0c31b486d60a5e7f43ca3927a9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b2c845148096d11fde70ba59e566383b8900f0a411bccbcfe2968e57813e0772b2bc6e7534320106943f39712a7ac4004205c561643f8fffb0156612c6d9210bef2b0e00a79955623e341c8dc900eba72c91ebf32f24bdc5e7929d0999eac118e2e0f3e6168f590cc45fe746c369d40fc6353c89ca64ccc38c2b23169f6571f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h405201c981c4495b6ad16ffbe1ab3c6490ebd497a36c1f61c731bbcf7bc68fe10614ab3536304c19581c24a54e27d26ab3fe33889ad8b5db06592cf01dc40d48bf509a078bd3cd218e916d684d909928e47c7e8d1cf1a4be8c27ed56f2a69759e792d056fb28f4af1284f604f15a2d5bda01f75397cb286bf66435b0deb3481;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f37a65c8d64919eb0f85afbd15bd49b37b542d5fc913e43e768cef9bfccd6b988ba19ac9f52b20eb3ed467e8a42f6c0b0c82f25c6ab2941620d11c81e242c2eafc0773479bb79e6c34b776be01d002a5fb7da071dff17e0299e5c46be98f4f3db80e3da2f4c1c1fc02373070c68ad203cc97502fb2bac58ca85d5c0df03ba00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1445e5daf660794b0aa77ea4dffba3e7199284525af4c95dda7247f25704c85c641f012ba92ac1c9a879dff89f16669e8644d80ba42eec3fbf9e654fe10b05004530f67ed6dc28636ce8d07fd90da66ceedf2489f47e12ca98df55b2bde487c20b8a832aa9a94b03fb111c1a9fb55c835a30fa5b54265d9a0988d21490209300;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7d31197ce0bf4079f4be9d42a27e128a698f54cefaf1ae935c0b038fa69494d20d7e0b0cbf09513e4d1e3bdcd562ebb23cbe21d07be4ce2aab5839c14e442a257c22b66c3844a808f85a2219ce3e4eb714ee7cd65aa1940437f40eb4a746936ab986974955faa8ebbc31e495a2998e65ce43c82cf4c04d08cb54cc75978ea3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bb2da1596a3fb67d99af1f2c436676212890b08582f8cb256c007c536bcba2bc6034e0b4f602cbf9a2e0b9fe3f3473cfdeb9ea8cb7521ccbbde9be9223a51d7512c10eb8b050847d1b65280693a289513400a7aee982452d8099e0c68036d7f45f852a164f8d31e8248ab15c7bb936de07ce126dd3b904d4703e53fe0d82ac8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c73d39f0b47980c9e3da53ad2a1082b3416e4bb64476a47fed0d4662591713b5055f84cffbf4c976f2bb1f7ff1826ad2245a0248661dcbf0d92902ab7ec0e39521cfef10e7d3645c01036b71e9fccc61ac554938e2755c41a1798d3bcf515786b558f3ac42da9344e745f7022661d9a9c1c75c837bda75455509717cda22617;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h409c8543429a01a1fcd16e9bf1d50b27fb322e03f0404309ad7e02d746e48830744482930702cdb2f2bbff83ddf0e95091020ca91f09bed61514a4298bd639da9b203caf3e5b3d5db4594f0bf7265fdd79029cc314295119475dec533fe497eea6bad8dd1bcca484b8bdb2625e94a0527a8d061353209a466532de99c1d5ea77;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f79c4e5317a6bf5e65417a0468df9d0205c586d4e0c5da70fd048fc6ad6d2bc90f337f3fbeec027b16685937050828a2038b8399d747ad3ba09a6af38e1a872667569ca5c3ae07118b4189b01656a903fc9b56c86970a7b6679c9054b7165513cd7b49078208e1e8369bf03cfe752ab5ff6068531f7dc629465f594f15969ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9a368bc51527cb6ba79e62b49403b87540045f2054e9522e87d1996c90e9fc419c474d8ba6ef6cee0279a3d5d20250bcde1f575dbf2dfcef29a062b3a80ec0f7cb031680a84625a210ea8a35c462d9b19beed19069946a0049129c0fd84a8fcf1fb8825f89bfb1b165a796e4b592045d71346efdaf604c50d13b10d8a6d370f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c2685748bfbabfcc703ff28497af3c9fe8592dc82869afafeb0a9ec72396b4f6d17d3f829502f73338e50f6fae68ae2715a2f17f9e72efb866c57da835f943b139708e058f5c9bcabd088527bbdbb1fd8e5d5fd7042c9fd42e184da8d925aadc7997652af2b1ffb28603688fdb323caf4a24f26fe02ae066df9361d8b188be8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2aada2f67ae2b6650aa1b73310f81b297918f14ed20930f419f9b0eb4abf01094a3bb4d1ab4e648279c7fd7fd0b0a841b2703546bbe2ce86bd2c220d5e310be17e265c6db5ba8bf56d644ea3152ad9af3e4adf4062c1d0bc28707ceeef838422a5ce10b2664b14580c6631c0e947f363916df163518764a46e49a1c41914b867;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf570bc15272d43663705ba4dba00f16c40062203ba7c7f996837e53fc646a25bc4e7de3fa894ea45c11400d4ed8ea9adbcd076e873852bfc032f466ec1b4400c3b1070b322f13612174a42c152379e878e92d55ab286fce1d002b1c50d23356768fe487141d23ec8b77a28d1145ec7c0f8c9637105948d997232b533871cb78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fc3528df3c11059a291fbacfaae31d8818d89c5f492caecd240120ed6094fbb711ea0a2c2b9ec582c2b6503d80c15c2686887a3df025e4cc1a9d2754b29bfeb58b20b3692e7980875fb862b288d5f0462d8ea0fa095d9c53aec45acd95ba649dffec4e7bbe6caebd9b2cc3c0b46008c1405207a06ba98fb582421da52756603;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a747732f1f67c373dc1b65f5d7ef1902977990aeb210b60354bd0b9f94f3a9920e0951e0f5fb7e00af7038bd546d540a4170a1e584915b5c0d133eec6bf72ad03a8acae095b3e40aa8d8a6c7e12059549b21c3ce0cdd8fbab0f5637bac5164385dcdc39279b5e22af14123f5c36719294a4feb4d7fed10b9ee270243245a250;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee46134ee773f7fdd8f045f82f53058c27df0e7574a95a2d1bff92cb0b468dea219b18bddca4040752895eb5ea5da57f5a52dec7ae1ffccd332913c12019f1affef4af066bd2cc70a478338c7f702d4d42842cd67fe287609ee620d906db9883fea73c0cd49491623b2973d26723d0ce8fd6735516fa668759ae0d4e00a19c2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50bd24faa49e569926692f213128b30274a0d70132e7fcc467646aa185a2e029e707ec61b7912d5944a414d0d0090e715dbaae8ac07415467c6b1cc8b0616d554e9902331b83f062e9d61824a6776e4b9a5a8e85273eec72b6528586abc01aebd08608937f64b42fdfa6af54bdfb2cee39ead2adf189dc599d5e612f94e4959b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbe81bc1f85655c6fbc556ec569b4f3464a443e6c8c2a2939317c393cd9f267427f5b9fcde234ec595daa2651271722113f14211e6514a921a483504b6cf686448d456f1413635022902e1e9018e1c5c1c792ef736bdedf2e2d237afc883530d8e99909ec6529bf41bd607692849268f42d0329ce17db0b688d72703d74931b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb87130df4c34cdfba0a915a4eb1ee4fbf2e41cf6ca372bd8e942654968c50592c0c67b18be62afe0db44e2236d0fdab8cc3b95bea8cd2c466bcd90a4b902f2df8b18bbef4bc5550065c6ccffdfb62e58ece5c9dd55437f2d72a314c8e65a119a93aec3792261f913e5aa6e2cdf782baa6210e0dac15253d0070e2d3705b810d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h284badbdd7d62a447d3c10287cfcfe1cd3e8837209442a0b46af42aa6e88a282096d79fc1ffe10782a77846a278035409d69d82ba1e9721c4ec7163a395c37eae8db9ad4da728e5f2b4aecba4b6e8bbee8c3d726c05ed138ac2b2b91166de56ac9376342064d7a8d415c75972c68ccd9462fd0f7c45619553a3cebd2c1d282bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90505dc621543e2cc83b4df54fd28b58fc6751697ea1374b523f1ad8fa3df6bd7bc8b16461080391fcb6c9e7bdc5147a17ee9a618dfcc369efc482f753f54c850a7483bf6fa29fe67687a07ac41f33e494853a64637be474565f5f98fa66ab4feb24eb995b1d8c269464f74fc088c810c52cd812988477a3560093478c62f978;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72a0284ab3f793d5bd77c6860291effef18253a3bde4ea00cf1022e53c95c21534248af3258c42a4a58f04059d7a9d352a31597337c292a4e63fb3bd2888f087ca2c403ffbd95db630167eec36af03cd687dacf344690c704070c0454a3a245f10c38ad74089956abd8ab3b2e9c7b55fc6b3d9ae7e04f41027383e0b0949ec5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc473e0750cc145c5ec94e9280ee4babb5accbe82c2a713afddf6f795493c29a236bc36f05d38f22c0937c16b6f27bc0de4769c64bf36ef03f24da50d1f2e44e0eea57583ab5ec96061a95149c78e5f7edd65b1aee7d3ebce1311505c06b58bc29754ec4b9530a69310cadd4e6cbde47ab1faff9d183427d8ff563f28155f21d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e39f69bd8ad424e56cc97153c2f7737aa0f0ceb3ae96ee10caf3a827563d89f2cc0c77b9a2489e6bb581675158031a74bc2095e28bae6450fcbb2e32a97fbfb3daa435667d291adfa8e0cb2aae211625a1294b15340be72ff041f992a08ae86346d5ac990eb07c6b05e89f3a415d7d12d2ebd78629f3fdfe2f3121fbc4f4efe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13dec7ae4a550ecd1c66f75764bf98f55da8d5ab7717c122cb3ce87b3c3813309639657ff2fe68cfa4bbafd75e5f2939a9aac94ca2144fd3154b8f2912735fb1f2cd1c594c05de986b394f03133400a03657ed869a19aecace27c54ef753c38236ccb55cbd57d9e84e2d8598fa45458cc144142e250fc7920725c0d85b284e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2712a84d73366e79dc6a6eccef887fe6ebf044871e4173c5e0980a8e5616f38345bc0579eec34e00820c086ac1f94510b53127b16f90289cca314ec46b274d147dd93cce68be6cb777205048bd89eb69f31175adecbcbe25c9c2233f539e76cefc35c6465b2b524a199cc1fd5f7fc464ae0d92efe2ca4c64742c7c00c8a01d4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c2d4cea031152c76f64d17781a26b2e127528e3cf170ac40957a8e7470dfde6e035a36948847706800486bde8def10896d546a741e07ad1f16e89f30c42df4c65589a212f6ed3579c485f48ed2bba30ce6043a370305c923cf71e7dc110daf582f468d965e4a4eb06fe892c79ffcb3ad755c062cf1a38cdd7810fcef9df5e31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3edbfc23badae97e5b2a6b857a03844b14a9b676e2e85250f0cf3abc5b8ba91f48275a2da99de2215b6dd6f06dc14240066e0c13117eae94541befe5b78f3ca7b7e9f96db147976b85c7010bddd2277d2b3009a71333ee709a719f1b7d705e26824a1c6be4c533ec4538e3b2e305af0716bf7d20fd751dff3e500bc00d4168d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf99bb3889984a6447b9ea977f23337d04dc45e4ee101fe0e0fc059b9aade81b612967b9c56d9b818093970ddc02ed4b11cd91a77d53a881e12df7b85552c5e8a20ed6c89c4a7219ad955e26199b8885ce78ec7baf1d9d8162ff7f1143e7a42e18e63bf04aa597f53cdc94354cbc3918fadae7f331550a8cbcf8125b8efa842b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17f641f4dc8468b1557eda2a8b059e39a643e42aba6dd8dc8f8dd4e4eeb7725624cd3532b61e37c40866f3acf94fd3c6d01fff2974f8dbcd8770ed4f1e7519ad3beb5f3c71a0b43178180d60fece778809a37d7648d4f8a33010ba0236c5bc958190ad41295e8064f02123bc2cf27029cd7e57f99184b4327ded8ba6383d9519;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h763f96abff2171fad24ca1c747a9a4b83c56e6946003539e2623e57a67fc591634e68ed74d96a8e5a972fc4bd59e37509ffebcd00526af02bfb3f5a7f94552681e905b96be5c39b8f3b1d6fa05197fe0d8f106f36fe02cdd20f6193daad661895297f1321bed6025379a76e270ddfca06c2550753ecca42bea7be759f112f1a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3094bd64dee654bc2c7151607b5704892520c13c878a5557aa98c6a8a3c438df76ffeafb32797bef84fb14a971df562d57d18ffa5464422dfd5314de5200fb0bed02f3de4ff94c3671429b82adf42e0b19d1a636f02b081ba9dc2939ac87269417884835b34427e7d124d98ea148778fa38f276ccfe682966b397c4d0a514d50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb0d618d94825e78aec7432cf884714b985d76319c9f7fd803fcff03cee15410d628a8897ed91e99740ca65b00ca91438e6d52615847b0818534263788744955bb5415aefa9fdae6369a6677d2f291f6f39698fbb8ac0e63b0080f03c0304362b57b2a67669a4e7df6354420b1006103dca5ec7756acad2ce36b3c0b43f6f966;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb604b239c72c201a85f121914a0d79aba653bfd4a38038d74306f02575097bae944517ea53b1675c86e4ee48c2569dddb69006447889efef92478d6261d3cbd46da62e1ab89fb8564c429fd73b6a3cc2e3e5bf044e8d6c22cd97aa252f4c96d918566bcded4367ff076bf062729c769e014e80bda9483c230f17badfcd2f53c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28ad3ee15f53621bc116eba1b07e9d249323403a357ea900df0aa4d7090231e0cfe1bd046cf9bf190d825692984397f8261d5e74b95abb19b2b966fe7075018771d35655ba1a100b15a90c997b2f0e6d7f641218ea3fe998d66747a99e167fdf412068fd9495b1f298668876bfe84d06ba0de96e32166a1fb1713919204fa380;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a623028324eca3556ae4277378b582f6639ad2dd89950e3c21b07ffac1b45567fd22cd51af4e9a8b7300812e0281091bb00e8952c9d7b750ce37d8c9733e5c0a2e6c8667f3cd08b68f757ff045ee94e33331bd914e288c9bafcf8406c4f0631f893820073f9b3306b54dc09dee60ebe9af5a852fa7d867dc8714b86e4c4ae16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80974f4cd341d704b28e545e05661404129cd04952136d9bcb5624d5247be977f4cf50d2a8a887a29f770f5d5e9899eaccb5d420b90f52f197d5ebbf87a599b8f819b0647a96b5a4d0feb76b5c4ede73cf5dd15609cfb20544f34c0b512c20f66fa22a57656e1fa6b04f646fc5262bdfb2e598897d285761a3ea0dce16cecf7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5218a773bb026f984ce04e536803efaef3043e9156998434c16704dd2a166446a7620499b519c3383d18ad8a34578296a01293824c55e830583cc440490f32f94de8e03dd446e47975e14f5b718985e823ed75dcaa0f6b880b9c6db320bffc62aa75d2ecf2611bf0e2ec1c439cb31a2bb6a527bb000f46746f94b99dbcdf24e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4154011702157378a42ae36f60dae4d634f412bc7a754eb8e7b493a30450e9af65b8845349487c03d58b76a8cebd27731fd565507bc1876fdb99c5c76dc7c5e104fb97c76ba36b32738652b92971bb49bd9c0d0e8980f480df009ec67bd3b09d32e6c39d81386d98402a989af788af7c347d22e2c4ef9a2ba3fa8ec815c9f1de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43379063441560c6b7e981da53d49fb8c11910b2bc2aa264682982652517bef47b41f56740cebc15822358fb4821512c0b395ae60d21d1bc3601c88d64108215586ba911722ac6281c0d1b3ece0f709703fa394241dabf5efaba235f8660145535a2353b54501d67a89da65bb09b75df9f68b42c0b3f1191607b3c181b8fb267;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h849f7f6d7ec86e53138042a97c4936d435cecbf7e19d39bc70f51e5cfd8c919379dbdb7a8e8202f3ed62ad41dced6caf4f5d77cbe35355ac4031f31408767944384c95479398d5b63b1a8a6bd992af393920ba19ace14ffbf28e1084768516e62f2b67b0835480511aef4d2d91098148a41f82ce0afda425009e1b197e4b64ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b393326278e48f6d3ec2d6df19ad81f07620e12e4fe641f0664b9721c7f9c75d81239c63ca98a172692da7451127b37fc2bf78c1c1c554e4ce6f8b794b9c0213994ef9c5f87e9bba5cc7cf8d76bb10b12e3c917fa21a35d50ff65eea8793ed98ec5ffe507c7a3fa05c82ccaf4b0c999ea3806444ecef3579d6a5ac17dcf2088;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52c6ad713491f256315df27ff2d29f4d1cdb89ffaf52c4f7b032ceff985ed2588c271cb12983a1dbf76817071a1439bb15262958aa0794f1caf91284e8efab4d1e95e6e5cf1ce3b5914d56fcedf09259255cafc0b6a22e6af182dd79e2c2e232b077096cc46f2017e7f0b425ad7e274f6f8d383eb33dfac345ccbe6b49878906;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cdd76dbffd89b231efc44173b19378ddf179d7f97ec2129f0f0e675ba9c51ab67be834d004b0fc0676f21b8d252b90946dbeb0592215b3f43ec23533ef88a91c3aa57022bc061bd3a4bee370af6b896f055f0c29b734fa71d95ee083aa71024ba702051be0658b7c3c2d2b0331c119788ce5392a0add52921d5fc7cc67226a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5f9f7f3700e6b24329a1ea6500f33a84e5c29d3ecf2e9b4206f75eec056118b7aedebad52b9c32092aee3e75aa6430b2390759b8035726a255e94e249af03166fe21d76cee4d2d83ec9ef801dd06f81de0e3f432a8842c37ca472a528f246a8ec5d935f92700fd3e34efb9349611e3ff8283e7c59afca3c807dc0cf820219d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf63b0ccd536b3a04d196f5013455b6456d4029ce9aa709fc9764a3c34651c5a947e20010d377946abb2118bdc16287dc9761e811742373c8eaef42c95e3c05f7b3a723bce294089cb27c5787a9ae752beb631f11c4cf62d8986c3fe091df5d279af44f23386bf233a9f6ca921d17a729b3f4747c236ae29b7e1303c811c88fb0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2d6d4437bd5789f8f76b9ecf82a4489773621ccce9fe71ac3c1dc21d6c5eccab7cc7348fae9a91c11669d14c6b66028fc3798bd28f22685054be165510996dac36e11b6801e107e3ecebb931b7828fa9c5fba3954d22ab8d92e8c09146b93c1009a3e5e05b65f227791960fb4e9faec3d714b33e3ff4005e423aa84311b8763;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcddd0cf107740e367e9b9990aa58b16f7ff9b4d4dc10a2180baff8f6e5527d7da0a647e3b2871442ead3f27392d4bc68111b8e0abbcad0ec29d0800bf41c8491064b4bd9ef6206ae27c3bb4af197689d9e07f9610425ca2687222a0b1e1321382e0f92f055c02cec04ab50ed4ef75d5c8d658255e0616b874dbb89138548881b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc069cc672ecee8bafb3b0308660f4424126c06db19179cfe16fc52e59fda2ae0a8f5db375dae7456c357131fbc32f49976c6a8246a4eee92f5d586263fe3229138a103a27375580d3d3158851d2bbd61c2560f64d0f1943eb16ec18e5a0fd832a7c5b386a71619bc87ada8d7d2edc7d2af40c14ee90192dda69d70593bc51fdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bcaea66dd7321297a9c76837abf4d4661dab9467be6bf58b8441496537c0503edb90a5b50ba97247800cb6a1109283ab0d7aeb4c8e15cc31f585984a74f954d8f038b34f919ebc9c114b68dbeb237bd5bc79e7f13dcb10a75eaa0513ccb9c98da7be991555f87694c7efa31126af24281b0d8b3981f6b9dd19b823c5ba1a224;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h373ea7eb9d8dcddf6e6e1f861e1678e67fa1418d7a58ba443073dcf01c6fb867fb781586e03ff79da094384fb483ba296f40498435c57cd31551b10839c8bd1acdd85b1aa0c155a3b17a7dc12854e3495e47f94441ce0640831bd3254f13b207359740af7be4b1b95cdb056b29b925bdf0c6eb4e8645f0c278cbefae8adc876c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf09431a084152dae887db10a6113ecb587d22436b67986814bd143ee322d6ecbef2f01aaae9eb0ae0687cdb6f9af6df42dd641a542b9c1ff117cb3998e9139605926c627ea8eeeb543998499cf668f8d5d4e1555eba70c1a8b22591953e0d0698f175f52ab8929448c8415e7c6f10d7c8430e09c66627497626ea7dc96e0ac07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h210a0e2ed31bff21c424a217fd1e4ef1b02f5fa5650a1854340edcaaf863b4f42df1460256f1ccacceff58bf206f9512a017c90ed613c552e22d9ff74aa014f24ab1f8c1fa4078dcae36065e5529ee800ba3384062d76520e69af2aec0be7336013ed130ec3a874d293660846757cc2c39d7d2964122d769d060b05d91c0f9fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5799b98f0aa25ca9852c9a99d1cf8dd201f2f450d3bc4e341fe963fbc3611cdcc735e32bb4a54c2e97141966bae3071f9682ec1db806f95c3d1cc37ea57dfd962ddb73ee6f83dcc015dbfb647d9c45d1a35c5819147ca5b02bd1fb55f8326ac3f83abfca76918f7fb6d897e2cfd46fece6b8abc107a81e83d1721036c4c00ff8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h845ff6dbde6a35b53893e1a7181b8460fad02a67d26d6d1f7b72c41644c08ce3c672bbef67882e1dbccb76b6e2a1198b48fc3a9081b5df5d15051ff96bc18477daac2639ceebe43e29ebdcd2e4a51424745369c4713ccbac951524cdf737669b6dd6d276b13f4cee1b73402234d11562902de352cce4f961b2f0f21cae407188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6265eba2bd338c57d9ca9cb5bf84a4442e5de4b647733f80a59c7b8f1c021945d6413a9b8ccb104ededff0c53358534e878e473aaca19c44f48918e84d20af3a3d5188df2529d540e0f94d8b34f018d64145bebc55f9d7fb852e7b67abbb483a257208cb6b902b5a10e7f7fe127733c421bd05a4916d3b26c74ca9307717ac38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6302bb656978f73213077b334daba14d2179818522593bfe6129af1a0cb44b49ac96b68623dfdd253cce7831b720f1ce47504293bcd1dc8bfc09a774b845da88dbc471f79202c348d4ca40c1cd4a3bbabc600d5762881916a869ce731cb95f3e34120c2ffd7467d04abe0bb5bdff9beae956c6f4aae378db1afbd0a43e12d42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98f4e8228cd92ce93d7c41191b8b2adae393bf87267a08aafc844a682ceda326c66c58a29899537381919c2bb6480bc2b68cb8200393301b7baed7ebfe864f286a3bd25cef1c96154f1c72486124f5cb9ea31f9c6ffd9fe449e619b6f56424da24d5ae8be50515b9ef354a0454112adc83cb114f4ed12de89c7c64683215efac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc84f211ec6d6c55734193024271543e1adbc74da7ad3a0034f50dddf3788ce29279f424b3bf61bfa0c7589f7aeac06246e7f686cd4d8d3bf990868523b8d40ee08dda4f3932ab3ce50e5fdb3c3daa353286fa76e87d7bf3d84b1b1e60c2c0e8f7de0a9fffbbedc579353c6fa2314d8b9ed4cb045eb78639c51d2b6eff87a643;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4e08077b647213e9c5cc9c956d4cfd6c9059c30091717244608531ee86340095e8b3152ef97d86037dd439c1f896449f217131d077633a45fafe2ac0345003ce4fa4bae58a70af8b47b337dabcfb807eb4754203cfc7832a2fcfb272a3f372d53e28a9b068d11d13bbeb7df120ec702d63b6f17ef451bb91b23c818ccc64b04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he497f5fe040815a952631fe1487dcae32b9ba9879356665d069259158f1bd39530c436de2b5deb08a7a25beb1f5be9ee137308aa76ec7baf4bcef136d81c414a215fdc00184fc5791edaa856dad7ad012b434396903eec7a1c9b383fafc9aed29272ec92031bbb044dd33403268a10029460eb6ff20f42ab355b50a944f2e815;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2217ae1b58a4d83608dbce9c9324b3dd3c2c91a83fb6caff7c419ce5c36ace4d2ed70c35bc4065a79919a9e0011da3b6332639253dd839c394d930794b04616153817786468438709c5ee60e032d47f002fead2a6925f7328c047841289e21c493d4e694c3a62f05e187b2e799283f1954622ba0b10324fe6a2aca8b1be32d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h149b97551dca2886bfa3f3d3265afdc8c126fcfe98ae1d82e24af22bfc2f39d3501e324b3669c4b910bab18740e962c481e7680c1f4216f9c00d93ced6b53097e5420b646518ec8b0bcac26dc8f775fc8735c9535cd9dc5392d47fbd8909ff504aced216b471f47dc78e03fea38b3c52b565b2add654bf331cb11f0ad6b4bb94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62de5fc8234c422fab7bce4e3807dba545ae4b0fda21ad02979ace4c75b6fc65c70e69e4e4fa30998e41631197ad4e54f0040372f5abb014fd2624cfa0eea1dabf671e6320d729f499871e6df3d4c732bacc3345accd2de9edd2bdac8891ef657f11126c630ff8349423f6af3fd757a378c6b6506c4e6f16273ac2fa37d64c0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ff98a622c47e24ffdd5715a72174289cdd78f6867517675544d98b04b57ff34e01563b0d3c48444b2389af1e08514ca02a1416a4240043190e6631bb6832a8c367b8a174de44fb5f0e5eb31e089747523e457caa519d84b0cde14af1a9bea0e41e8f344da7acc977baf3686e561e441b52e95c6ea3e96dc52533016e5e17be8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf63d5e231438c4d34d408a05e436c3bcf15418dcddd4b1abaa234b3ebdb0f931a50f014665dbf4913329fb8d883f3804ac6781da24ed5ba1c1b27ff28cd74bc73b0803ebb36bff7c3335537b95bad1c53e291d7162ee79a06fdcee0c608114ccb7dbbf7748cc3280660f8d48acd64999239d1db9ef0e5df974215d95d938e2df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58b748dcaa67cf50055a27e225525e60c395900fd19eac00d2e5265672b52c47143a8fd1b3fea22ebfbe6a301bf94db0ec18cf1ecf94c5c2c954dc94a5b3bce762ea6ac49be2f5dd845247a11e8de5003d3ac4975a9eacd0a7d1e69e31c460978c8a18c9c41bed44966b0c151dc1cb4482d8680c2a91e9ae1b88744705acd5f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb203b4a9205def7cb02b74bfa180dc290cfbf75252d0c366615800975022da9dd4d2fb76e8cfdfe978eff1b636f179722ba685fa838ad5995c1bf14c21769b37b020f9ef2cf7b26065a914035f938e58383a8425f16678d5c4713b1bffe7b9530542b4576a8866009a9bb997cae7f61ea4a9ef34c3acad300009d52737298114;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e04ec05755a80c8e65ccba4f30d9a92801a5bd87cf15acdbbd4653c67f9d2c15084868cfc7a9ddf4108865cc30af4a6ea4072b2d241ed5f48f39995bafb36e927b6c19534d4a59f17b3dfadac0ce973e5bcb0d3c06fccfda068d94323c5c386af21e1c98dfedd80d20dca76149b145aba47698429f2c4aa5de82dcd20215902;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cce803a23a184dc8de15841f5b495ca939b5c3f909a51e07b756543926d1be4fb1b633a7e037f2915b10e5d66fde58cefaba882f58188d42e862269e55906c141c821b2474f690800f87855c532430980f87ffcb613d0531f8071afe8fed92a65532af1a3d6258dacbb922df754b50efc0bf0ae4fc9977e806f619d00407206;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h144a21533585889e1945e1d3a7b258e63fccf6a1986b59f6844ec747c52af30c2ec6f7f36f56c23a294589d88eeba53a0fd84f991a5ee738534915447207bca96f2d4a0361453685999c2f5182f5148a350f1182f0d9404ec229e7fd1af011d91355e342f7773b240bc1c9180201c99adf1743c97f738334da7107af686d655c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3edb7dcfe479522dfdc1565c6e70ffa28e259b107790453c791c842f4fc75d5e12204e365fba40e142e361658c1e8fb73e54c3f1a80e96c10f3afed783e8d0cb9d4de473b9bbbbc18e1445692a6057ef66930d107b6a8c210b06bf6efccf806634e756ddc8b63f1a2a016d03f28ac5484b231b94a70d14d8c95e4461b5099af4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6aaf3cbbd7c04f401dd4f6cfe785cf86d2133cde6908f23d5641d7f5b9a94f852ecb75a192a024de05ff735c3778294cebbbe40a40bf13a0aa028766c7edb61673440a3b877ff18c20a3df1c0a2d6a9692aa5345d4a542d9be034eda059796702d311651bd0126acc1c63a698e44a9f23e25b747c127d51391d121009a7dea09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10e426fb4506c3b9ff13901c246118247c29c28a55f8e4eaf54b32927d86cc4aa5d5ac03f4e0511d5a20aacc381fded909f52785c3664eb7b29a9189257e734be1db0edadbfdc6f1517eb3abe93fd095019cdf96cfb5df3e4d3b23a729255d65a123228f6f4950c810846497266f282149c6d9598d532f5c3adcec26c6e815c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae42e16642e564e63228ffe1e3940afc131e8ca9d0f1bbf9c87230a94f1c6e863c2651877b0d19c77568606af79ab49dce03ac0ec1fd92bac0297fb66238a61069b30bef71c2d0fd60219fa824161aeffa8984eeb4103667dc87917e98fe7d846c4912104a077c0190124d50ee223980002df92d144033708177003b92d29890;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33d47a34b0cfdecdd28b3a11db2e0777a8de7f9c7aa34b7150e896eb0c1f16ec70c03ca96b758a617f7649d16102e03679b355836e1f383671e4f7a50c71437639290946dafd92ab1af1661a5cef6095f5243a2d03b7b59e8fbcfd03f344a833c7e1587797ab69cdd9be626686c9a9a17d59e29290009156bdbc18bf48cf8c36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he17c185abc6542862db292cd08a02b118ef0ea056dca91260b9a67fed021a487e1690ce830ad515cbbc59b9b4f2141fd0edc4972929280c024697c6c59bb9888c7f6e39ac87ba64da9fc670ac05ca1e3245a9b63b09798f07339427a9ac9ca7bb6b32b598c7470f854d21c435fe04efdb22d6118df8e6f40c5fd1e9fbae93603;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21e1b9ba62ec2846b19278459b6a314845c8c0a922581313288f5f5d924fe3cea982020e5141e77b56235b3bb1c0817bcbcaaef56dea0872a3b7ade333d1376564464e1c22a6150196d5acb2c567bd0fd0db7f61f8eb734bc82c6a470161aba725d699915beec39ae0a1bd048121c403841ec388f74165f745a8e74cb077f303;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99b4b0062ad0c93da225ada64b559fe1a68b422360fac10024a9aa2786a76fb61c4dd45ebe38d5dd46049a190ba0f516ae58490d07dc6a4acb25477bc42cc1e2167053055d5ee0a6062e6e9e2257b9039dee7f51d8f3a2a9a52973c3c99b903281f1989959f39f4bdf77d7269f49c93ebbe11ac0559d4c2d87f8d2f52ef12666;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc38b72f6bc7a96c3fecd384144600383135141c544128fec2f56f91ac3011aac52491158269efe3291ec2931e75f24b61bf94e3861f381289a46fb1d6ca38455e87615e00ff3620c39772e31d796e8924e51f2de1179f14481e298cd8a9eed7ceeb8579ec2004eaa5ff98c2f517c12a776248994868ece573ccdbcda40261d9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3801e9f609c13103fc0301047b1603237d86ce8e2c62e1a7c30f9ba448ad98ae5b656f601f649791ee52ebc3ecb387b9d76f93ae08c931d26fdc1310757f0a232fbb9004fa4e9af2a5bdf87dd3afca07cfab934a24cad887d5a0a5249bc282d823645fe7802db0f6dd16d68acde5a916f07b504812179d4b58c6fa072e89de9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96f7ec8e4c3ed646e6b1d5cd5c1b31a51e79b70807c39de416e2d6dabaa4db70a2eb09b61793957f42bb16b3fa495be5a95ae2efff09f25f12805bb406efd4d98df2ffbb9f4a648872d102cdc6332efe87bb9d288ecc82da88d2a7153d43ca6322d3578d8fbd43e46e922b70258e1eb6a65b37197f4f8286310ce648911e5b3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf973eda40f6b327eb96b142026bab8fd6d48d5c05e0d61e1ecb50b132225e83051345b01dd00f29d93a0b0e87d2a65429d45036977af9ea3f973e5a32ab9457a30411b491b158da0068b0596e4c1038aaf88f9b3adb38dc9d0803c962153975cd2d30891119e2ade52da93a08eb3cdad187cff5736850ff048007ef48e31e60f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf40a1cf4e9e56b04c2556081720c37727ba3b5fa659f510405248b045e62effa04039812a3f52642c87c150b845b3ac3a7e5d648dab1657f3dbafd1da244f43ada137eed60677b3da1301815d6affb50e3a7be450107f1881c9ac80c8c3bf1fe2aa39d4d805a03bee3a4c324bdef4edcf178cf43b50d22c9bbb6daafdbeb99e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bb09ef21539ab0dc32b9dfcd5bd62cca019edde09f1ae39f118d48143da1e2465d4683496db0b8c5c64c9961ccaf999caf7ffc3e77e9715a473594894c81505c3381013af4ffebfecabca710e78bd1acf4d65e5b33e63e890593c7f99e47ce71600a64088006262c155c8732e259f706126a3c9a033ecbabfb32d204802c5b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h974e44320e80942925b0bc258d233b983f153f818d947c6622dcd01fc2e8892477bff04cdd2fa662bfbc906f22db8b124622b917e627b28900ba0401794550ed291f99cc439286250f8ecaf75b6a0f55aab2ae99359115a2c391c43c9e637a410566a2e447b010ec88d7ab6a4200eb9ed9b0866f67c1b02e6dbeb56b29240291;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe1043eb436e189df96cd74472a2d6f275b6552b6f813c835538a2fb1d0e9dd78ebb12e749a2e4309a07867698394444e28d7af07e1cbacecadf7373da10cc1ef46538268ad2ca49439947cedf79aae81a2edace40ed7298143051bdf2edd9f16cc1a20d8b16db5de4953392a540af1d53ad1495087842f6a63531f5c5578bb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde857cf0eaf607ea2b45874b7effb9ecc74e44971584c008f09f7843f33f0606eb20d4930e8f54deab4f7f6232b16edab33bfb64157a896a43b4a5212528a074a98aee9e0b7ef9090d1adba94eb73c4d94dac82abeb156387d1349ba5c3790fc22a5fe6dbfd893107cb16fd745334a6e1720fcdfb6077f2a93229a2aeb8bcfdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0ab140a400ea73d40ab3525f34690ef2a32f464ce73c95bea135fd90ebaff6dfea17a409a4f9cb5e223071cc55033070a96983c0db76135750d236b1f77ad8daaccd2542765aee1bf49f89cba989777bdc752561f667bdc2afd6a78bc609648ed839b53f882d16728ae90eaa38af8b717e603c15db67b30a85fb38d77fc0ced;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0bce9111ef08f9a3855d1ec3f397e51d0b80daf1a0ee053c6fae126cb4e15ded53826f48c1e70bf65ae9b55debb8884b0798dce3e42b79506a9a8dee1828584c556dec141f821b114948ad18e864c2992322cd6ce4bc5353f0a22b55b4782eed68314380f172699c9381fb14c262fb5d2b7e7823858905cbef79e1c8446b38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2db0417e20cc44b6ed3c17eb77af8cc33fda22f9b8914fb9e546b2cbee59bf3abd6c7d6d0189999f2874d1c0e667537d29b4b580b53c942d4dd128662ffd85d5402d6980d88eee54a8d71edb421b8c8012a6f58ba045d199e389a5248804906ec20f532b010288ff623e137a7aff1a71f674cc92b9029772b50f74058707d69a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc1ccac6e9b88792079d731790b38e11b564014177e80d7e028939767db4871a68a417d8655ed83c6c28e6bdd5e499be410b4f0fdbccd548b59d54972306a9f90310bffd19f2ceb3a577f5f85e65c08d3f330326ad48b59b84b1cb281b542cd29f8592511cf42cee60347ecb59b9a9dea3176ef1c6a45ab731f93fd599fa3cbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd4ca5f35a175d6b7d4525cdc682704795ad8e807cb5f69db90a9cdafaafdec63df62a304c03be384b1f18ac7e1456f172ddfb4e83efd2d22afb93abdf36c81cab3171b90f402ee4099803c3d02706475d45f59d7a7590aa7a4d469e150cfd3e319dbff50da3f540b58ba7897101593a37eac3934ef6f237b48f67766b2c113d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f95e3ce39201c08fca97ad0595538b3b62cf07062be1bef0d49f77889c408bb123d4a6a038aa2bb516997a33667e31bb104012050877398252d4910dc8a1c84a4dea14e240f50752fd54d1817e896e3afb9d6fb54fb952f0b201699c07f1cef5686d20135dff3604a0b300eec563adce88cf111f44cfaa1bc51f9fd3e10dbea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b5ea80c39dc715cbf43387779c0f98e02c98bbc45ad3e956e187eff5e76d33ffa1507854f1819c8c994dbaa4f2320b5a23fbcbf852c81dce6cd1d7caac905ebda5fc9aeca1bf3aa3e89d601a976c70002bb10546725fc9f5c70e432240bb3a1d46bc80c85c01a7eb19ce9d373594ccf4115f8caf29ad0e8c01bd5574a3d0ffb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bb96cb1641f21aaa938ebc9ee79696cd1d3a0c1812525a9dfaf3abd2e0304d7889ea1577435b81dc5285535a7e4538da9d5bb36f9620eed959afb449fc4b83ba8db5e08d97821171cd0a43bff6bc4acbc4ebf61f3d0d9d9089c671bc7e62e379273d4d906081d602de7980fe345240586ceea12bda079e98aaaa1f9a0a20082;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7a07ba24ce8878d3dda63928cf6b91fb56eac90a84bf6a1b59b96eb49dc8fd58fd95c0046b9b155d6c08d064e35c2451c221c6b48f86170abb917061c7bf6f5de71580ed395d44dc27899a3a5865a4b92767767e99b0e66d37541e32f3962ad1ad1f85fad078bd45dbb8d700beaebe78bf2da4280635aeed75d076f330a9b46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8acb062c664bd677b67766773f2f14cedceeb154d970a452b878fc8d0f4155022dd283db18176b4a6cbc8456ed9fd486aed39e76822a9d3ca21782d667ba0e024b9557c4c50586b8cfdb21c0646feb27e470bcebcc9c3ad338698f096028441721b58d1d252a1396548eb8a3b829b978be111a46de4323efc56c5969c7fc6a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfceecd38975ba0838188a3299e2393baad11777c61b9de430c23eceb3dee5f80e8d60b32cc3c7cdac9f643f5f66657e31cb017a86df80590be5b2d13b624ce1f1ce470ec9951ec64879acea9ee6c049c109320c29e08e2c991cc05486095d6b4d6bddc1628c417844db46d1d3e087b03a4ad61913ff485237278bf8c58a00f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h100ef1e69e9071687eb71b82c22d684348b1a0a60ebdb01a577f466991813ed62ecf28765b363ff09e716815bfe9590eaea5a58d40e5f4353fe58fe1153a8dbdc76cf947ce939192b41fc9e61ee739c7298a4cbce73d889c56e21f727bff771fa2d54b5e7c2462845feadda755ddc9aaede1c90e07d63db66c940cc8786c44e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3647a558aeaef4d13f631edeed8e267656a9512d24d19bd24e5d20d7c84648c925fa18c944f3d683d874b4543b58e9700809f23ec65c930ed9db84261d90df3fc4db49f005b305275712357564f3163b8318e2a52e22ad5b3bc79e83344c510c94c148330d8a8f549587a4d87eef377eab1dfb1cd955e34d12c14a50a99a4143;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he08e71e0547c29b841dec5210a7834f5fbbb0ec3e39d6581febc39f3a4233a6221a6c8e9717864c7f4c295c574b52d2448650a67dfab219be3724afb45c3c7619cb211081d87f0739643c12e8275ce63facd00e09107899c559b448f2d70d2fc652eba9ceac53b49021975aa031c5c00550bc34af129ec7b50d34f1ec04f949a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f423ccd3cb4337adf92a2cce5445b13c1a33e96bf53d36c4179c952a7e798d3d2e5389e0081668cec340c90bc06f0c32cabde7b2fe9964d773a4fc54f0f54d5674db3fa8802b33aeb54c34ebc84a30cfcfa02696c3fcab7cc3e07d6631694d1eadf8add6f2899d65dee1954eec0e905da5f79b00d934190ccd2ddb0f44f4eb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2312b35637fe1b2c458113120b185714fc2a17b80c63af6604c2c60adc41becf1856d38dc935b0695d3a79501a8d2f89671525de79f648350c7949331ea1c973d801b4a7faf272e0eb962e4d5906def33ca4439319e341009a95f9093fafa7f416c1bee2292b0776946ddde7ec3601e61e41a179f877183ae15d8b1c171a85a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3385b5733638e1c92070c3d0d641298c1dc40d46168d3093cbe145ef9e3a56222a4cbe47a9dba7fcf63746e7033540e6a77b53bfdafee2e51a468c48c460d181ba7ef573110699fb14bebbb4ad21214a0ac3c88dd5f70cb0de279a70f92a0a9769c5099e65cbfe68b33e8c605df35e4dd26f046df7245ea9fe3d0fdd3d8eb3ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd104dca0c832ba40c751240c8556eede32160aedeed06d9803502c1a1984059b40d39612c9a8f93859b0683ed9fe84191e6010fc1c39e903b0e086fde95de166803e7a2e7114142a40c2678a766abaf266cb49175962b779999d5a24a41bef06e37789c9142b43a3892b3de3c2b14fc474ba8fb6c711ffe1e70b2c875f77cb0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0168a8687ddf6f6f981f7fc1bfc5b8f105da6a8c7571afde12e70e27e48f32fcb0a871a98c2bc4a43e7fde1f60dc5f3a1d44b87d723f43e38f35a3396cb44786a9085527b0e0cacb29fe544dfc1f5c6d35ee079636ae2d48133b4a161a9bf529e5ee7ae72ad6a4ce575c8d4f5cf88881824938ae3b25fba5c99cd46224067b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97d1f87baf3eca32ccd577ee1e55c75acac1d316e7c0c3ab76249c286dcb9eba2dc5b28daa9dee347022246b9180ef4b2a85a4f10ee8d5f0cb0e74da2eb17f53020b7183fd1130fd98ca8491206b4ecc78e954813d7d88875fd539f0645bb8c2d762984149b6101b48aa1dcff7e537921e232c4d7fe894e227bd0f01c4210c53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7328987795479c59fe67760d04d2549c884aa010d00dabcc6944d49e32cf17d39b50a53363035689a9825c707fe28fb5607d5f20931f9b662309116d55c9a0748f3357cef2a4bcd3f3854a631654f72542703a951568492b009d29a01ba4a631b1b89da339e32bf03893fe2c86d83bd4f4494ffc69d965489a05fb3ddcff6b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc49d25cf73f09fdf144a8e6724233d6f9bcf57f5ab4809c4678028ccb95e3798789d0907b26e10f15c5b4fc3c0e918d5c22beb2c2da78d60e6398121275eae73be433b7432f45735b06aa71052d0bbe1bcd27d71f793d99c8f9d0aeda416ff1b3408a93e317d66f2b432f27f6c2996ca05497d56d589c065f7a8c85007de490;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f29f7c0480ac8d58e1bf64a50ba57c3db7ad8fa14e258281f1a40072bac65c7ad3dd5d82aafad2d7fea603ce4d85c97105fbd06103c36d9a687e063511f778580db420595caff604b5cb7eb04aaf991a14c514ed8a4fbfc0bd08b39ad7bf6aded63bbe796dbc4116b4a4d2e32dd2b23ba01939e9a58cca0a93578e1491c9c55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89eb57fe8900c3d00ec41c78e637ab7c54321dca7ff870c908cc4ea99fe6fda8103e9b1a4c3063a4990dc1b00bd6345e4db77b3b3ebdb60c5aaa785171e46080f19e557c2210a3d98ba1a46ccfd79c4f15db175467e4741873f161015c0c7febcccea73dfbaf61d5677b1e82fb986a8bfd61ae2bb2bd2787ce77f15540a3c55a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb23ac751d99d0136599e43c5a017da35164c2b4cae4540e9ad6e0d456d1f61a640bfd3c97aaa01acd8ed41ff561a8bb97bb9e74ee8dce904abb7adc4ee061f18e92c05b19c6da95ddc0279f7337e9c5069b97804f18d33a9f231c05dcc90eb9c1f052cfd8839a1bf67c163c178be9a986a896f713d1310cb70525ca182a3b388;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8144c295e0770a9394bc6beb3feb7e7fa1832bc397bb83815483ff7948a8905adf7431c52a38b06b44d0d35f98de142c472a7b43a5f478e03705a18fa29fef1b37314998c935f302d81982212b9e4ad5c66a44f1796ceb0fe36ad450a8c7df5ee0559388f6b365db5dd7fbee0c2ec2b57b52da3072bf63175bac2ff5779b6ccd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc27630c6f6759b3c11fc56f8461d1e105198d1a3fce8745f9e58ba0967ae0f36962e55a93497b26282b2a9bfa9f77df40162ed2a7bed04062285f52e275a94ce13beaaeb10bfee8ed0f49b3fc65bfd9115a1afedcf3372d833907ab60c55a789eebe0ed40afbb286d260432435e968d5d1992d1f0b8c1612fd0f377993053d0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24e42888f026203846c253ce818a4ae3f035ea22c5fc653bb96114b02de60afd3a1bed361e06712ac497afdd47d8b0686f14a22482d8d81000436fd6e05132daf2203664dea439d1fffdeee335aa05c020b70a3e2f55da61db07d8f6a40fd9d70e31b859d3fbc7d8ead5ad2745e117dee39bf1a4f8d0eb8955f813d45b7dc13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2e265ccc4a3f39e84af6592c3654e1230635b7b33c786cf61f6bb7d46abf76bca05cd11b40f636c2cc019695033f74b22ced2a1cd9c40d94de5e85649868b9bb3c7dc2f1b8016c6f3f0716f7758f90be2891288c38adc37d0163a71dca56e893debb18bf40239a29b6e355952ebe2294ed95f3ab3b513322d00cdcc3734d100;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9594842f5e75580c0b1ed400b61e76ca59380a7578e9a742d01be2b7aa8edd21fafa1f96250df661d9ab8ae361d2f19fef1611dee5f6738debdcea9866598ccb6329564314e6040187189a130a3e6cb5e21115fe20d18e65bb9fac694443e43e7e486778a0a0aa9042716e044d24dde38dbcf27dceec501d69adb0989b4b6eea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e6d7973dc1252b60fa3efcfd580cfff8df9484cb9cac65433785307cc62b32a723fc01082536f3616f3856d8e7fc36a01ee59e5e5e7184895e0fb4c3681beae5bc17ba09ca22d50b6e0972cfc864ee5147d3a9e5e3ac56c6fbb6a562f856a8b6577f27efc7cbd8fb90880a51455b600fb74401cb619ea8c8bf7a2a069e131f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee34f21422484f5abea15a01f63048586cee7157ee70865909f1bc0d92705ba851de4508bab40801b1be5041f9d4eb25d6e6db55401cdedcab3db3e6830793f0ba1118357d1d8cc3546d0853e06c94b239040761287338d9da324a8e7f7e7f7197855f401301a28a2a30e942503329d548fcd5f67eeb269eaeb19daa048fd7c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87a2dcd6c2d41a1dd7cccff0c889a3071b1b96fa3d78fd8c88102cb31c0c709133ec462f667cf00f5851c21fbd4ddcad5cffa3da4b465a73d24a882671b35ab16fa31a8cab55d95f8f4b263258cd2edcd798f34b7cc36c4a14b4508127fc21f2484ce8cd2326764255ff8d09d58d39ce8ee30bc9c2483156dd7a57cbf5808893;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8223dd8891619133aa6fe8c8dc9e8e15bce0c79e6d0e4c10bd6f8b08853f4406fd0b9d74d71c4c48b97bc50a612f48eb51e239d3adbd06f7bfbc7da58cccb0b96569c46f9bfa799f19ef0bdffdcd76e9e44fdebfac670e72e0a978cfe9d62fa908059d4fb2e16ca3e5bfda2df0fd5debe5254395cea0451c8356e678e184885;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefe6be5d2fabcbf5f64d6cf376a6c6db99302c871e0c51a4a511a2dcb3abbfacac143cc5e138a76cb855b3d949cf44f9858dc0b0f7b80bc717b2252ab841891bf0477b138df26180ccd92c550cc278a9ff346b1614e780db94501cb2060beffb1263b2e43b7e408bdf03c94e9bf4666bcf5ef2592ba8397912b4534e9ee5aab6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h449736f68b0da42c567e1db6d88ecad09a8478072895a8b045cdc44f5f9255c638cdb2d6d45fc59d8b5d49c5c890a315b2b92e3ad97599f39007cc5d895793ebbbc67f3386e02121201925d355b1e9b5f4ebac662fd96d2919ecb35b7220842db3913b805da3fff391d6c83b852c4eea561b24804ca4224786af1110b764266e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ccac240b29d70d26467ff7289b0eed38622af2b07bc790961d01d6f4bbc7fc43401b43a635f65aa328e8fea9d4b8294f0cd5b4adc8bb206908ccef1044e959360be505518d2f1a19fbc122ba74b62edf2678846c75b6c774df3242a7f1f03bdcab3bbc6ba04cd00dcc0e77c0f6811f709d91d5bbc615c6a7fcde1a257a93f7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h165783fd7c6095ddeded4c2a87c63d4cd704543df216c497b80ed95f1e499bb3f3435f95435e281595781eac0d91746b7fa6fcf7637ed8e6d4ddd78dbaa00fcd97db4f0f58e36c5a23d40a47932ec0d95b8303585a25ac8779f7890607efcdce95b3a8b5a303a7e63737a997b392ed0cb85fd4f1d064eec113ca83a125c8413f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16bb6c931ea82be1fc579cbe8696ab6394740011639157f4e5ca5b5635b5e524c90d7ad511c19aa37c242289208fa8d6106625fe48a890b974574d608aba1620d1ac0798070c5ae15bf2b12caa0735474b944dbc4024b410f103f8990827b868c2582db1f2d8ed19f0a52abdaa6f35ec02d8444454920c5ad93e6f91255a1ea9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7897b8c5e6f41d6fe0b11400dc24920170e872dc76fb7d68bca53727870564de23c36be215c96b23e45027f34f56c6eb5a9f5332f9abca0326aae91a4a5735e43fcd38aad6457831f05c9dff15ebdd27ea810e0a10035590fe9dbe9019b11f65c88a0472f955f86d5b4091e79b72a5374778033e49631f87f6fa20ad76dc5bb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb719de6db5d51c7ed4c7527048740a316513d239c9128b5160f117ca81a7c1ab1c68ee4d78742a50c81300aad9b34d7702bf04f1aa394ca4b1d7350f60273a776aae1eccb4411112220468ed4e6c1282792d6866dd2916a0c88e8425a7703b6327821986f5c1b1d41afccf5d84133bdb7d4c4c6f6e41d9d160600e3ed403698;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h117e151c8d68b8664220dae8fff5cb6fcb7f87e982272a6cc34ea9eb2d44e5a3e05ee83fe9218a0b513ec32c0193303bd0566a47f5c43b08d3f671839c1e449944665e961709e9a297c6100db5afde4237876731d304a68362cddca44e6d20da1141400fdfb904e3d66b8c3210f27c7bf16ee1a5ca617bc4ef558096bec267a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21fc8800d8b5109016340bc41d08a0b0e46693a4d3d8d2a76510b65e5545f2f49288ad87ea53ad41f9b1d3c404f4d73b2e0f2c909abf425317fd06af0a9d84ef528c0515e7c4b19de5ce6c972f95e1f5b70df44f4ae79452f59dee1c54fe0f51d871e7256d3be21ff08a4f3a473caf3dd88726c445217463ef5fca65ca91ed9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61b5b54e89dc8c39ae4285475686a76daf30fcc4382fb7bb9edc8f80ef9e3fe6a662bff21423a36d817aa17bb106423dce5b2955c67dd002498b1bd6103a2a7c1dee71033a5801d3fce47a1bc307352c50202b78d64dc948c55dc252b31b84976ad55fa227b76ad653e40f00d9f0f49ba3ed5d51ca50c0ec7647bbf592cfa65f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fb9f1226cc3f4cce54f2f5dafbf9477710a14cfb61524753c709ae7c8ea42d2037d77673df9ecf12558b91b3bc082f80358dbbc0ccd0a81c833935ae26095a1dcc5aff8e6720960643efffb19b20857fcd43ff8721ff75381be9bfbacab6dcc895d1d45e0fae7ed6a8f97afa80ab72ec289e329e8b5c084b519848013f125c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb71670592adf32326f725553b6aa65659dc7594ffee3a6ceefa4d65556846e27d792e5f352242d209e2b5ebe5262864d5d1e87eae4acc92422ffceed9e33bd3acc1f1903f87c692c5c2c59d404d8781f4c089c0936ecdd543fde1ca3bc9eaa0430ded7abadcfa4343353b0ef1d724a8b537971032478741c3c801286970543d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h873a05d2b4ec4814f544aa73364631dc1175ce9bf07195294e8322ff30c5970812d2030bfef2bc88acaa537543e0ea3429a045c3d7fbc0a238b5a5f4f016b4c59e9fca6bf50f8739a8889adfd8916f58772a6b7a3a2c94330add4bd06585abdf149645257893e9712be07aa395452d19011f2f75e8d3a72e1c246e543b9824a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc74eb0c7dce57bc8a2e2e030e2061a5fdf667e23f6e5d3dc745e725c13a25fdf3140d99551d7154607a9ecf0780946c667a4c84547f06f52ebb609f715aa3785cbff5a6a58da92ed475e8df405c5c8caa66225753c7b550918a8ee691ea1f854af7e9d5c49dd84fb4bbfcecbd8b9cd546e2401d8fe58b05f7cff202d3b6f8a2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41fb6e23c35ea1daf4bf7fecfc45b215a9556cc6746cf08eba49f6243fba7c6859f01cdbee578bb7e631de7a73f36e23b22238753532080442e6f3b1ab95cbf9de30fb08906814c38afe2609b26fd5ccd8925861ffc56cd4e3dbe5f7bbf6533c952f4351f2e8d621e169f16a33db70baad1f7f07771f1a067abac1246024ee28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12ca1dde1b5c36e57a47b7a856278f609cc9fae7dc252b000e4dfa6e7683f1e912975335cac0ea0b809a9b925d4e97e65c468bbde2ceaa2bd10bebd69697d5d38e2a834da57a2c90f3ac9ef308c36984cf34b1a0419fbc48fa2b108d6540748997fee373d790751f2f742f8559526ff72e7709a7c5d6718541b2d1761a388dc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcd8cd2289b41d894f1d1c86e244caaa902dc34b797bad92cc0e4bfae171a050a91afd4e3795f6b1e9a37561fc2a6282b001a7e4b60d7703c93104afae0f4f8d199cd5f83483d9d90a1d14848757ce1a4e0165ee10fa5507f42aca76d5b892718c36af309fc3345a2a3a2f762615961177582ccf4b3ec8b14671136382454202;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he699764a4fd946b54d5e1bc0c11d7d53fa579d455d0bbd3c58d37de3e0bdc5975c2ba85b40e4b66fba20941bbf423e9168945543516ac98177e23cb98c6649826c2b9ebea82953e78eafd29b810216905cdd943a22cb5faeb552cceeeeb43a59a0c9d3ac04c02c825dee9ecada57f15653ec2da1bcb3537df11f89018bab9583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h569de403d55100005b79f3b7611690e8f0cd398a05ebc0a3cd2d1fe886d771f4fb8445c783b20b8f7f8deee2e7e03e0f547a9ed16150b22fbb45da21e8e7775a2039592a3d58ae3889086a1409534104f87008d675100203d146125710f5c1e5d615abcc373632a4dd48e950ef77eba54cc007f3b9c54d2460cc9ceb233da5ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde3bb06e7ec6102111154a5a7a1295e8ab0f14b1b5cd4d2017e455764e055a764094272a9e476ca583e59b7416a49dd1d08034f42ca795332e3e2de0f5e026f45bd7a8242c826cb0cbcd813b599e9dfc38f40186c007c18601188d768b50e6c606ddb3b68d72f28f8e6aec2cf593d5c136de5a83d4681d99c24947a52a2447c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36dd31f8b0822002beb5d7356a2098f83a082fe5271586a9a41d5d637877671618078e8c0625db6b2a5fb41838c11e2a63aa8d275a85d19bfab0a8e912c79e24f936611d245c60f2a6528069b1d361a09d79c770e26e1a11c2c2cb7e3aefe5f6e1ea1186d67d775a8a70407bfda2784eb6f53d3c53c9c1dd14bbe97709c2a67c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2761b363dab999a0c79b0940307651eb4fb250679169e098700e62d2c39e67b6c659dc2ccf9cf381d83cfc8a95585a9abe12f890670d947dd0e108dec34862ab1f51595320126caf6dd38ef3816fb92bc018846b89d75d7ac75c51f51336214c093a933f288248b1d02f2f99ffcf99a4decb6df496ffdc5380cfd620e50c4786;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef6879c763cf194ad6bbf83dfad1c19b4bd2b11e667f2ce76a36e496d71d0ad5236d945a036d5e1709ecd80103624f304a147b62e714f4903a79f6b982ea5fb88480403529d74cadb14ac8d82c0d3ed31783f552098d3a8edf1f263c6fd537bc3f027f8f5b2aaaa162f5bc9fe9e948c803bbc8d3d28f90f852aa65181d0d25e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee13ea53cdf2fc646e480b2b306b3cfc99e83b4ae94a1f7d07999e0c34b918451a24854398ff794ed57b0ee78ea14c0da440d8671d90f373e2d30447b5e37ebbd988cc5f3b365846191ab3b57e5d24cbb958b38dca528dcb05d9360ad1bc8833efe925db06bf6127cf25290d4d03b728570717731831349b70e50f957cd0b078;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h940879185005abe481c53e74e027158608796a55066956ec0317e6d2e523364019be11debff2119c0ac3227f482167ae594312b46b6bc136170934862da986e11bdd7df17a04b6b23e53ac4540e62e2c0dc39bfabe34e32860cb19438532e7d318d48cae87ae9c40d7a054c47ef52677251d3c0ad338b240a2d5e373ea886d51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec305f9eaad782ed981dc8461d6aa8e57a2e58c1aa21772a75acd058c803b084a7ef4117011f76d205e690ab32c483cb428f07c1bebb81322a33f4a3758057e86b15558a27c34b05373e51567109de3f7ceac21a7cdaccf10bb8ad50c9405fdfc180c8c6fc112c6c21046dd3fabe90b132f69d8dce505ef7b97e0dbbe2ae5490;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3d6ce88c89757e5453c0052e8058acdf758d4b6e209582d1205cb2d464cad7b2511c96ec5da0f517335cdf1748ad355800cfbeeef0665b43e4b533d62f62755f23278caf6dab806d9c651af3fc7c7c530121b475c4a6914cbc511c8ae2e0e3b1a61eb0085fa89efb7a63c6725a98ad04923785ba5b750afbb3c913426c81e37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27c5beb401707620348a57da32f2633843854c63e3d86494942b04ebfae8b7f718b3510b7c31b9bdbaa92aee6c62fb769363717dfed289fd69041cec143b67c1ecb5cddef6ec1404642bc7ec70e78e58d64326cdcd2ad5d35b5855b72af0161806611ab2554465a12e39fc965d8d5aec7db5287b624d460fbdd7285ac14e332a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4c4e070aad88bbca291e05f08fb5e88d824e8fa025137296dc6671a83acae4d0308d279245156bc19e1e0a5c2f1502cee939ef51bcb8a51b72d1ce8e5534eb17755ec3d964ca0c4b0c3d6a17befdc8de63dc0ddba34f2e656904fa66a904b647fc28230b924fa0b8831037ced7c7603763bd5efc76f7cda31e5a862e5a49fc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25eb1150b85a47c0772fd3756c5263487ed358af869f45d03051d49cbc473081c38bb4fb8213ed41ade410af92c102c31687efc38f9841fba5f8b4b91e349fc05542040ea42728b4817c383565a24a1a786c6d8e2e38f3246e0821bf2cb6f53b5e1e67b7b05b6b2fcd6359a13a931349853c5abbeaa55401d9ecaa05b68fed60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15431689304c4075b2f21b2653898009834cdaf0d67faa2c946f77238bc2700b7d5f6b5aad37e32482c02e027133e644ce74c611823a14e01689be71f13305c9c3f975290c7947b570f65a13a9c112c30ec910e0c087821a53f1c3db3075278fae5ac7ff30d8b26a5d52794f6c6a5e30a5a073d4d32335151ed298372601b256;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1ea3379c90682a55e49d45f1275dc842a2bcae9fc1c766b8bd1a52af698fc434df53307fb3271f298f21ded0fdfaa32aa724472e18da1571ddc6ae6367caa30fc3292d4164dd517349bce3191e8a3f98cc3e60556b6f06963c6910b6434dad320887a1f02529fde95222a85cd500b8309f3748017217da447a2e0410c2b7034;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60c8df9491896b88b9425986ad01a66c329ef92adb956bdadb594667ffb77cde482775a7172fad0bb73a962c5b8525a45b3a1f4ba82a58dd086f151f4a34cc155dd746c1ee6046072bc6b49f9ddcb2f7faa5e384dbd55ffeb00b9e031cbf8c6bbd2d459aeb89db8afb6610a357e201852e4ac44fee31e0d5bf34437aa9ce551d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbf2484af983018d6103b46c42a46c46b1736965fdc7104499c32d973d1ac4e3a20c3254e834a81ecc0935ae09288360d98ad19e25714abce59df2b59ce40430b2f48e4ae04a75712406b62406f0b19ffc6046497f4ad8939f712e14a71b4f825e98da62ca96783c15f19e9cb2647ad4c288301874507141f0e6bcaee2ce5b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h759876efea23fb7872b874e71cd924a20539b0af343c4e9c8ca2f199c838699c498b5cc086aa5e77716453370f4822984bfa259e5d2e876d4bafba188488341969e5424c0d5cf1073b77695a3b9009ec093c482e0254890e8d4536b5342b7bf95a7f2f4479bf8ca7a662f9920ee0327d93f293d43bd495c7bd0a9f037a7a1407;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61193d1c932703538e75201ae0e4531d5766d0f02cbda057b91709542d47a139834fd6acf9ecd9e48a13e9d42b0c1ee9d090644772c622f2c090a74bf37829f70a3945d91c879a29e35039889305bd48de1a853560ba4451538cce32025d85dd40caacf87d058ab51d83e7b169d43225d5e10623a8b43b8f16135158f4836ad6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he66a6b7cde65db9e7b3b9c56cdaae3032ba04763d3ae16ac5000b95e460b7689e221e59f3cbac4ba0ee999bea948b4b1c3e55cc83e32134535cd4957b913bfa403caf98b2c3636eef737e098e58045465f907fece5a2a72e4001f9a965f190a758d9f80708b4b179f0cc5ba946498fd64808b376c70fed9ce7c7f9fafae990c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfde2830940548ed4e0bce641414cf427f8e8ce57cdc3831de74f4c5c4f9ea95cfdb7ab1f96ae74b2d151b024bb626941f3643a2452e70616cf174ca328acfefb4237295cdcde2d61a34d19ad7ab6444296b8b106adac0242e4eadfed1902185d48149ee9b3eb3dccf621fe63e5bb69003236bbd43a5011f9f5d39d6234510239;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdc039ed99d90e7e76ef86df1bd7a9d98668e545bb479105734d2e3cba83652b5bda4bd141ec96cc40e260b6ccabfe08532dc446e707e158599e1994c55df22d0a8d8be95244c62c51b945fef5c670bd6101aa388e508ba505cc0c4fe3674f28410fb965074df9f3675e55f58f1084b1459486fbe8174b582606cb853e06e998;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15130c75ec62ab73ec321381cb5777459e66e7302591464070c13992f1548ba6071a2ce29b639dab56551dc0ff9450556d30c8c9c870fa76bb91dbef41b2417f12764d11c719daf49be7cf2d4291fb32c4884c277cda70d7c6eea52c303fac6bb104199490e9edc60c91fb83cb0256e2f826e075505c3617fed8c7adde5e26bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heeeef9fdbdb9930c814deaca5a4a60aca4789d8a1421a47a5431b42f73c02a318dbb539b023a33fad77b3004ab1c70880b910dd05f979a882bd07014a7d646212a5f17ac503b05168d8200669101d85b212113fbb10549cba370e67c2530c33a950fb98bbd8426dc29736ed895d11f6925041e90fda064706cd11e5b0cc1ec02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98361c945e2279d8e76728751c05a8a1e28d393ae51ab2cb14194e768229e4eb481a6eb5509849b7784716ddfe97cd3fe6cef870b5e9ee0dbbf6d1ecc60369290952e31db49a560593bdd2d05eeb60274c90c10d72297ad3d842c28f4e6eb1abf0db3461e95a872adac606d8d34dda3b5b5ced931756c688c72368e26c1517fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h277bd3d31d72898ebc734db42f22212a2334f47f3258965509c90e51f8f29d1cba5eb6efa2486411e14f9d1f06144775c3d7d4f5ecc4e310d56e29990797b27540677e7ace6624f8affb217dddba63c9f3f06fa1c946a467b5ee9852f6113c126aa55f36f68d7de7679e4ea952093b52626dfeacca564680aa910ddb0e263d51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea1b7fe1f38c88fbab85659b5946cceb44e081068e7a7fbb2373124de476d65710dad3a3258163ffe9719bffcd96832dc9fd2d4d9d4e288f151586460e8bbab1eca81296ea3d2cf6e020e8769750db876251cd51700db21b77e06cec3d12512548c4358b96d43a327ed13c0c45701cdee1bd82cab354fd5484221d29243d9d2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9080e6ba497d9c8c115102e58dee442189aa782e6907cc26de35229c477c08c314e0a1a228e311fd9e531fa31c99918457bbd51c3e24f399d15122295c0b92660172a2b5a80c47507a1e73a3be195b725ee0174a2c4d88be822b1c07281f99c5063094285f3b97f6a0a427979f45d703fd4d3aa8f2ca1bb1ae92599ac4f96e37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4508c410aafc29ec94983c6385b8386b04160accca643aaaa0b4eb9e5d0e20ac88c49412945e3d934d77ac2387f8ac897cd6030993dd6c66a7ab7d0bb10a0ba75c2d017386e52de0d7387f02581f94a4d98731cfe6802e3ef53026768605fdc66a24b9e89e1b201012052d36d4f0fc7e5aa8aaa90093bfad1618f2640cd7dc1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8d2fc70a381cce315860893595e8e82f37ec0a59602e99db337d1b56329f1da572503b4d2246f0b10154db0c17cf243cc27b92314f1f298f37975b157b1132a0f2a6601777b0b2c92e3a54630329189fe03ae6c996644aa0f5bbee001f43167f66d7ea2a2d01404c4a3818f68b6cf208eee481dd97d54bf9cbc6fbd85db78d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55ebd47756aa78f2641524ef23af00c9325f96c3fd2818ab083917c6fe5c64fdd211b5ad9e70c91890d40a5d8553ac7c293df92dcbedd08d2fa67d12f4ec5acdcb2c65f1dc9fb5c37678ff7fdf84dc5c0138b5140b97c1a70d60d22d62232c91540cda5ad0455245f7d93a9b148f00aabe0aeff8f382adb1709891830c8b7121;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ea2df449999949d552c7477ad50d2597825758ddf06a5fc557779b4ecb7c18e60f20230e577bc7cc374ac80500b91b80f786e3b9be28a40175100924f9ff00d90857f5220b52e2096f283caf0963af7e8be39066b7badf796a0a692a925d97d0237944a706ce207601759ba54d21e60807703d8eb9dfa0235cbc984f66eeca9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b371afbc88bc502de7bd32bb191656c795ccc3e54bb9977c7c707458a0cc0e4029fe9af7d9e3caa6acdd9c42126175994970af457390ec18804d634c77ff0cc84d0aed70508363f743975284285f07c9ea650f5346af3317922e8862f159deb57a5f4562be802bd36ae58fb70a11fc71be59d4cfa4cb20164a641da254227a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a5389c7654431022e91784f25ab570f5bbb575cb36ccdabc9122d6600922ed4f1f92c3d862e10fdcaace755ed632a6bdf1f0a89f964bea2f580868aff7c95d2958383ae6e552bd956634a0a1e385063ea1f1a626b85bda7da8316c235670d00f303577ee018128060494d1d517a58cc691a71829183b9b7ae556029ee39655c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9b8a90f622d02f33bbfce8fb437476ef421aa49b178d9d5f50ab02d5e28c927b781b921becad412536b37b3049f2724a94e19ea7490979ef78773bd6fcc937795116638d44b9900607c703a813aebe4fbc3ca76a5196baf0dda18648064faf4749d15a40a7027ed9cac727d394cb6bd53aff95da8cb94a193c454048fb7f29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac51de3163afc4b6e17c1bbcfbb2f6d7de2041cb4ad761ebf401b439529355055587b41ccbc6a5fcf6afb0189432a10c3eb673107967ac5f4fe359796a1f2f4b2b9d7ce2323edfffb950a0f53b58d3b34b4fa3e49b8f683a6323b797033c41c05cee25b856c736ad85e431df841be55ead96620b6930d332dd2d0ed98c995f4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h308d851a07817b00c14cd57e5616ab549ea71c8dc9e9f0fd2f5b980dcea464fa8ef93e976ea8cbe0ffd5e856dde34a67f923d1cd58a4bbd697343e5d915d8b8be7a346a1576a2b2d79397a780cb1ab3d29b8ea310f49d21164642e81482974032a6e1552fc302cf2b061ecbb2350c67b284944c58c36d490211733df66738292;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf222ac2b17be7dd69a5e60ecda59b8ae25795e486354c6e7fd9bad5bd5b3d4d9ded1b28a49fd22c0429f2374e73918072295ff36b7cba34545a3a4b9647300ab6d37c36b09fd1efffa4a4bf96250c3c4748abb088bd247e9794f4257f06f403123e8bc02b902db2395e0afdcf36bb4d26c2e1417601a313e59b263179749737d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h398e382880dbd940fe19c10f15d7ab051dca62d3cf573c21d76f4c696706639e7df18054592a62ae4498a39e422a18a5d4abe29ab41466aad8cedf12f6b18f34a1305d41c4d42c72785ee2e8e8bb9450123beef6927eb586025b24ec1ae689efac43a6de933737cb8002c5105074393a5570d1447efef0bfe0c142c91af50e0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1a852876f2f2098526d6a8249cca4eb9769b422a14e22f35252420a0605efe88c1d3a5afdee1639a3f8e3d63300f0f1747257b46889da7e52f5e79df4a894aac4c4de151e3d71936e1bbb5cd714c0a349273f2e28d6290f2a0f3b615427cf12f7f2c5ba1e3e0d42deb249f5e56a67f68e35ef954c2fdf6865e5b0bdce0b9d60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcff8f367ea6a953ab35b36f1ac73e3bfbeca03e0b4b65045b371b388303eebf462e64120d447b4d83fe9ebd4f8990cb495e95b64e5d8a47ded7fd02f83ffeca7a24ddfca2add359a3c5c1cb99c63ef6e43ce0d9fa023a1069d9dfe2e59bc64b515bf818f689133175a2eb208ce08dccfb75cffc218f9f2d1cef9228e5b3d06ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf753121aed4be55aa87508ce29cbcf5fff7e2eba32e2c3641d2ea74575d3ca94a2f9a782a9e8bff8fa28831a45cf85f3aa76d23e2551bae0ddff0b98d73a9a93017356fe6bd7adb0948cb74f29685d963cf5b006c4b40096aff1e2eeda120003d3729cdbf7e9e9c6d1da7d88b27d3bb0b4c08a2468a29c28571565978b8c686f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbec0f6d22ef5b371c7b2755c48f39db2fc3e4e46ad487debb6cb49e1748778a04656d235d4441dfd5d06682b518a1144f674ac83a25730f747b4bc3b7cc6d8087c97b19f558b9efb8516b1432090270737cca55d62506d6bec5e49ed4a1c3f2cf3e5a8965f48f1b540db8f071b34aa98d9fb22f305f1d96d1657a31db96c5c0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd1967c6e2f3a7b5b37dda5ffaf49d8ee957c71c4831dabc20f31344c7b0ccdfa75e15918015f1fc8610ee693bba84bbffc1b16aff66be4eb3cca284a760e35de04194d3235b9a47647012186083671ec41c3054f8078bffdb2aee9f99f08ae5e281e7874af71c6fc641b1b9595f33efb4eb8e24658156987f9ba15af4be13e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f08a5782783932ecb757755dc2f126f2ea4558043f44f5727fff3bb8a6bf108779957f200c218ea7190830448a07e51accd9c588784fc3dd0a56be638fcd41b058921c8583f1b707f0d5be0f1c4492f525b682667d7b92400815242721fa2ab98da1e24368564341f54bacd85c039ae51b7de2ff807f715466bc704c89e228;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3781398746b74f6c696aeefe80917c914597b53d03012c70e6d8a0ba35e126505d669f99d1ffd20d1fe4275bd8b5079750db2bd333ecf0918052e556b62cc518c7e9794959351f9bfcab84931b209be4d436a2d47215fdd0c3c90b525b4ea65e5afb372e37c7e95340dfa9dcc0e1f6b69d61aeec56a0c27d0b434bd2b80b5710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45cac9763e81c66ff631dd9dfb2939a5cad104f530c2aba588448495dc2a98302dccc4af5d9e9335293c9488630dda3d8d8ab214db3afa5f9a8d61cf4b7a502c76323848a0ee88edc4aad6288a1a7d2a6d12ad27f44c837197fb15fb3003a7ebb6f0d46e1075f40120f1b833e5414be9bf1e9ae36290a594093dbca7c924f8ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72897593b5232cb8f6ef15294ce638f61227733abadd16b7eea4a246a7a56c081f939557940adb1bb6d1b524c9913a2724f13f4aa264707d4eb81633dbf957b1ab1c7fe1cadd0ce74e22add14d88cb0a42040726f70223f031efc6bd7b82241752e1e146ab7661eb0f4dcd3be6fe2b93f40968832519f1da12c76ea301c3be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55d868c2e5d2dbd04ecffc95681676978c634ec3b9d3fc4befe01628a3941b4b60be9eee53620b08a64b8857bb3e3e777158502cf447307363341f935d2900bf1dc60f7c96b0c894416ce1466b1fa33089d403ea416177e3a523be6771a74709458a1774f5c94894c753cdd75f5a8bbc7301b43e1d362f94086799ba18c857b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h302b5ff7d364a3806a6c41794731c2b55931eba1d654caef4f97b3ed1856e8dd596f3b85df82e310a4277fcdebe838e1f783f9d7ce3f28772ccb4daa118791b697b3d96bc65b76160ed4552cd7e7ce33ce972e5f53072506c30f132ef8a1c670e1431b1c9fb7087165d7885bb119b1398e487c40ca9706c2a80f5f20a01a9714;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdd8c8bff264bdd815d601fa09b97fd68980f3cc5998c64471ab4d368b99c13993e89e673df907ca8aabc712a36298c3b74d89ac6cdd9c0613ea6d4ecc42c2f86d634ab646f21c805ec7b483fe511b1185e13ea4363109561cc18916b714ee99b2e586e45aa35eeb9b6abe6de8fee58921920671732a607eeab4e89b2c1a10ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e7222bd88248ee8fdfa914b5cdf8430d92a34d44c6ddfa8700d936b9362ba80f66d15efaec3a96e5a69a2edf0f2703bf6ce915399027a50e67e8d5da314bd4e33b62ea5f745860be23add43b9934137c2d6e3d9d9812b2cfc498054617f027b12f111136e7b75ab49b6bbfbe33789df7d80b438564a6a95baaa53ebe4d28a14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha88ba74e1dd8789b3afec8e4ea8f6122863146403d9aa010378e8d107d0cbf346d397b0eeb5337fb903602ec4bad0ea34dc4377fc8041ece01e9e4c263e451f146430de187deaebebd4e4aa04f4889d9f02e3b51e28f2be64bb60df76cfd9fa462b5adc96bc5994065c43f611e52749040c8c089747a7871ca93d51b7ab4e0b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b86a52fb34875eb41c3448f2c3c0b0efa6e9cbe989afcee2b95c953d0b883863c11159fe8a9aa305b10d02bcdceac62641b260c08d654e8d2ab7686c87d0258f6e626b7a7bf4fe36f0225b2392e0933c7b14c825e850721a23fb835a1ae9d290b0016516edc1a0491e6f90b602e8fc3f65417ba4119ca29271fa5cf4b3bce94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafb670e299b4a291fbee35deac476aec6a29b839cf548421fd5211cd49563bca7c4ca86a460484906350116f8a9c4c3cf0d0bb02c03d9646e8bb3b1299d65b0cf0d43cdea73178af3109b781a2db76d2238a64a3da1e2cece605247709bc13c0e3022fcb1157f6dc62600ce6f2a1c1a26060c3df16c132b6cc64fd8259c5783d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38f125ca34fa583907f06e95dcf7741952d84b6a7cc2f33e5194f54d84f72e66de63aef1abc3cffc73807276e311473e476bbf82d01d5d322b0f6a4a95c6ab26b10b49e168b8fbb0f1fe4fe4887ef0efff36317bdd0fc1752b75c0548f40d654d261b650f5f461de7607ea9890972bff0604f34144aead46b1a19c74f47dd47c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c64403ec4448e0b440ad7fa80f8e38d3ae39ded71d854bb5318f5d7ab774d230bec3926ae2388e625e280a6a0829f3e11c3eb805410fa04f313fda25c3bfcc7b868b25fcf4f1689ffa9c7cf78acbd30e2533a48d3300c1875d91c276eefcdb254467b9a772179dd080ce25bf2b7aafab54a1ec56df520c83a4d458971f37aea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h551acafc95415c6490538538c08e9e50d223c78ca0e0dadea804537e571d8693a922dd4890218298c0544b76a8b41517335454672c412ce61b8ea2e2fb03db0d537caa14cca7c0da9ab34a45409cd7d3eee30250174267216db3761c83272f2f09945061c3fc6ca7b7da9f0a34344bb588f976189c8254f698f9d53934207c68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h419f6178520a1f7442b09719441a02b3d81e564060b860d641af7dc9216c43525ee84454b12266f82d6af7be46861b69f154ec9dd0ea5b34bc47437f426ceb1d05a6b2339c4fcffc22a5423d42e6f36820ff4d65987006dfc91e1f17ce20b0734ede09e288a8f7c227e931c5e0c1a1d893348f8b7416f76b7461ddd89ecfb3e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48b42108e3bd57a3fc8e9e56c675d2e6195683ab6b075cc2873c5fa56620efbd2afba55c5de8283909cb0b26ed6289905ef5b23dc1d374c2d39e6c7677ba57ee90f51182e1d0cb99c6ce3abafb50f75bed428f413884f25ffc00e930692280f72b4d8563273b869c800ba2916f7eca4a8426a7e694d25af00091a02f18c3fb53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha39d3adeba396693d1c716f87167b149b5a4b3c6998609092b34b4d46fe8c64ced91ffadcd10374005ee2ab8fafdc675799834af6da007e30e09ee8d543186058d56002e392dd8d20d5f4bfff58e3c649881a284e39c65e4a9bc662355a3ea98df2871a63bc925d7ea78b142b9aa1632e153bedeff5b5c9726107f496c55262c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8b85aa2bedeb82bd09720915c62a8e4558a3ac1f8efe861f8e5c498c84ef59213c8dfc8187690e4fa295cb76493eb39c0da5456e62698afe872292e414dad930cc945b80a751d26ef64e872bfa970895ac0caff1a1823666e56dfa1aa8103a343909f5b43fc176a8e50ef31572d7dbbe2a71c89e9f98e5dbbb1b44549fc6278;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c67427d9cb6a90dea916a2e85ecefd678c1c191b65ddb39a560c7a8d1ded37aaadf850647591152991ff4fa3bde6050e4b8293c9179a6da3c94da341b085e99ccd6acd9e520f64b37df6d9b9001863d5a3260c8e9880ae147662090e962207fe5234cc6fd4e52916a9455054a8fe8827b64bd87c02da4e8cb9c2188e54339b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40a1ce4aead6301960f721dc8f461c7e923e27407e858f2e196d2efd5f8cac155be9873b94d0b7556a1c3dd8f4732d3973d1c620699ea438902b3f1505a3d92af43656fc37629d970ea0052725aef8e818fdb441fc2cabc07021753a29e92ac253b2b44920242225c25993e5ac142cec5c501b1f4a85885a3de5060db8b62bcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f2e27784c0d0d17f9be9946fd17338dd14993abe612c118446ba53a3a5bca6f9b8678b0409bf711b722b69dc02594d6554926d14d2adbe4300f9ed08676bdfa71a19e977c48af6350ef30e4fb99b55dd28bd8d5f0a8a1c749f51c58f52dbd8c6c6f5b115d55fe8eaa78e18f3c7ec58852d2ceff9a17e6e9a86992e1d5262967;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4a906801a343129519e0f2575a16350acd7b69df623e226915ecdd6d17c0f705f0932d2cb2925d833f021c214c46d40a770d5fa0052d5c127006f87f21e66d9ec944fc0a2d94d3486e94d6e352165092d5763be3122984150ab53bf6194c85bd91cc585ec5c664c68a79d66587901abb3622cf0d42d4d3937a640c3051704a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h531e7413dd03aea44c084ce160d76a1bcd48efe8e8931b7d835876a93e22642d371fa558b76744d8638e9f63b9620790b93bc04d0b6c4bb0926a406cfcafd855f9b3e8141aca41a98782b200d463bf1e2255c9c6958a61bf2f5a50064c4f2fc527b1d216f2fde141881c0614903330d7066b42f5f1e9ab9ef229577ff03d34c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha691e1678e1eda25db592cd0c1a310e3687f373c32ee28ac996acf4b11ede221939926de36eaddeed56fc8a79e9a91a424cd817efff0c4f908d998968d71ab3f5622dec889c096d92b44125e8efaec50444b4302b46fe720e0860025caf726b29c7557398b5527a38e1be1b45bdd4dc789e5e9fb95e264f73e7e82c9f732aca1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ffba8e479947b9075e5586f03fddc7b0fd9607d6d7a218cff7eed972f441a77817d7d17858f771a2b94cfa2a5104ec9853e45945b812682bf2a3a8125daaabc327a7dd5c03a2b191a1beafb3125d6595017a4591f9d65f7cdcc4bcfe33cacc59732f8140e8008138cb0c64c17acef2baa5603b0cf0acaa233e535a93080fc8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd597327c2b02ab1fd64ddf069ae4365f4cb61aacf6b168fb66d324204e62228bbc95077b14808a3b56919910f969dc87769222488254a16d018589ff97c34252e25ac839db2b27be2f30291becfd00fa41d4689b1bc67686687396872222d64bfdeff9d747da7a80cd5dd876088499248847937fb7d5e2bf9348a5460bcb3b08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaf5de92d45707e22dbf9d5623b57ea9bdadb051a6754394e8aacc6b0b090b979d32ab17742b8b46a1a2177231cbc61946f2a066d6ce5baab388389811ddeee75f70b0662f968337d1b275ce4507845e0edf4ea3b62f1db6e19ed7ede09737006eff1cbdb0d6067c8b19f4b23ba5a748dcad720515d8fb95b92e4569148c1137;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc5751de804a3ccea79c8a716b18d9dd9578fd3118da9d871632774d0b7899cf03daa14c5447afc150431082aa06f80bb3d5b99da617b59e97971f0b84a1d1cd36e373ae4e2b76f98920cd12500adff93d413da4bf515b756e62d736759549de452351cd71cf7565aee432dc40739314ddd4559bdf415e923c1d4e0f404a5cb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab4b4bd5a1f514784201ab9a76188d52bad259b82619291788918cfcdcf1b552bdb0b533236fc7717a775845764efa92034ddaa97209909bf284f534ebcac183e2ebd73bdc796d2afcea21e3207c1330142598db45a9ef1206a27a624f749c12e11a7eb35e4229a69d2149bc6f7d46e44f6aef409dba65836ee1153e28484c72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea8e16f1082ecc176c94b643d0e11a47016f789ad366d55d4d1446af5684c64ff5a96ac1d3255814c49c616a2927240928a96c567cf50a6cc020a469bd806a5b923d21973010aa857d16f84fec7bbdf069095e7e91c49bbf7246baee55d99a3bf27eff9c3a49dc8f160f730256ff5915671686855256889abe9e42b738f65475;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab928f8aded40a471299528dddec225411c0d4a42631a1222500c2f53450154674df259d271ab118d1835c108d4738c222db1f7511be3361e9b8e16a74d7e9cd36eab0e9186b8841a679e6658217d2f86e175f80a86ca588f05301c93aa5b2a135576a639a830e1cb4bdaa417f62e16709100b48020cb9e2d871afb800487ce3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfb934a6c679aac118d9a176e684f9400d4d340ea914b6d5a96310cc84223ba98f8e5b6c509f05c27b5c92f6af8a45650fda169dd9200f772045378beb486e9693de2e54f7fe6680cbe415c605c83d74afd6c875900226b3cb3f9b4c4a1c03050974361bd3fa815bffdf62d080c0333dcc381e2dbbefa0a567365931c60971b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h808a93b90d28374a7566a4f5848770a7322478db1ed4442a496c5f500c217677e04fba89a754eb2a943850963756bdb1969f9f753078fddca26514e1985933334f8e8ac3c441e0dc1454e25261f64a22d3769674203b09059b259b7565178eea43ebe9f54791a7bae21c8f329442a0084f53269d2c3bc235a061e5fc4a93f127;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd84e43d8747f399b2e461a89a6673926bdfe9e5bb2e7a54e31e81518f43dc805b2afcc330b5313e04070a83b96c40e048167bec0eac9f49146b7a1fc74d24b98043a0cb5646a1c3fad5ced3963604d96858e39de70d8014f7924e4291baed947ea63332382d1e9e2943ed264153bf4235c84c0a924ec713baee4a6cd3a88cd34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e102169670012ee193c4e9479c268f76429c8eaf6c1af4065f4831c08c50561a4ae309635e516aad2d48c353cc1dc583ddf68b0b6ae3682e6f955964689819d96dea7fdd46fa6f11f0994b2d50c5205fed2a054551152215a9e686b7a3b315dc68450dae1d2f77edda444701433d17a99d193ec3a3ee8d560feaaf3233a556;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h448d15ade22ea7387ad83aedd122ef6142584cd17081b7495dab7e3b7c47b22e6a4fa94be8c4faea9f5fbd929ed00b3068e8f5280c4979efeee19485f0bf5fc4c3738ffeb6a07fb5aa11dc6f911bc4eca46fde32ed7ddafd1b542aa9f103a8ab4b98071c1139ce767f4cfc226951b6d7ea6bb538877f079f5b979069c5b11ecd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haff4acbc127928962d375a569f29f9e80d82a19d4ae4118a61b42a8ce26921f1d64080c33afdee48a1b6bd8ba8ef0f954c0010dbed33ac3095a0a1402c5a160e8a6dae62d501c95ddd76711b0227bf4ee71f16ca80356f69312053090d48ce90ca38d4c3a1c8d501e21de9b317b21e6ae71b3fc7ea79ababecb92122f32b7c3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacdc86a5c2361db2bdfa759ddaef62f7334f78fd328ab8bde224e0ce1e608ddb751c7a1e0c0ae4c4da995035797c2b4a01ace19eaf92aa297c7867131855eb45941a0b7e5ac5bd9412652e58d12461a1dab0153e0799627001579806f49580ea9e1326be9de6f7c0eaad940c6d84a84271c2adbe70b6bcdde7d6778d7c92533f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc49f1b4c0938ecbf6ebae0ff4e13a46f6b81217c4ca87b76456f61776179453a973d6936cc7548ed00752a6ae3efe67d6826dae2525fe102b2aa24de5110eead48af83a65d063e540220d4916c042d30bae4dfc8bdf8b4c61ebc1b3a4337f80e7c02cfccf9a37a95a320a7236e30d7a17d15af6086173829bce146a6dc085607;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80f9982f6301bc2629e4603034bd0a812ae8cff6bf0d57040930ab6ebe7dc4cb2d441ea793baf36cb1dcc88f1a7423d351693b8e6dffae8bd7d53fa5a84f1f028dd0750cb72d24f296c2e87568830280c16988cff0f454112fe5ce06eec2c06cfa75816e0888c8b3f7140ba75efe6e03fc7e7095633b9be6b6725529bef1f3d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb654bf6eddca398541ad8c0540d0197ea263211e4de63fabeef6b0e1932868bbe74bada5549d1f4cf9969c995653a6aa631aa17366074f8482686a2f1d2d4f77d04155d997abe2c1234a5710d164d8814d47a817b167ae4683e2233968cb4e1c810198592d63d476b2410fef2e09aa210bb0beca9a3f26f66dc50047edd8fad7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80b5274b38dec9eb94e1f9ee0a057f77c9fad312857232babd375fe1df2920320114a42d5b65d391ef77fb8013b4569d7f729bc18e1aadde58b0743222d574bb36e8cf38d0e3a9ac590244e51811cb15fe9ff6cdd191b45e9775f90e8abb0d7caeae3e0f83eb099e101dc1eb0b5cb86f3e6212692b4bb15a0f592be060699113;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h822bbbe4cae026d4ba4c72bc3d831089e01061dc4058d6b6f5ded5d34a55579ff3834fa7c2d0a4f797eece1b2c3e0bf4d7ac67e09a0e2bc15f373582162f0bdc2b6c71a94de76099aa0a8588df1fe902f9ec1e0c106c457ae1ec1f38c3d38d4866b3a7e0908bd951bdb676b3198b1b02c24f7e6076e407b8f591173199449e3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8624d080472fff951ffc97bfd1d3ce993eb9d68a03d0488808d93ed3ef8157833d392b0f55e65eb3f3b324fdeba13c50f95adc3bacc4d4573cb3d4607151e457c052f6b37ff26efd89af3b45bba32b32caa972cea5db11c997888cc13218cd2d8d8923e7921ad6af0f732af2603c442668d7fc59da2197a823540b0251be1624;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2332f7dab96e4e0c882382782e54f861acd30e4ba08cef1c9f9a5417bee059e35074b9f1b979789f0569197be1259703e21bd30245ff70771d9738b94351abd8822ca7e51d5963f907b4b489e122ea8e6d6688919283d47ffe72eabbff27d956bc9b2aaf5201834f0f239ec4627fd143046dd3922968764a25048c3cd12ab3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1e7bae36eae5790cac56c74b1868f1bc26a2b792c36773512d230b69a4ad4bcdffbb3c93614ff5e7e4d7e89fd34dd2433ffc3ddbfa5c816b0f11704f4e20f1a654b076f3b7ed8784e4f901801c19fd16504316d9752568e0ef1c82f1f9173ac006f042e9624980c01e071453e32db716931fbfc52a9496ba55a4b91ab9ab12a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9e23e053a0facd036a1a54828bc486a0947b33a5763d7ac9f61a0bf98255168b72e1fd4e37c95414ca3fd748d517486d93f7053d924a88b75177e696d4f625705adb4054aa903981e45414e03f894eafdc5065ccc0ee1d93b190e73f7eaea422a559c4561610dc11dbe1c1aec5ff09db927272ba4fec20b92f29644870c8399;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f2023326f94417d5c115d7c692a84065d6f86fd9d2a72a834fa7cea14ccb34394655bb1abf4f131bfdae14bbc827ad53057c200957bf0b1fbb8cc1bb2cae8f90224d4fcb1f92c4629447437cb28d3b98ea2d6e3435d371eaca14bed19fe6eade44ff864a53d49f64f6226df612a6051a055d7c63f0386b2eaf9d5fe1e045103;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f1e58c5f2f4e30831db9c6e6a749fd686e3e45bafec95d7fbfb3c710c880550e068eaa8b157d924b524b0af91e4d15206eef327dc9ec29f393dcb7bd6a3d4b094572d49dfb0e0c770ae898557bbcc6e1f0cf405b4b710b8880d06707a991f00f2103742a7bf01b0a9583c4ebad8a0d7f373a4c4a58d7a28712ee66e5c020a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42835cd8088b74992d7c1678d017c7f23e77aa15471a0de4765abc9efe75feed00b049891bb730fe49d0f14c878aa1314d114e2e0dffba5062598b7856fa59e623fc36563501f941195aa909fb42f7a9117b38b64abd7257b4eef0e104717719079b3c334873345318f7d8cb6c34fd5da54a33add0059ea68cfbf2370d648785;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he862f458c69404a7d9449af602e344f03d5ddb866898ba360036287ebcb7d8e41a9b8fc3082a451de36717b2c2c8df12e9290d433f04be9284bd9da024516eaa83ea5126597bb5caa870c80064ae3b0f1908a51b6294907fd469e63fe5d82b342b75a3e9bf145c64d0b3c82ecb4fc9a692c61a06b61a926cf2a39424da28bcb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he46e1b017f61fd66aeb1d56242c68453ea42423b51b6debfc3111853654a5f72a1ccc2abf8923f56b3e8b6717abf651852210872f8ed8a27380bc286cf3bcf6e06d81fb2a58099b3d226e29abdfa2366d44f9180700b841325b97fb2d06010879be7fed0785e61f372a7bc4f0202dbfb6698dae14c744d9980dad4ca64199959;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e44034eb0cd618d279cb094bb98465fa62df2534f8650f235680c4aa76547ec9de5b13d924bb719d95787fc20002731c655e21d903e42b60228535082b0cc835e433d5dd0f35575128dae70b4a252c39830cc864f86b02ce27d6e476642fd9c0f9f5466c43c8e0be97e891ef8b915eb80be3b5355fb67b65eed4b47ea904cc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dfe95c5e6a4d6ff3373aaa8e70193df1c483b886d9bc3b9c096108f9587bb4fa75bddb74cfde6b6e3155a57a8b3b70cb0777f276a0745c881e61d608e54c6ef7de5a8be775dd4b8121fe6260d6beaf11624e8b47c6f57e1a0726c005f2a4172eab1e83fbef26c2e1b0d76faf12e903652dc405dfce9b82c2f44516e9e5d540a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd77621002cde25c265f7f461f407dde081dcba9c98dd99122389a3500671f94e72ce0338b5c6f3dafc94e8f4497c5748c4b8bd76cf4d3e0fa92ce31ce433f9d32320775f71eefa501caa8cc19b6a828267895a954effcbdc6d7c115d095e10dda694d258d1aadbaf7d8ea08b2e6dd86822d65d964fcdac76bc7c154ec51f8a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ae1926264d5709ccbdda70014f19b482ca426516f8138f592c542c1451e8958047e9309518dc7d1ac7ef900516e54fe463f96202e1a28991ce7f950ef848ca341212b124cd0e3d661acdb886ed947e7edeaedce8f190a2430856dedff18d4a945f31b60d78e1ed03563fa59c8a9b087c1ee0001fbd46d6ab56e4d62f3183ed6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h924a161d0edf112ba7966de74d2257904a5a6dcd790644d41631883bc29c7bb08bbbe67814c964acc21301d0f76ed8e41e86a9bfe5b5a0774cc3b1be61c4333c54d98411aae7215f65b26ca71340859ea5b0dca752eb36f603d15e5351cd84a07de288e412a49b8bc75963112af8e6dfd8e9f9690a149a0b697bfc361061d379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5470e10c84de6af9295830fd66cd61fed16da036102af387e507e12853067692702bb6bff33f75e659c536465125789b69aa670cb3066677b3e47f59d40e90f210bd459b5367b5dd22e258e532fd7d53546a1df6152f03254cabd7c1e81a48c9ed67e50cb06a2d45ebfb1a220eb11af5984de41b6cb70543231673f8429027;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85b35763f32a612be6a266236c70573a3e2afc8511a0407b4af5c8c80fb66206e451a3e8dc53c0c0066e9b73958b6ef347565735f4500e80f30fe0ddca43490d109d7415db595dbcb495bdae6637490b09b3d800329ae35c917754afbb179cb394719d0c50a90a1434422540c33477a0859a68d28a7450edbf3397374c18f385;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7576aa9f9d12db2cf433f84c8e79f8caf24a53a069113d13658be25f0fef920a5a49b9a37d53af14772e17877eeb836a70dd2220a81b620644e607c743adf9f127b1fd32a57fcfeec391693fd144c4c54554c8c629df353a6be4678b6084455c5549d11528eb68dc5fafdd69cc57875733461edaf00f964ede3bdad848ead18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fa9bf5e6572fcef45374fcb4a32a96cea9c03a719c3d4d9e54b9f97b7b8c3a052a4d367bcb21850302e53a37ab8f5053b24856ed59bb010a490499e8841c32ae231cdde720c5e39195277d78d2cb93f60b5d245ab12a98e9f604fc2f6457b7dd9ce451d98607072300376c687cae4e8d5ab674203c5442a7fcfa1779cb7a9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdadda696cf79fbfe4d9244b23c6d3c5e45bf0d40fcdcfeb8521a01a32ffeddc3716c0ab8d9a1e9a4149dc8f6cbc05a73172957f2ac53147b1a79facd12fff28b4f2fdf541bf9877210c8a3bdc059b56767072d56722f9efab6cdbb9f7857a5a527398a48fedf792613348786c9275a14ba897dc7a569b2c9e380499b6085fe61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8c0bca8414cdfdd759699623d127287c38c85486474cc2fe53507bd9ad213724e0d93e7bb07fecadf27baba80d498fb0355bf3175a3c552c0ad9e0fa73a4c371c4eff0977a75128a7adc555e73bec2e4edcdc4523bdb9355989db165982012389cc298cb084d2ec178d24d9ac17e7bdb152a38ee5220af8c289b386837fd499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86bba3312a5b7b51be419e8bcf82c37ea05ba8521d1afcda237400df354e069374c0ad6158f8ccee62bc1227f25417c41941b90c0e83ef22864cfb8278fec8c72f3dc7ca5b7f189fcd2fed33861f65ba00e12f046f8957b5802d9cd4b1a18bc4562d04e98449cc56408fbc08c5f419f328fecbacc5a5f7f561cdd6ec120980dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0f5813502409c049cdd86511c4ed609c8dd0439b2013aa34812c5db8ef7cfafd209db3126fe0ea7cc02fdedba3fb6a977c4750227c956b8b0619026d7c0623c18b63714722d78066ae98179a55180260c08ce01ae47e2b00ce7a5459540d5b53ddf9b70dd960a707b8c8d7ebf7b40e1589ff9d4f5f57af0f35e7ad37bf063ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h307a5ecb7254fbf4742faade329115c0f24fe879822fb885a612dc4f2acae0c75a8453a8a673e99d60b9064eb49ca08bc004470c92ee147054018ef5679a6b5ffa048147e23168e38bf8eee5f6fd89891f8fadad9eb2224c436c1e309f88ac27594e53e8e76143a60d15ba5b337c3f139f57af8cec8df8e180d12c0b2f18bea6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc8ace742bfeb536a21571228d719d3242d90277297128add2f7a9ca27728b6b8c375ca0c77cb23fd63b5306b9cdb07f0b4560de162ac3c6ecb78cc74644381cfc183a4eaa22ac45b577b906c9965ade6e7d657d40ffa6fb3a7ce0b054622e585b16bdcee412fa2f34b07b9350061155027629b7c831e7b41d5647a1c32abb75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h806e21c99095c9e72257912c9c85cbacd4b78cf744a2fdd7aba1e514f6b191c24b3caaf86da0ac2487a6cbf3ad15c21ab8543f6c44a749649783d08beccd6bd973191b2910f325f15fa81ed0dae40d3b7a502f6284e09c3b1a1b11eb35410013b953c1edf58a3087eec74f8d70dc8ae106674e27c262682b92045c478ac0bb4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58ae2a9a54af61ac4f9ff9b0607b4d1f171a049c84092126d8096618dc42b268311656057df7659900fecb7e945e57d2aea2ba7275d9a9a48ce19e840b5ba44ea47a49ccf8f30d9bbac33a9f43c5dbfc710b22a985d8f16edfb96639bfb9b10f67062bb95c3fe798042df024ce833f57c0adbf3ba910a85c9d032729b30c47ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h227b38b35ac96b0e781f559f934f5fc336c9dd6ecb4e16a14ecb86c94e5e761f52d99ce1ff9d0c9f643e697bafc3c7a63655059212fe38943943b9c87238d74e66f0935828f0a4be7130acf71a5eb1d73178648c0ac26042214650724828dfb4af7fb9d471d9dff882d4d5aa0e227347975d27182748f26eee52f461135ae7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h848370c39c7d2972546ee21b2ba6e77c72c5defa904e1140eb51dcad4a9972e31450eeee005495b0ae7efeb6a950608c1e7f59958d236dd957f3d1fa27a25a4d20944d9a1426ac4f26158ba57c51a6904f455097915a7cd15cbefff7c2e9a5f0a32ecfc26d5a5f6a45013607a94869d4b18c03796f56f53dc93d6e23ee6b58dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21a02a5d53b54348dd6cc3d114e47ed3ca36cab34be45a14a9c37c6a30e0d1bfa3012df1e40321ea19f152e796c800635f4221f8f41acbc3a69ac7a3e1fdfe1bd22d2fffbb524cc7f3761d606fa8ea0e65cfbee34bc6b6763b7d3c85acd0ba2e4d74f7282b5b4925327743ac66e7e8c7e350da9d3928597f2d98049cdb95da9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cc789f123952a1f9fcf46058545a5f7f415c71b0c4b40effe42e27f546ca9022a9e40c18316fb75fdb4bc4a05635df6cb1f12359baddb0df61c621916c26ac6cf991c52ebd307179775ff42fa705bf891ed4044bfd162a2ca4a7410d67e76259b3ed439cc65c2ac6d88a51c1503170a4df8e6de6c672d16e71c860be6a9a92c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h472dcc6da06c8fbef38d1cb3715855d7389cb6a7867724009df45ed7e572d432912a34f4ae2d06161f88cbbe22ccf5c5b38d509457c54014afb7bcbdc205558ffeebee3f3e239cf53c638eed59d370cdefcd502f82e0cd40991033e024d5b26379f64cd5de24c0b7706aeb7708b9568f03e25ca558b5f2ae14736e1d94c70e51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28b79c04a86a8703e471aa6b86b14f4f34ce43c3b87e25456643fb8d7f4c918e7d2a488b34d7171c5dcf86a58016210f17ba5cd8039c774a4839a8dc495d997b28ebce03eefcf4701c0261514a101d57241c441ef883bf7a77853afe3dfe855f07894ed3c9e404f2e72b66642fc4195845d5595c656c9f77e87b98844ace36b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b978a2e657ca245a63e190ea9c8130dae2f9119acee873c5cd645c5dd64a027ec6a160d0c58a607ecdfebaa5bb3aa6b61ae932fe27b86af58691584eb2ffe4442e980cb8a0778664697e135446c94ac6d2cb39377e929141f3a42155937d278def723b8ddf1b4f60bd48d281483e4b42a17aeaa0a09530c4ceb30a231a01d79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcda24392e4f5abebd50b38d67676541d2a9c5e18954cc8dd0f41dc86b62dbbbb59aac59579ef9513429842cd286a98e2c6c38d5d160157de1039b776a698d3ae21cefc321786dc9eea464d88c8682c9b7161fc6967565098ab2678a33b8b9421b2c669c7a5c0790f7ce47c444bb95004dac240a8b0052d9ee19cce7036d63114;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76c8de92d7fdfa5892c0ad6d0f23f7648af4aff4c82cfd2e3485e81cccd69acbb990a689867f79680ef600d198da48a5e21070ff0030d806945d8ad633284684e3a5ba17b87282fce919b25435cd18055b5c1fb6a62f117af1b15f361528b876268c170e4c71e52d3da2281c2005e1ba72d4466de1c60bf847bf712ec1bd808d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6275520e0b6b63b43504e50832c275ad0bfca4477138962e990326e0ec7fa2cbb2478eb3c7496b125ef03f44b7812db2a9e36340affccb4320fc972d616d79df836f430831e3087c053219e4bc5a7fe155af5e3be21843a4c5b7424ed02db1e04e2d14d4b6fce2441b509134a9b4dda90141973cb9257bfefa7bfb48db93f57a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc77f9079e075b4d1207c2e561f446ad4ec60dc2f73d0d814d0f8e96936fcc69890a0cf0a5f0664dbaf5fea05963a182449321b2bcf5ab2a6948c9578bb996ac84c4f9871a37aaa6361b53adc8cb6266419cbad2f774faf84372e5fc34d75fd94208b4ac19840b24b16f2e51270b2acfed5f892b027f97b6a47f02ee9039abc8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha73e436e6379ec0c84d8cbe61ca2f4b5ea5a1328993ccff2cab6050890b62db59a8a7620a84af5a6dbd2798e15958477c2d833ab2104335dc838e25df4eacc52d3e40bcf424071afb1a79b7b666b30e3887477f29c5b60531d24fcf360fded1771468ee34fac67fce9f18d852c0501f9ca1768ebd3d359792886671a1f0cce24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92eb39a4df753537e3819ce5bb80b3a79eee32ef424b35fe49651268e44ec870e6a2cc06750d36effcfb1666bd2fa46b998c072f9088129f7e002ad44389c6ab09127bb11e8c2693456b1667e247eb8b7c2eaaeaa841a69db14878c06a26b252f1414b48d64e79cc25d7941729d58d6d97737543d60a25ed7106d8e4aca6d306;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb13fa97816d31a8de08b76348c8925b14d59bc4ac37833602e4bb889e2f27d72baf6e6e914e6b40c260bd334bb61f73ee594dbb117c650af00ebe2bcb10c3464fb19f59209a39e05d3c98824f2cc8f1ee7a71e20bbcb1f315f20a7167d559695d6ebef841d413387a75f5ccab0a68fa7cc938d0d1aaf24df4ae4537744785ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdbf124916fbcad1e3409a6d56e725cb637aa556e46217a67a3aaedd6b40bd64dea0d3d826ab8118a2741af8c21ddfc224582eb8e1112e26ea7de13e8d35b5f7f9773be5e7ab894369e5d7709cd02e4655275264e1e826f3c88ed2dd54c5ae25d33a7ed422b9f476783c145616bcdc11b67ce5b78f8cced2d16727081989322;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f00e5dfecf0eda2af54b13080c8ef5d1aada66eaaf2b4e91cfb221af1675b3a2d0cdf92d36ca08bb262d0462d5056018d5638bd23d9d6fa378497897f4929791ab1f3949bacfa4a0004c379f3bf5ffdc60bc3d543ad4c42dad60e61f72d79e68d2ace8c0c1807c2f98d09bd7abc087c3bfdcafd7a00091b95400b223b77fbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h864237d65ca10423cc4cb62bf0af614c167d116dd6a52e4ead3e974ae1a41118972fc95634588af0f8aa2b634e06219493d77759cb1d2fa3669608ba35aa8c807d6ffffcc6942109f341edcb74cf28fdb452a0992de34bb295332b7059a31f201ba6d36450c43b4b172127776d8fa9ab8dabff30ddeeda61cb3abd02f78efa78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h582c48150d71da490c8185dce52b99075d978b533b97b9abcb0f66cc23380f21ba7d2adf19b2ecf5720c317524a4216dcc0f1842d20144e737a51d9318ba87bbb064300136ddd93999a28f3fdc3f64727055d4970473776ba5d5eca47913cc719927b46afcd5488c3c807a035b1fcd4606cac5380c1f2edc16a8be56a41beb49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac47f973fcac86a7132c229f14e59ed86fb404ff7892cd8380493bf09afc977f0da57e20b4f311a6301c9e627efe39421c7badf6a6cb954f391d6ee4153be125516708af04e91ad3daf0c49b937f23b82ff5e03b01dd8116a1a21bf9a1cb73bc07377186bb8b99f063baabd77526887e5d2d56daa9d8159885924c8b84c16964;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95ca93c7cc4862cd8949a789ad5b1c8bebbc9707a43c241825550c9f477511acda48a7c2218691fdb569c6110d29319f1a8cef3629278325aaffd447b759a4aaacbaa60c9bced24d41607af71c6b61b21b7f0dec7f5d945672235ceb677c2b1cf0b693e960f379ae08216d9d8f2c69bc5d0e82b9e4e9b24b0e20eb051eef2d7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89a6a5cc142707b6b933c18f98eb3305088b57d4cfd7a4277b1bb40959a8ef7d6cbf7fb830d624a408a9998cb1888e44dad2c68301ba46fa6a47b878a933725d279d5548932e2dc36c83de7d1aba46b21e103b45d496b96817d6ac1621622377eaaf9b3c26d1a33e4b8f02d86f60371f7fb2576a57df527c07fc4e0d2ad10079;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4e8f69ca005450c1524d79070e7e9f93942a8297f7dbe754cad9ca85870a8660d9563232dfef7d2d7c28dfc75994ec1bea90f155c9ba57caab7668ae91b15e96e432d2d8bf983948205bc337a431c2c939d22909af29cb1ec5538decf522d5ca00bc6aa42210becdb39e646fd4becc86350d724796a224db8bc21b3c3bed8f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d4ddd0e3b2def6a3d51256149525d534f85d38cd78e6f2c519d171837f1331498fcef7de97f73f3fc0d0d8fc066869800c5af728bd7d0f3bd0e7b85ff023d492ce08ca7b2c81c0c1981eae8fd042cc4472cf164a03f977350a6e8ad6ac8fff9e86d64e13ec21b8a7c00650c6d1321b2ba9ffba70dfde662f7905e96b4904647;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb39bf7b67a80185dcf792e5d87dd012f0562b68abc511e44b4198b9dabd57bbf5273d46025be33c4595313fd755d5236e7747af53203dd215dc22330cd66b5a213598b2ffd0468db7d404aa4bdd0d6411d2c9ea5edae8d5cf5431394a9ad25795e71ff427d8970ae54fd00132a03410375860090410c5cabb6aa2ec2a53edae0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b9660b689d4970c7403c9285d0baf07b3c17bbcc76232170e3fb47ca1bf452488efa4f554327a033ec841ec9e3a4bb732d1db21a228961b4fdb8645a3ace98222f76adcec01387ed2e8df479c6cb2022fdd490b0905b7638381265276cda9fbe3b23c13ff6daf1817231fa444a5bf482cdab6b0ba22f4e46a0c5e196d711a87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h954268addb9c044f507d77de4f5d0196d9b3096c62745e55fc0d69be4602d5a1558f3a1dce742142c8648483d069a9c24655dda223e9b2555166142c99631a276a5b5a0c1ee1e94a72ab2ba09cf3f209e7caf7ada84e28b868407ea8de4787670b7c853d106b3d51b78a46b6848c0ef2c5cbe51bf05f8f84bc6bd27f361e3f9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb357d388ac6b26c101311cca173e357a6de26cf1e000c8102c431a61d61ec75c950b45128b6ec94c9ad746b47f5b3ee73e810d87ce6e45038b340d657a5df662394ddfc30f84f436746f1698124cad950b25e7211c13eba83a9e3269602b7a5473bff2d9c5098256209c3569caf86fbab46320b5510b542abc14bad73c2b3fb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he863c3748dc8758e3c86436cd9c116c0d53b7f031edcf1c9d720f4409b31fc79e4015f26e89658061f87561603543f8c7ec46456faeb866391570103dbdc110a2b027906fda0d067a83adb5276e4c8d2d11f2680cd426dab13ed0094a70d9090488b2230f11e68cfa6109dcdd0f5c05c209cac711dcf4565a2b0681c84022fb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7929babdc728ec51c16507ee8ef230e95bb3b22f0812ae725987f2ddc62bb488ced607d4431d6804b2de8dc57736907be70d07d7c846fd1c39209ac63eca2aff6e8de498efbf5f500a32a4eca5bfc48431835098a8b28e3f94a4f829e41475e4e67ddb3b15636e545565b8cff7f426c65cf949347085b9fb9712c3ecc3d98f57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2fc0729ecd39fac6d69c2066ec2d4ab109cb61c82944e8eb5bf6599c4ee17558b000b125d56dbba37dc05c4eef7a5aba92e425cf6a48b33071ddc26b8af6398c6c01867a43fc71a84f0b5f4e1b30199e767734fd5ce1046198d100270fec8bd753dc29828b28e7c3f2908930afca35a7c88ac582aa21136eb15d689730e4bdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3822ff2ca82973dfbf3526a5cf074f29613fe216f2e2bd68da239c4714eb956c0e1d9f1b898fe25fd820e297e70c5a724dba78223768cceb777e8e7f81ec4410eb939b4998493c79ecab08bdfb7c0a4219ebf4527da2b9551764f0d66224afd9203904261cd4c2f92e345feb2b247dc9c7b948472203095826afd41ad018456;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf32f404105110b631ca2fc0e14091c14423fb95f37a668e2fc4565b5b107ac1e9cc78fcd50b951b62583c4ea277efee0a8da2a76f89e5e7bee7ef7e2a6122a7be982765cf8c3dcf750d14e1010eb2073a52f0536fba66f89cef8439a281caf6e5a4433fea79dda03367c8fddb6106300b1ba887e6759a10e4be15621d6828e60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9613073d07076a6e37c5ae066256ece3836926d420174e7517125ccf33d5a8ac333d015eb07e618397bba47f4f5feb18d17ed8d434bbfd04609043504dd556328e94021f84b29cfab5744b19389d24f279085192a53051892b10732867ccd77b6d52034aad07cb956f8a832c83d57313885277bd6bcb9ce1a6b730fb678d9af2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18fb7ff9c9333d138072107369724f5b05ef9ecc46d42027b3826376373498b1573defb94603e4f696df5e1581b86ecced86d66e6f23c97c7985cade65682f6227d918993c7f46a96e6ce706d8e0a4f6e494c76d953537b15079ea575a5fbd01aa04a18bc79c18dca11ef1331ce41a87dbf3dc9e9387e365f3ef3c4c12b63ad9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eee1688f312c73bf698ac8f4c6f41b960aa661e7d0f1bc1290d4324c364b8e3eb7ca90fee5b1344d399009eb3ba09052da6f38a28012ee21976559bcf7f631439f76da1d680aaea00d7882b755e4403a83145114576e94a88ea0eee2627f7bf370998e37f34dea60bb6d0156ed7b2cea1c42b3391d700076e78f5947d43581f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha892b91f615f192cab945d7c0fba3520ac4862b855e77a750f42c5e95cf9ba2e200722becddba128003b9771dd040208abb110ab18fa81f315c5e97c5dd2e1d96a48c3857e4dde31dbeb0771bb1087381a346438f3e3573c065a701641f9bb076c84ac169df349d3566218412286946fc5f57379a26fe643e7fd8c1fb07ef9a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdede0990bf7edda9203d1e0048a62ced2413a5e889424993310becd3938d25fa2730c6c633a76fabc46e4406478513555c0e8bd26dc8add7b58e3fda200cc1bf844c8827b351f3157ac63243894d5258563c0a05598e5537442c38466a3de6b8868a06af72c992cf07b97e17c9ce1230039ac502742f868640333b02e4762c30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ccbc0eea90789d666c9645863c1d47e5488683c39d4b7f7242e053fb464cc7530b7a4ee0c233970bbaf83181e0ece77ad2c82f24d166ed2935835074e6e178c36f89cafc920dd2e5e38332e26e4a5c4a53e843d622d8b762da1a82d0fd83c20a00d386e61babffd27a45fe2420c7aa4b4e51af525ae7535a4102ba407ba3d8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1567f03fa49ab8c33a5dc36373c761165a0eab934e1faf8d4ab5a4592d053e4094b3023fbc83e69277ade027930ee764b4001300963934782ea054e82bbe6353f42acf90e49adc153da101da342401195962bea278fcc801c11e55f9480fb75ab567e94f9d8ccf2eff747b7e1e48e2c81340f2ca3c7e458c4651ffe1cfbc2c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0c0e9d2e50e2f8027bc787b1993798b27043ff85caae01d731fd2f020a2e8e252e5fd870fef73225f72481e14d077dad2f17e6a3ca3e2c13314662abe90d066a7e90276c5631c11c2c6bf45ddecfe862e4f93aff4fd2ed712834f4f06f9bcb105f7364a22911cba7b1b097f6c4efaab86d2f9e1c30e08449e7508e1bc666f2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92a96bba5bfb2e7380ca5b149c94f581a2a6baa5161109246149de1f15ceb2763fdaac55f7d6f0f4f63f22c9ad393f7971a6225250e7e64f850e3c260e8e9f176cb968ef65cc92c569edb171fed923de7ce92cbd7a766c6918fa32d57d4db99a17782d63300f570a1092cd86732ccdca6908f32d17aa06ef43befc22152c2f16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h226d2e8d1fa69dbc1a628b9bde3f343eb6535008f7cb89ebfa4005f8b8d8a2df04850de43a495f17764c35f13372de7224d50552be988856986136465dcf4a138e49a538cf59288892804e259c0d9afe4175cd88462c18f7a4e92a464500e390da1988e52518b34aed8ce18e3cdbb153c5431e95e1d6f58174937f459454f3c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87ec6d26c4c8f0dd03e59a85e738f616143a41876e6a2e21844866643bc571c39d74ebf30e3f4163d8cb2ba66ac54eccff255f4dbcb8dfd908460df5175607dc57fb86714d49560a287505e0f51d6839ed2a61ad9e9099e6752befaf67728ebbc1e4cdf3bf1b185f1ae661af2192d749d8e9d27ab268c9efd7eb54265ae2be13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he059778f635466d951b9714d6bc5243b5f9534c35d188771592a877525895c7b14889674434f2b8ab5bec427135f937d1b7082b93d1a85cfbf1fe6468148a1279a74c682f8fc6f13b8be32cc1b06acc59b28f2df6df225dbe62c8ce114d74afb799a411f3b3b37143bf4da70a091623e14735b9c003e9a2b12564e3064791bfb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h523b1c463197dbfa0437318283b603a6ed6fa54e54b8a1f8124c1924670c216ce71392e78d768dc9d52cef9d40f8f30ff457a4f58d9f2c297da8a41fbe295334161034e68b03d405dbaa8926e53940f0fc9fa67b9fe23b58f036ece4f7291ed3b932bccbe631cc5f789861b6262c534da854bfaed6c5948688acabe924f14b46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h261fd6c9df7614c3d00304b4aedc174df3bc04bd3800255cf65066fdc2b7738b11be760f15c386c71346c7b11f62093668d09a967591949105d7c44039cb12166dfd6fb69dea536e8582425f521a4609347944e98139e2c90153490efc66ae50a2df7348afe17b9d54943250b26df10e21259e5f2b1c04ebb0d47fc0baab3da7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc57765d3033bb4d1e067c53748fc1d2ab26d7065f3e90367a784010795dae86b4b66732e153d4d404a5490e76b741c7b81c2de8f5ce8f164242bd240a6acb6e2e59c0534f906233d06d4cea9b13b00efa248aa0a72ed1a9963fa6061eb12a65affe5f42d9fc1cc73232006d19c8208226399265ec908367f940d4f5d14cd34f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb29fd67c2aaa9cedea04d9313b58d4c8ad341799fba3ac043edb408c583404953326dbedc9537c296649b6f3d1fa46ddccc3b31c39c06ce69ff4bb53d30a433fe2c63772b7e32356cfbcf3c68ac2370ad1f4592ebb58e5628288bc2d5ef4ddf72a1d2c35d063823584560da9151747d7309cf057f62542db8de132f84552ec20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8152aeabf9ce4a7654f63ec31a58907b697fdc5287d2a0b1bfee8ed17c818691ce1f5803fc6d964cd83c5d5d746043339687e452f3d17b55fdacaf4caf42de112c5379b2803421c79344ce6904e9c914cd403ae147ae3188f6f03de89e1b0ee28ae57c33bf69c612f8c06d7f1161ff99f65883293d8d87cdc25e79ca1cf1ba2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75270a443a12d0cb8f3a59fc3ffec862c697a94e1a7599e4d1661e2ea99c69f5aceeed01216c6fc967f0d66843bd5ca76afc0589e52d8d4994d441045c1b23a2f3079965d6ec9a667f63bde9db9f83d3dfc7fa0cea63ed8a9d407b1ffb11866233a5c0f19a4a7050f6a34fc6f2877b6560a1f00b584fef5cd9dcbfa1a17df4df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c642a464402c0c0451c661bd3803bb55745ed8c3f2b3397098fe4e8106450cbcdd8f6466943dd24a1c58efcd906f6e473472eed94762cdafc620d38191cdd591efb629e05c285dc830f5bebbdf1d72836b62f27e69937f5a23a69bccfc52ff495df285403eae684e6e568af3cf8cfe1216ff322a3537abada4cd293c3809711;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35c08efe433af74c330224bbdc42183c91d180a4dbfd4a8349d786c94116e8e5e76fdd5fdec1e71e8bc2c7b3bdcac2046301d2f69361925fdd8ad3df5447a148e3e2f3df86c30b54791912ff3f382c40e239eb8aa2400a1ef6f05fb3225fc1914ac61b098231bee6f6ef1d89f3cb2301d425e06b7be0c4d6d6cd2d7d4622d7ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha52b1b738e73af30b6a84090fdc17b673042c00acffc38be81b2b7cf4a8c5da67ace6a61a3911458455e8c0baf620382be9434d9ec8da6d7cf0a97c939ac0e5affc68c00a8d9795233e0e7a4c0da2491f0aada499dc5d4cd84287426afa4a867b97e4e4651cedbbd378a469158c5ca166b86254d79e665906bdd3a1a673e86d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha35ede6243845cd986cea1a617acf47b8af165917cf0ac1623138173691e52b12b86d406c824ec51d6dc9e1183ae6344b8179ed6ac44c14f62efe2bf5b3e67fa8bc63854bcf2c9f7343898eaca81db4c10b1dcd335e89d49c7d8821655d0fb015479be2fe2f4524c9c890ed011f20ecb02d8baaf5bce0d2068ceb678c6572112;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h249a0be8cdaca09d149c4389b5ab5021cc7ee9ccfabbd1682b1772815f87621817c625bf2f4d871cfa7028010f334c9b6df9c26581e5dba8f23f6bef36796e6ea4c6607fe2e6a1333be04d11a385ce0519ac3684613a283d7f25a7198246598e5398ac6f19831ea0b34c6fd486d23e9fd5946bba68811433d391dbbdc0718407;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he424419a665423c6034e5ecf4f986cdde5a3d1882cd36df0ff2177a034cdd5abd4d64c059b65cf4264620d19d79c25543828cbbe0e728a60574e1c69421f164f1531a7abae31d1f83ac465d6972106a3fbb38aa6b834eeaaf882bb8f93cc2ffa437a3ae1208dca2e18879403e2d4c957a256d112d9c0396843278b481ce2b341;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22cbfc80ad9c0b3123b18975298870711ac4575a5c5a018171b6fcbe5237f2ecef13a98fa25ad1dbbd4fb5e513d91d2d6c997090a1e6fb014780836b6c04e2ae38de44aa99aa2b5aef59b1211339178687093a2a12e723382604208b55735f1f1b44dadeee19e6cdc9f58610771884c832e4916e39102856b83a2521022bc0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd408afaaeeae7f20ecfa76260f41c8650a4879da951ff1859c884e35723ee426b2b2c826ab60fc689a0e5d4145b14b5ae3cbb4a24d268fc1c59bbaf00c8122ae306dbd4619dd77574448ba7f1510f106f99d1161844a7a848c6e09ba78a368f6bb6a712b4a0a96a5ff64d6be66b27cecb52f71272e9a48008ddb1baf1408e800;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff96f887c9eae566ec46f39b440a60c35563ead1f7dff21531aa5e46c319eaad357e9245afbd667ee38d089cf2ce29fefdf93b285703e8e2114ba67dfa19fe59406d0a2c1a3c466b678e6b0b8b927c13f87ce8237fb1ee6f7a45f55f971729113633939cba6822343bb6743351ddd24d89a80d8128a66bd5f6bca9182508fe2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb6b633a0a303ec003f566f104d1207939a10dfea1c163bbe455ce17e1a3cca2fd82a73079c4a1b5e3eb070e433c3e74f937984a8b90c52f9b950e2684071d44cdb848613fffaa65b87f8e7cfc25e1e3c653d3c91f273390363c38750ab408c465aec2e2b75ce38a2e37c285064848039752db111f2cb953bb5d8ffa66aa6a2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6f0800ac764597611468d885b73705d4cba96594ee9f007a9610592690f10c63a60a87ed4a65cf8c781c106826ddf40036df54eb6294fef746a02e0236a6d55a1ef6a9d109d6c748c40fdb587aaba5a38ba74f0ca04de1e0c226187816dcdaa6a227183556d2ace20a3eb77449cf585cd5fb0154c5dbc3872b40f524b886dda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e111565b51c4501b87a7db5ced28c2c6f64a3023db62cc3b8f1bd7d4ed23277a636c7afe83ddcbf63b2e8385a4b07ffb4d83fe2d5d2523b6bb8ea702d8f6f1f124a14439b916e9caa44f52275eb780580709b7a1f679bf644f5d4af69f6aebfd0a8c8295b138e8953eba430ba018d0f5f742b363a39da046774227678e4e2cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1e928eb8ce0e2489127bc586b2c386425d801ae6aa149df7b8bb3f3bc34038b1eba9858b01fd67a5b766b1363aa76e0a19fc32d000a1523a51d49696b532af8bc41761c87b33c034ccef770bc78365e8f02781c495670c0c8c9f5f0879dc1cb6c78802d52ebad28bd8544d33f9c6dfa6f2db8b0440ebfe1ad107d7caf5378f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6b3d90f9b3a6df8564d0cd74cc2db91fe571a2104c74aa25d42333bf91706b9e511b7969dc46dfa4843791fe7324b97be34d35aba58108cd5bd07207557bc70389ae9d752fecd738ff5a8bcf6bdbcb10398da7d4b902d18f19cb859b8ec5b185e1c60d05f9a1aa4ccb068f57eb15c29ef1b6628096d2bce34ec8ddb631e83ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bd358fc4cb80fe78956cd2814ffb808720b4cf49e8fb3ac1376a70a40f125e0b9e1677fcc2152d7f6747b2adaf0213cfa9de8d9624ac14ee328e26c78cfe571c3e31ffee310b616c2a49247224a0b307d3e951aae2d76ab49fe55e095f582f1c68b81d91547805dc7a25870c1066d3d6fdf9d6a299d20fda900088e80bec4fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8040203752c3e0acbba450a8640c4e3d2075c6e199d86ecece13d07d2dc96e7bf93ba5cff8213589658bd1693eeaf8998bdaf9488c170d10284c6afa822bbc46521b7750b37634fe030c2e43699a6fdbc6e95607bec9700a3b25720182b21485d359e4bbc28f21a47dad8cfb34a90afcc1505477eb2d61215d4c2e885c244d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf45071298d675f691d59d9145678f2ae0898f7c1bf644f65f16e221aaa4b754dcc088f5e82694095716842a202546ca474f3bc4aa5a85b623c23d7f5c81616a1a5ce3638c8f2acddcc882bb2b6ad29959c2554b21aec3634e281082ba6a34e73b99524350340251e962aa3101517e84fba9136626228b324e5e674af6b69c842;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5086c18f888fcdcd8a38fc227bf0d625ba221f58c8c3a1b1a504eb664867c5217b47198e00046997b7b59ebaf534c97bcf6fd6f4654ac823acb6ab4f5fb57d6668fe4a09bd3e2b587ee417f019d697a658bc736c25398d0d21bc03e1c142b2dd42e418888eef0795b60bb93e78ca199af088de603cc36de38bd79ad0ea0ca3d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cdb31b50e2af51205ca40f1ca42013ff41de4c4f7151571861f60d2cb30302ab5077033f31aaf5d7edcd2cbff5d01bae6b6a6a5c94fc8837667365a0fd335038b8b65680015dac5ced1b107ee878f8c9ade344186f604a3c39c435cedc7702e1a5155e95e7e3fccbfa0f57571fac5146c78267715e698e2a580abf7d9184a08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85e7c04ece6d8dbd010003fb6834cae0654b5fcb9bd22d3d094691020eb65b2c984936f8207dfff76a9c4cb92a3297612a0ca00b2c5614579e8d2e3be4ef059a876a1a16d2271d742555bb23fdf1a3b652119ce4f9ee2f7c47cc1112d8761b8b7e975b2ef729b714976b3bb0da874148c130f4abcb3f3f2876434eb8f5b52d8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h706331036f29a2ae2026adf1598a9e14371cf887fa70dae48402f47c5a2241e15289dcde4f56a4715b31fbceb7171690a8099e522bcd056f54e0990c3bb02e7b546c46bf273df4d5ca0874569c6b537a44981a90daa7511777c6c34ab7856bdde95ba21b4ac4e79afe06f28e2deb9216dc5e6602a960aa6733c69c5df525a939;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h946edc560e4ecf7cf6c67fb24c875e4ee461cd578cd282d2608755d789e0a710fc02b50b787dba19be2c9715f2e912a83d463a6818219f5a97f9b6a83237aab08c95205fc5a409d06c8339c006714a4329aa1666c4364dac81c4c8119cd891f5d21cbaf01c1212a277b206d5db143fc3e4b5d0245c8bb5ed028e463ea70ab549;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82879c8b0d2da5cdb03e5a4566ebd909f84d73b7896575be7635ab61eee3990d7672abc7d3580f9c88e03f82d85fcdac2e7dcc9e902b83e3539deabc987e6082825881acbd6831d4de0b781f5af7420f04569665711e187a2c9711032afa02c62f25806dcf0cbbb3aca0f20809ff064f96cfed5910c21532cf6cccdd1026f2e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c88a212e326093bab752a49fc83be154d6326f026b7e6d7118a1e4f7109a7a8674f6e18b459e69fa3d9950e23a47c962b60cc136083843e42947a14552f057cd455e1a53edb4ad79e8a95b731a54e01d3fae19ac5f449e19f10cd49b62e29809c4eb603bb6be826bec6a1e6c754af37a47d487f8c348f153e4bd4416f26ff6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaad78307a84c1d69184c35b442117dcbae202bbec45906e98696dd33cf56412360c3cdf019d6433294b8df0f44f39044f4fd69c432ed0175aa5579914bbf0628096c45edbea3524714bde29944cc3c74d4cbeeea843242b8d228ea91ada2eaaa97baff902bb4ef623155a63e1337c9605da2544c70faa3ac89d4c03ae55a4c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d890c81c50ffeac97a4ff2839b848b301386976cbe026b902fbbfe24f454260666b184a56ae420153153bb25ba34a588a6091d9bf38492fe885b1bf080be25f7ab97702dd91ad17580b6038f008fe66faf4141dc2ff082a2a33b196dd04398e2a05c35540f37c04558de68abf99d7e0bb5b2ebf0f266a7758e249610d98188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec3aaafa0c1039ab681d6fbad44378475853cc95ead72dbbca6a2c49107a9cfc8a350024b16c60e6d4dec4acc7dd9a9801f412f6ff4119ad34e73ef46336de1423fed1f4f120795e50fcc60525b46691db0e8d8968e3f57d88df55fc94d141d2509faa429c049a531eeb81297be346e29099c076325ea278d0750bd030e4b445;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4c08e471e721fed2bab6ffd7bc0f34fa4dbdb45057b5d7e79df966450489845be1d085be067d820a3f7f2b19bcc8b6929ef5a678ca6b2f7945a076d74bbad1ad1345a3d7877b4f1c80a5993c49da395dbbfe60ad15bc72b8f68ce6251d0fcf3d59e392adf57ac6dd6a0f2fddb44b4fc46493d275575c0093633ea181df53a5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h652d0aed8d904b6d91be74c225ea7276b597b01c7b23e1fb87261f6aebc873dee1983e827eec9ff16225d329753bcbb4087a63932b919fdc68aa011d6ecea79a47554c77b55898621e31cb991d829720a44781b5fe178977bcd6c679709348f5b4a4aa4d25f2534450df04b61383718636deed7bea62ce412ed3ce533c68cb19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h247d2b23b0fbd32f29a31980b86b7d13a3ac18d97bc8c67ae9d35ed3df9df5a127fe9f05f5c9fed5110c4927add8beee6bd9a67e986614f79ab9726848dbabe0447a36d654e8d43dffbd5ca7d568df3219fe3325278923af6f85fc41ce5790307e9fe5afb97612b4869f2fb6c6277fffc3438c71266c333a6540f741386a7351;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4656e6be9760e64364c850f60d198bd11a163188e387acebe43d39a63a2fd4361c7ee01d13e6356923f8730c0f97f8d3709015264e8b1bafb2ed9bf6267775c4ddcbd7000917302575bfca4b06cbb25eba427533b90d8a4b99294438ea3a5760f74718471a084e152da50fc6b7c024df56cffbc2faf4bb1054a023cfafad6464;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34d873d954f7f781bdca5f5a5eb68d1feaa14792bebf7b0b4f81ab20d3bfbde09144bd6664fe052a8c3db523e5f00cda258ab32a4d8622bc8af7b127293cefa5c7dd07a27a142985cb3c2409155e7dc58d21b54e6aa27424db76cfd17ba1b2289e96fe2339c562bea7daac9fa6a897e304a3faa22a6dc96a7d1ac0db5a6d2324;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99f4a1f44c09266b845759ad52252b2cab7d13520677963e707416330f08615548c4896cf17d27fc36de1897eb838fcedf6f40452d88a21a96f84eb929d1f8ab91ca5be917499cb662cdd35fb392b63dab9efcf65f02343d662ccfe2c42f22ae63853b71c50e864b8c61b987a4b7ce26ca8936ab1e45538c4bbfb1f1777cbeb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69daf1e52a69cdf03bf1431aeae27c5084fdce29635008fe328896da5967e9ea2f33d0e226e759e298451a6e7acf2652029f0f35f52c5f680f4ca520895c710e17e2753c62bdb739f5da94823772cf528e218a108006a20a0b3b5e8621d61c77d585c394c76edb9714a71bd56e6c1b1eb0a5f63e39f6bb0806c26d9653208b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38c24da74cfbdcbeed5531984a230dbdef1ab6990ca99ce84ebaeda9ad5d793b06f748d2762411c255574f5cd8b70f47436061151308a69590489220482e9433a2eab4af5748a7171ce9e98c5f704030c6de2c1c0d54b03d456e80bc81749c44cc81648435f55bb08b5e56aa43613657d5ea9b63b1ee4a2ab9194d8d23879723;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87c3fc5a87520b16c2d89ddfc0c1e68f3e60841cbb8fb4cafcf1d95dd294bd17f553aad8feed09ecd70ef434fc724bfb73d00365caae97bf6e1c173fd8dd06dc1b44026c9c3018b3af857e5e073a5cda68d9356632766ff8eccbde3d5e3dd25575660ce7c182b895c72ba4cec580a14cea8d4b0201bed236e7177f591882b120;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdadd759134b6c6abd6e7c60b9d8b6cc62499a5324ce7a68200781527b4556f2ae4439b7d4145e2dde723f30077466cbb46d893499977bb034e1930d3a26de603c3a84044942227f5d9db86498464ad512f5ad45b2a8594e015ad6f5f9659899372bd35e5b39e7a60791c25b2db9b47fd4478d6d2eccbae3bac5b0f213a22468;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39c587afb1f15a9e17907844cf7b59943ded94d84c648f2b0dd136bc94c055d87d327341544aa349c6ce42ccb06916777099e6af79efe692fe94e9b26e62d2a2e13a647869b64ed3d176be695ad7709d0c290f1e1a352ea743625d0da71655cd8acd18315a484c029b6b9eb856e8d2d2082b5bd7dc11e8bc661229222bfe3dc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba4f9ec37df44a7c0bac8ee5cd760cd84e69122524d7ad1ff8700dd48f369e5b66795d98999cd808a71f12a09859180111581109d5aeda4795b0e1bfedf44596fa1801be4f032b9763e16dd19911c24c2983394820be1d794b67ef9730fbd04a4233287ba47141fee3fe2ce71093d7e489e9eda2b000536e18e959d1e585c488;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd21dd27edd4463f15a780e71661823709d64c35d58f690c49a6b4347a8304096f8fe04197660b5ced1b1b3b9980135bbc2dd0bebbdec70ee7a9798c9d77b01de545f9a86f1d20b256c1fee60f829dbc4b87321ea9358eeee885d3806b823cc1d9474b4e92a4b7058e57f25ae2e45c8212717adef293a78dcefd0aaf39275cba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6a03df317bc773ee87b6a64a98cb3655baa2bf4f80bf990b90bca545ddfe78c89d9edc7d1cfd8d62f64ec5461053753c469c5e8f3c73b8af5f7fc13989314fd98b3d69aa448387655405e7d161a89926cf634046a9cafeb2077eb109ee7fef8cca8c51bc9b7eb5095b8ee77f832e2feed0757147bf1a4f55ea2a3fb7e82586f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72773a77cb0831735e9f4ae1ffe6d0fb136f895df2a96de7e457f422feced8dbc4f460773e6168df9747460f0af83c52bc50541c919e2c0e92cd820c70177a890d543eda9b88e39c60edca893366cb155b67bfe7d177fb014b901d2255c5a8b4f76f9a190c796d46e85cf864340d09134cf7d6f9f3d13c42402e23bb582263f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0de0970d39014b8744d72af2f432cf81032b0afad722394f8b875a6e83f15183bedec5472d22963b4eea8383ee51f1d941e68109a21afbb8c63eb81d2073380f4945411a5f2888ea355a7cb71d1a66ee9ea331e94f3379ab28b18bda2fa4463f59e54c3a0c5ae23211faab4294b9036f4190b340ceb4f7b6e4ba9cab16027fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc662e4b4630ae84007fb697b709114cdf4cdefa568375f618b6937b5862abb576337f855e46fa8d1527afc1f562ed1fbea1b1890cb1b1b723d1c7f133d25b34cd53b1ff37dbac5e02f5f4bb3a3b123d3eea0b01390cfa0e5e3ba3a7ce9c23a01140ab03ab4b8d4dcb3d649c58b513b07fcc9e982c398f25f53cf17656c1681fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f7a236af0cb3d72aa750c69513ebef4702ac2b729417dbc27b0ff7794ec4b3487a06b59f7c5a08c22528b42abbcccc3cb1ee248b8c5ad637c441364ced67c4fcedf1de03006eae47c8e9b59339e78ee7644290d13d766cfca876281d34253271576f904060f372fd51a87464403862e53be580efe97a425aca136e54b0ff9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb61d850308f201fec10e13986e600f245ef018889b02dbd54364f8c4862903a74d6980d658c61c5e0c1869126ab5e1e93a691e871b3c24b85c1176d1ea296a289d884e5f265db2205e2f494bda6a3c8c6c055561ec6a98372bb3c5a1b9b49f2dbfab8616163221d9e278e99c6b4b2877b8b36af91ad77437bcc24ace578e10d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c0fdf67e1f2d923978935c03ba67436a645adaadc20bd5fa8a75cd878ef59447a5c6b7d39d793b54d8fb6adc6681c50eee12e441c89e690976a5cbd3e01abbf07472b80e00d99e20ef76b32d99fe787b6f45d0f8d870fd432652bba2bc61f38c37832283d49aec0ee739b373d9f2cf6cb4451e80ee438c3b609f8ce3bef749c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc56c5e9a6bccb78361f606df7b0dad5f9eb875036fedf6b168dcd021d0b976bf9c49bccc0803482dd7b61d3460af0294780738184d91a163771f192835f89374b408cb7e67faa75f34006beeb65699313784ceee55efed25f383d5d428121e41e2dad566aa707a1fee8d99f88fef37a7d3e3878bfad9539e0bd744a7c1672de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcffe8be6c2e4f424bc0858257d4cc8b58a07c1b7a53f6b56ac8d8710d4004b15099625b678bc860948c7fb97db1ee4b869d30a1d269467016b4edc457ba0ea485b30c41e5fcae169ae4ca43dd52eeaa81df1889ae5fc3e3e49f547ba4c5710d373e6f5a0d11c40e4927c6db21e55a698a001a899a6bfe675d942f32eff82a217;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57b1069ba7334720295702153474405f7d6f51f56d0b688d696806bf4ae2fa51952287e8d40368894483088c63ea48db58babdbbdd73872b131577c269c36caa2ecfd58df28160e8656eb8d3fb5f7de34e965588bcf897b28b720c8bf866bf6ffd7e3906196180ced3e8042506f836bf86e6c0c646008f48134fbdec2fecc20f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f90f2027f652fd90f2fa568513601daae940c652d18c731d0f745eb3194aef05bc01c8d3a7ed6c82cdf8a4d7843689bcdaeed198dab41b85cb3552de63b12045c91c42199be38a039ff1b66e3e411eabb440412f6b718b778cbef222da24ccb078edfc41ce820290effb45ab4887142c39fb0002e352bc1d08195474a4863fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bc101fb03707ebb2b302e86bcd3a281c31a7a1ff7b516ac57d290410deb41043ef3ad7fa292a86da89070edaa49125e83f0de2f7876a1db485f1595dc6dc8652c924779f78623c471a1cfd5699a711ab008a2b973cd0fb4314fbc668b1734bf07bab979e7f288b1f99b46b79ba757628f7971f2e8d8233597bc43a7ba57a633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e52ba1f3450cf76da2a9b3ec6911b7bc2400b87f7beb5aad668970d855173c93de89626952dbb0f2484dd577b1224e560c6b5b442f2131dccb77217b55c1ba318b4744de43041fd4bf8c9f926db653ee9ff82ad3febc0be16659c3981c5ac648cefe98799cf29b0aa82cfac46f2752e73e9f82305e564646f5bdd53a15b1672;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1be6a6af33a5d0cacb9cdf7fe279af31615e360e14464424394017e1deb94144928f7802d01b90790898c59568cdee79e850c4b174012735cb5c99fdb50fcd819e75855b646e3fe1c807ec249bb206a7c3534978f61d93d8fd274a34af7f19f2c71c9fdae721db3ee8a7b7a7061eaf3cb98183e16bdf30d6dfc6646f679fb4aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb168f1bbc951930eeab14b405d5d0b395529c6ad3ec2a9f0eb64115dda8a3d7560877032660f4e10fe44e242be14ea627f2ec992ddc8b76e4be526485492612ce298165e78c66c1fb12f766143385f5ae1762d63b1f4684430a19dd3fbbd0d7bc74b58f49eca8dc9a6031670e0d4671d95eaa41d66697842cac06d07f7d5cc98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8ed7f6b58935308679c187028a4b3d69e075f95cdf658bf96c1226766c25a2f29be1650099f9085331e55e6922a3e282a1a85f83310cb2f6d0420ac7da1ee1be67ad140711d0469c3baa3e55fc757a21205766c04a47118c7a3126f9fd1bd4d03e81b65f67825c163755c0cfdac9d33af12704f20f89c6850a3e94e0dfee04c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c00dedfd764247f9909f7bcaf8b7f16813145dda69b933c3a89c153777b6225282676725e07c4467951fd7039bad9d2aa0af94578d187806f3a63869ae031d145ff467258c3eb603d8a56e6aaab4b4e8c1159ded682c0f03fa4968ede3cf8588e2923d63f4eb21042e1c7b325470942c7190a8e28faac761e4e9daa0ab01788;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9655057068f5fe2c927e84488c0059184d56799cf5de1b3400ececa6975361afa39d5532bb1905330547f5572554034895bd3de7a00f1c54edb0c3c99577ea683418700abe6aab14753ab826925854097bb9635a44d4b4229180a2f00e25ec47a35013f32390b0817e4c72ed5403d93cd1e70fc0fb5d09d71976b240cbde0662;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf6486ff62200d1689ce2530d45988215ed631669e4d83a6233df9b23fe6ee71567728a79fadf140b88ba29e0838d7a62fc92194eae9068090c58fcc01cd76b8e76b187d475fd8db190ca2c8787840804d32499579c0e4ee6ba7f5443ae80497256008bf91072e2b56cb7f18ba6992e3e8826ffdac3a353c246d3b3743bf9a4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd230bb8cd4ca7118d67091510f24ae319d4db3af53fc08ccf3135f68dfdb2c21a37e5726e55d07ef22acb075becfdbd3536162737d9b1e4a587633404576d9d82ae5ccfa484b5567e2ef86031b01911c39ec3563fafae58c3999a806b23958e36c249ddc950fba693dc3edfe76c0446cfba37111ae438be5965ee6eadb0e8a6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55377c0580473a53a63b9305dfea56ca38c3aa795ced089d35a97290260429f6c03137025fa064223d9b7e2b27aa76fe19424eadc9ce21f27dbd8ecd5c1aa8169dfa336e42a1dc983c3e57ba398cac80785e684e2534e42e590f2b0bf46ba38aae0f54e9f9f8b8d32202e3301a9c3b288d86fa384d15a48b4b2e8cb787cb4fe1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc64779f513b9d4e558b0ee0a885d0abdf8744481cb5fb99c9dbc29fa16618fc7f41cf3d3658bc552e23d2fbcc23d607fe4e304f6b675b3e364690bde82e26f4b24c9fbcff0e9a9ffbd8c6ace7d3ab1e56379d272e56656ef9fa02382233fd446f1b7a7f7d62754cc1994f0fe9bcf2141b83c488b4f98b5aa95b85c62341b0716;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf21b0dc10cb4a247b1c219aef84a3b32d4f0a8479cf74145a5f22607a6012a118953772a6aae7ce7f73e473a0b000638d0bf28e4d3d037757bd043f56291fc73ef8d2f5dc43e6bc61e4edd6f07a7cc66688863123afe708ed15aee9f2fd75f3b0ec8e90682c171339717f6ef56c1ae7857b2d15297d54f1ea428f082f67bc25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcc7cc33aafbf5b611016aca4d9f91f4c8724500780d46d41799d934492fe0778633b1f697a6da273ea333befc218a8a9d1ff74af6e267b1ea9fff6f957e9e3baf77a74b9247480b9483dad40c22808685955d496cf419df736f569c494be9cc90fa7b46ac5f078407e187940ec1628c744c5a27232775ea8ca21e7981a87f6a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6bc336956e0a8e0e6ac6f2219fe639e0ee17dcf338978e031fa7071ca8dec876335a91e6597b1b5acd1fb92253158e25b5355ac02060028b2edb8dc537cbe21d85d6603584c2f30988884466a61f91830330777ce4f947afa9a4a281b880d5360615640a278b3d31155f43997fbb95c0e3ffa7cc399e901f2242a4eca041b0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf3e9bd94b47051fc9425929ef86b3b1c387b0ecba23e770b6e395962404e3abef6f7bf7c325ca8f8452843dd1b37ded651f0aa157693634997ebf7fcc22343349e4312de9b9d2c53e6a7d79175318fb553c123179f9f41ce3fbc4d5c5492e46088beaaf65830c60581dde157f2416e4cc82c08879b8b12523e69e2839bfcbe5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb283ec1ea8d2dc382ed7173dc0c0d3ddc4687cc4b160f47d6bc51ea0c517b85eda85e1dfeedef02f93006df5caf58e19f79771eb39072e6dc024f44c53f166fe61f3cda17fe63a523ab724aad02cba881602349f893abd2dda544a783fac45850cc2f43cf02542f6d2b93f39594c3f9ecd328287aee89a149311171d86826af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9df3f330897fe5bdc6749b387158fd2a25e977aefaeabfd5b656c10cfdb880733cb1c583ba0133a27ea2b0b67c5410285a9948bbf5780e67e141154a366e6658ff47883af32b32f3b4287c9fb73b583947b3c86d7ec46faacc5e0666f989d2031b905e1e3d906e8eb8b4be7adb4bc3d87fc9797b3523d0b9fd2b2a290eb7638b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1985e53ef4bd562dd53b182a2811bd3c3749606ecf1b96463dbf7539b60661a504446c851149fe1d01c537e44463ac678d9531ed8322ca141476ba62fe57320b4c7e0da53fed24f62e8b8b8da40a727f239d410ad911b736db563f76d45de1262fbb344bc0661eeb362d48247f1b97969777cf79b7d0cc4ae960280bcf9e5177;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3adb413c522ab6582b5d60cacffc9e953f4ea0b0f609e62f43e081d9e5f268bf03b6476419c0e063049ec92ccdbb82eefc063a3e16c3b1de3d2a7a4c82137e7f2e39823fb8f2c8ac5a40202c926097654cfea695e73a0d992655a934607814bd1c76f5d1e83c11e9f91a1030575c8aa6d05a40ac38c9d799976b477ed9dcbe66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d7f873186e063a346ff76096beea0a907236bda123c3359df43b1222c488cea5da797133b226a6bf83ad33e7b2082df1e8f421df8d0efe0de185c62137e9dbd711905a6f19d47b14cf4e75fb1f537b800eb318540fd0ada441553b625a667cb86bac6277ddb067000683c7a25d94e0c26596f90e825886fe3ef8d17ef9b6164;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h928d822605c4e4a2ad60e5c90a1757c0ef280a5c259f9db9c5958a6e1e959a6131f296be082c501b1508728b720c888ca04526395446894b43cc4e89222b828c03c274a4d86e1551ced8eb27c8775a81106cc940f54dc8a42cf5ad07ae081b58406d007a819a800d43b2d27fe0d7ba3b46a478261394784b31059929c2cb3445;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e0f5625abe55b427da2b77d050e63e2a5f57fcb8da62681823432fc8446f0497ffda2256cab410cc7bcdaf1dafe8b6b9bd006755adc1cc57655001d725834b76de9e1b2c3d488ceea4cc1f0a761b961fa99a9e4928e611a6ebc92c70481c33f5eaeba1142109ae91909083df7a77a1472d5b9e6bc032a9c2c2c0b22b23e8b2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fcab45c2c261f76a253b2225d606742920cd626f32fd74dbf5cc0db4f7271236bbc8c468dba8e35a08c4c69842c49517faea5e5d084cb6cc00bb58988df621aa10418c6cefc523550587f58365928145f8d1310785e33310e4824a171debe99c2962eacb2f361ed54e53d0874ee8f22c078f2256771589b1ac128fb8b3464c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5f8aea2a77d9410d96e7468621df61b37a89d8c1e9ae8d99e06c21489cfc8cfd5885346200b265daf3c5a4a1377aa42b52c3ba0a8799866972193d27f6a9fcb5ae7306403e594b7c5cb9cfbb25d1b271666098e708d9e7142bd800c4147e90de0ab0c0c8c7d8815e2ce5007ea7d9694fe439cdd16024c4475beeb83d26f850d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha05c9be0582098027e7502591a5f6c4ef9b55dda8d22df7c60776b91b372658bd9f087aa2a2c3fb88fa67c394add0383cfc2def98e0d46385abb4159fe2beb65a49ee4b1a7f528cca520b7b4ac5751f472cae68520b3155558f6c35a23aaf35cfe671b812d53ba3c8ad8a17d3aa0d3f24748a5e2b0070b1a0f38c5e600d8233f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h500bdf0399d3eff71cd48f9da75b43f5e9279428a8f0b8571206668ca4a72d6c83537aa121bb9d5013f49e87c5787b8f385bb62c4c129e4f1cb04519775ea038949631491d8b43fcacc9a224259d286c1180b46aea0c90b1d2ee3227ffe3059f38b8551b4bd2f14188528efd2d2c3b74dd71656829bb0494bfeb6d944e4be469;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87d5c81e7bf8dd4308f326280627f83cbceebd5930218b3b82a87a6d1c3465d137b6f150127fe6e57869dfa95760f93a29fbe726e3d8691a4b371bb91ad16cee813114a4988ded5cee417c34d9b9feff6b869eabf8375c376cd7a7f50e56ccc127fa92b055f941e5e1f4ef8a4f394c964c1267b04abf85928c1cd73c96228ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had1a326b4b49c2089b549bdc0e0c1f7ac8417c6581f452b12d259d3ef3dac17f12b5f04774f6326c7d2d82e917d97470003b3c6e121d30b12eabd902fecb9ac5463403433156475c0565a2faea731bd5685e1a9e19d28bf34d57f7e333acbae0d60bdcc51c3f981884239114beba1635dc0c38c29a29c4626ecc6534ff287320;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hede84612eaf080eab4274b90dbfa1099c64c289096fa1f5dd972ddfc67467d591e5101f79e7d9f525bb6c9a515f6bedaaeefd96632b1b49afc40cecec298c4f9bf7b18f07bdfc91130007d881f37abe82b7de4d03de3df8a1cbbe630a49e4c2b4e4764bf5b60ce98a26724d1c50cf280079eeaa270704215eb5ff3b7f331193d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b5a3ec68b6c97345ce92f8edd5935c73d1cf2015557197bf8849ddef20de77c794d7d5d0567492c573ad9dec5da193a0cdcf988bb747ebd19b3d5690c5f252811be7ebd2a7aff16b14607efea34d28e1ccbccaa4d234554b7b13d793282f0b8494e66c2cdaa2a6cffc4ad80c380ef9ad22cfb28c2b3478d91c1c5363c461bae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ae3afa62ffb3477fe1225a45de92d744dd48ef5c5e667f458e61dea1919b019c9d99b42405eb8270cbf9c059d10ac9f74ad35f46704c58b95988fd87ca1c002ae3c349435549eadf37ee64d954b9ea123f83a33d096a8d7009b407b38c770f9861aeb7b7b6f1beb4bbd0a7a28db1a34f0a6bed9493780a5d2ec00d50c30d3b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2311230e84f2b316b6027a35291de6a1994f4d0770597458700584be4f5b9149053a6a08bbec0a778be373051089424e4fe363d856c45be5b92f45db8549fd76d3984b82c731358df00db018db95462427216ffe51b64ec87f2a28ec5a8eadce4566ccc3435adfd98853c2f523a35e7ec32b81eaffe7f62ffdcf84131b2167aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85b3e44788807546b05c63208812d2ddff817f8cda4f84a3d020cefd707cade8f1a525f6c535eec2735a8de50554d57c388c206c8a991ecff43ddb7a2185dbfce3ed48f5bcf1663bb6ee0da0d039ee09fb63a90ffaed1c0e85a3aa0f4f4d048f8ef697f40aefe3a8084bfa419796cc32a921fa168f77cad16881f1c8b1d94493;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h987a2a952794c9026f4d360833d92f397c015e86180533705b5c7d9727f3fdd597f16d4cef580b4af9e4e253c2b95931288c36520aaf18892511af8e17826cc86a19fbee893e8a0cbebc01fced99ab716a3a7ec75ad3cfbc3c67e8156f2d4036cc0e2b8e08c90769eead1a24e582f5c2f4d3d989663454c8f730fd9711d7e43a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf864f8dc34432d434075da5fa98227ae5738234fd3172d8d85bc666d8dbd24ea718634f273547b1e0eb7009dc5d122740327b5d63778c3cbe717d770e4943ca5d780f5f2417b719499d8d9c617dc29e7b65927de867d7be2fac90a5bc762772b9f2e202cd3c5b3b3c91efdd4d154dbb64e4d1d69dcd8a9155a5392a0417ad87e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc57f81b384487e687744bcac5c8e5eebbd2b019838b18ee6de3e4b57ce1cddea00b43e1a1aed2e1937595f58ca18c7029fb137ca35b2b88d25af669f2f64433d2b991bad9f82ebb037a47803784c813411923a86c25e11c2c125e48ff79cb5352f4140f6486874a9d062bf546ed1d5279b8b5effc284faa29be9ef28544d778f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4ddbb2ae4a8560c414c3e99370e7e2b21177c297916b300918414ea41788b7c987b4785a25fd8491274d78811f836034174940286832a80a3caec3077e486f10179eb0c0e7e21c8d4306989486d3e865cb40b7dd7b24accfff9971213d21a376dedac24ae5945988101736ec0d55ea6dd32bef462f148711b06da38b762d2be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42dcd010e61ccfabc1a9f6e9515a50f05a1c566c75bbee0903bbf6c468e2a27989a08d74974fe616bb3511375529c296c11c6ceb300d5493a1cee8fd3ad6ebb4bc47d1c3806a2a16d4ff0a597de1cbd2612f7b73c94e29d255e5b4691230fb87fcc3f062bf1281a1ac6186315bf0701a27adfd786d0c13830ae8b4ddb7c224b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b631482a6533ec158a22a98fa999210d5130485507d9ec587b2bd642a9941de4a6aa1ff66d77a69c717e4d5241900f2dfd72c01951ee9869ee5853b7a263e5813baa392d137a17efaa53cba4d88be474ed9d6441e396340dc83a52cb1e23b89a716831d10930261f05717dff5b33ceff58277db975a50e61f05929b693c83ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74d7fa957369a2c0c6caa842e509a100b637758771ff1fb858a873089d4d41909024379b1d483ce3a13a529ae8d5ade64ec9de04ab249bd1628a7b5f7006feaf4de5784c1d9697360e2691fe736b894879ddcf0bd877e90514712158990c191e511c252d8c7efcb3378efbec7d27f880461978f2e9da07d01fde191b24a26571;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb41c5eae090be3720f6d48efedfb61fef54ce895f95765c0e816bc0eecf03223c0ee8d4b0ad0e9d7f43492ef57d748e06db47c7781aaf08d86fd483e3c48d963988cf295c7318c748fa916a23ec804047c3f5eca9d38065765f3d921b0f6b01e8e8a2ce601a90818602bdc9a63e2fbe0542c1e67fc7a72377484d802ed1dcf14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef46224a5e76df8f25ae012ec5d24c205b481880ff33fee7457e49fc6a86e6560571caf7e91d3f0a0bb5925a805f0e1962028eabd6741a7283ab42bb147f09cd44e67a52bf2b06721a02f989e6dca7b9d98b98f73d828097716eb35ea0f8d1da0ead92dced35f18dd3762bdbca828a14669a583fad1ab54910815a92109ae3d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc532413823dd5230fb46f00c9ddfe1d2e0d49dd3c836539306de481e57be112a8c5880953b22f240de3d03842c2b566f0fef89f3e3c95b5b7e10370c26845a161f6f9e8b794b04a6f61926a444b381de79ad1e132928afe59fc02907dc0023ab939728f6aae28759f32e58a82c5a6e666619859bf8dafa4bbae884f60315bac4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ee39e406b17b5dc2d000f3c68928ce8268af50fe09576b0301e1cb5e1e3bd85e52dfa5dfaf5ea7a7f340a9f942187bc87452235f9997b71bf002cf42530ada97e320cff48bbffa8f07e0f7211bbdd96673f02b2b18d676de7796f8f7b84c3de75ac53daa393633798e84d080f55e67629c0a9331e5f0c6c3b9ff326be2adc87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f88c1b4e739028c2d477b70937c2443bca096355798519f00780068039b68cad70c0d66d3c32237d59c079036ae0cdc98e55224497f94deb29873828a14548529e0b22457a1cf821b814a254b820bafdad7277f516e13ea2e888a0c82216a2a21d9f183a0d52bad28358d41e8850f3a24f3c89e9fc346338427e83f47baa870;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd681b0077abba4071e2c91abea2b72a36a229570d8f52605d8dac45b3e7dea8d27ec9e3f47117500e59294b25693e9b4a91ff497d5398b4e9593ee5687e2d6914767484d55aeca5854de46a7c751140f3d111b9043e220567c0f9c1aa86059cd9c44e9f58d8a907cdb9bce480a8972e3499fe0a799a6e1837b567be2489f6acd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb77f787c5322bf0ddb5e2ee055c0c6b2dfee5e72abefc36929e252458f6f88779b6a1705d88f705c9f765b486bdf0b4e0cfd8326becceb765089bb2040c0aec7af76ac20f5a997d2282f8ba79a22a784121b929f054586eb58e864ad21a27896b6143882995bb00d83ed9861e87656f82303ab6bb7dae3cec16e4dc08a5236e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b762b31aa19d01c1ca810c829ae6a5e15205fc44e065ad58bcbb1522b38018159d697dde133290f9a55d5765ecfc6b60764febbdd624474bf78fe54cda079b8ff484c9917570b1cf4b623ce3adf6a77999a809a011fde2bc33dba39a032f39614dce961d56b7f6bc5c9f11db55b78b1304646cdbcef42d17aa0f279571c2a2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca3dde8f642ec8e4b9c5e034feee7588768479bddc2b16903bfda4e45fee68ecb3e31ac395f8b5235b54184f021db8ad65408bbb16444c49cc8d89845b14533e6c759a5cfb37563c15bdac885ae29cd366f0219791880949ea15a9bef7226808237d5bd96c2a7507584b301cf084f9f53ab34161b7d87e26361be88e16c6cbbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h790ae53db6dabcca34732a54231d72b04581b9c58aec95b2cd7ad269d31c7f27055ccc2d5b5349824f81d81a54674ec3ae7878ea37d631e7b700695b81ae2e95993667173f6c853363c2230331ff2a8dd34836b7888bcb063dc302214e4b36d1a17d4cad0d405da32cf11a0ade45961388a5c95305101c7796c8dcb17830cef8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25ae347cbd35499cf856de20b5017c95d9dbdd26b2a5cb04e0802697506acbe0c2441f4d592f2e2375ae5ac1ad93c9ce2a0da1c7914653e616e50849df6065978264f54c147a60ac1504a95642cafd02aa1601332e7fd0720ec2fee9debb73efe2970a873c4e469f22c46c46bd00fa02463d394c44f327a2c91a7247c3bd4270;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9175cc9253ce487b60973012b6f1d5da9c78831309e3b31ea589d2457d983eff4266672c6ac566378fb0ad66d6edfc5ec301abee71f8aa8c49cbd973ddf119d16b2e3ebcda15316a674bf354e74a1b89175b1cab9a1cb6aae61e8fa4fce7fbd56d2d2423cc19d15f968e5513aec2aecbb7c91ec656baaec3033368c10a5ab618;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he836ad5eb5a7ee3a735f589b5447517442eb9a3b00d2a54c86edf79702d44cb90eea68d78d17635c2428f3968c7dc86e4f0d7a85ff6c212c2af0a1b48f1eaf3a555ca69554083a3fed98e242ca89d74487f19ff68fae075b62ca062e37e7e00bf8fda28cf5d3c827b388d13961a4d54d8469531bef1ae32736b277a6cc97fb84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h849e097c5ab393fda132c1f7acb13e474057e579beda4571ec4f77f30db100709e5c8477d6eb92a47372426ae5818b8c4aab67db1869f36f8e2139d825bdd9bc5c38efc92015f1e831dc064a4c6671036103a7dc40ef3832ecf76ee0eef26c30a064efd530b12fee00e91dfecbaeaa122a45975bda503420f4c958ce901966e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h204dd51d4c208f6d5ef7243bb5b312126d9870b4b50c684019c400aab2a25bafe13dae36d05a5e2dcfa6815d2e542fabe37119e49542ab545f19511e5193e65a461d7d1b2b1ed3a8ae763a261725e8cbddc2db72ade27abf35ad3299edde16c6a674c0efccef1dbfdd9c6b98f910083fd0a2667ef6cd853c37d0596240ae88c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcecff616550f43dab92162f4db6b08427a08c481ac5c539f9296aba5683f736d12f52ecb73df20576e5420dc666029b8908a7023ce293f47daa0353d6ba1782706b823363a313c5e8a4ffc0c050e2b282df07a0d4d08f3d2d666885ed45702f634d12c2bdce5ec308165552473649ccfaa14fcbd7f6c99ae54a518367c08d51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3036968af80341135628d4554a9fa7218932f212d372a018175113e3424959cf0357411ab76e762b5f9592a97e811b3733140c97b8560c634944366667c8704d3470d347755625198d05455c7ae3012d00875bac6432a5c820c7cd3417e23291db91918762983f5faa77d88a6186dc3757f576954ff6b1e337b0f28d6f8e8d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7236bd0241f7ca282d50f9728e5019730433f5299865faa69ddd13eecda6132ed2a0c8e5a9ce6ac8544ff7926409391a01d36aba5a74eaa15bdc354355b2a634a3946cb10de5a73d9c42484347ff5bec9fec8bbc6773cd222ad85db3c9d0571f9ec59f3a6bf34a36e36d1ba5b022d31dd560c1bed7c77f426f062ebe4cd42daa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb80ecb806a43d820d4038dd9fb86c1d27d5ffc443d9ed33941c42f91ca904dddc6ff831173bbfe62c73641b9e92457dd5702c4ba22fcaa1be2a69199f29d0e79487f13a3727105f53f38122d974479c03b692013a0195e5aecaea6b80d44794bd36af2513446c94d408f03eb86ebe56da93d1d14155862a0016d10c2aae6b01b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he90636e1f3ad70d8bc2a4edfdceab928f0e9dd0bd1293cf37c90ecbc73bd5727305e5da178475446e3eb331e471c69afedc8488d4d2d2ed3b6802a5f56e649373e9efc7bb5dd8c9ae86ab44cdfcebd20d79e60633e2e577a1969c53c248a2d6bf9b7a9b175b0440ee66829d4a5dff6ea50d6c771b7aa42c1face0556ad18e3f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he095fb0e503563657d8d00bb0688250d9040643372f78a2a0fe649e7ab19e298e707e409c83377c862284c427204eeb4e127c0cc52beabf6c05556fb07872d544f1fdbf25614593e86672a10fa3b0205a4429564ee89e473f1ec84b763e4d5f2cf0a351a92ed0a2a89c88b24658d5933570485aee2f34da853ba9811b128cc18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cb6642dd87fb3c0a612c8e108f4e018ce36e949d8594b6b18dea94b38edc976cd6866d72b266ce04065f35263cafe81ee2a7060fc442ed7f4ef41a6039f2c63c869093f53bd4b81c6073d847143b7efa12c86fc3d3cf552d8b72ab5238b8d603618d99acbd752bd33808440c69213e6e246118bfce8ff7f9dedfef750dad102;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h752ad31841d2c35df356cd3ae4fe884361ef185f6899039be8973b27a18d32e3685a8a43f719b5e2ec6b90a98d7008a922ee19c6262da18d90bc339efe41efb6e87eba3b9e5ce2ca9f7ede66d24e985b80aadb24e512fa1a2dc9171bb53d54b332c406cf11b9c62daac611baa9be8b03bc61fb6eb9f9fa07b8f3fce56876e0b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94d68da69c3fa43b4ead870c05cd8ba8c60652f9abb09488e5fd518e63ae59d305afd356c1aebbae725340a1b3a1009778c40f1a702860d591579886f918f27572dfd50fce57215f3bc4f438a417109cece1f91a60d2883ec527a76ebc683948d0f7e0cf396509ea27a2727cd5ec73f1406694d3781089a9ee2dc91de9c11bae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6844efcd97bdab1cdd58e10e0d3736d5c8595e7f1e1fddb90fc9d8040932db87e220b225a608f677f7950776165ad1a132d7b1d047bd4164f1ece747f4291e9304d59189bcdb34186a22d174bbc504e1366336f87067d0492f8896334c53108751eb2178166dbe5f444c643ba5997a384e20f2c0b67db714e64a9924c6bbd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8882ffa88594b29a9079849faaa0dc7af0de69af4d8928a95ec34e4cbe60b80c17169f1458c5bda67996f5278f885c20b36257db8640246422cc80d48b1769b99f34d9f9a6212a9fa67434d3d62e24bc16c78dd60e90635602c104a939cc1d5a02d6a5204c0c682a9cc09bfae292c2a0615bb7923adebdc0168d107d4748b7a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5d7a867942d365a5cef04c9284fa7817ce72c2fbb29799fe62c480e5eb3508d33e35b9b2c4f0660bbaea677a3cd1838aa55369d457f62ea9b488635f1c48b64dfc0f7f4cbca297f3d17b046127cc58b51612c37eaab5bff3df3a2502ff11bc716becd5008bc93315fa33448dcce81dce3b0c794ba0e2d00c4dd61c0aa0d9338;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he71006fd297123dba4b20e099a0da493350498a4e868cb5e7accfa7eb4f711f22ba419abda1ffb324069f7d14dca9a51c38c60953e1ff7d4a53e97ebed207de287ac66a0f75eb056fdf07b37e9e3552c8b8aa4c585e205d053b207e7ed0ab50784df621f82cbd22e368d9c4f0fb946753300c133ebb97bf1206828e202babdfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18fa7f61deea283994b5aece889cecb27f6e27ca3651fd17b58242d75124634c35d68be8b2f4567662499b00824921922c89449e45b65a9877aee49b7944a03d8be957595429366b26f2a004f885c7c3ec9fad0727af4f20aaca20d0344ff52f796d33db605947c30b1ff0bf837f58a40989b6292b1a32d5fa8c13ae907281d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffa3dbebff27c25f4fcbbb993a6c7c2e180d8d174ec894bcba1940189ab805298145db4fddee846a8848a3396839547838602525749a089156ea27a20d4aef0261da4d0b5f9853fa52dc4bfa00aa2467541918ff6516a9feed8136628e469e016f616e955b89f0de3060ece35b04bedcb38b0438f2f9d231416dc3be25c687de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h217fd89ee80773be87e2cf0bd6b107acbb2649e1b5c853a389bf42a4c4e2315b5ef474c647bfa9b87528d0add94f016789150081922fe0338dfa2844d1ec01f4fa7bdba3242f6de262280898c81166f59dbd00c60f0f70ccf1a812dad1da7ed8624c858940cab30fc42ef0fb0ec398d077117ac560ffedde2207a4bde13badd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha333795b505a566a10ab189520162d9dee410e18ca68407839d3674fba31d9678943e3e5b64709a1fc09f5c6195ac9fe471db9b1512abfb5c8ef806ade9a06cdff39134fc70dcb0b355a11764d05c659e459a2bd643cccf2cba5eb821e02dc9ddee5c6c9125e22869bfc94b7b5883696fe13468bfd37f9ff90f750d6e1c4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f449f30c2708d8ad3570ab42b3b9347a44f0c5046e0ed8f1145745e56b1c0ae75062d81b078c75f31a64351e2486b71edd7230c80db5c56a4ea65851ef987adac1e4cf0cf5753cc01ed73fcd8bfc6107ac1a24984c2fd85006b6c26a3e59ad72911df5ec56a1970adb09921de401ca07dc3d0d56101d49dba9cddf4e8adf678;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he25a82aae342229cae5c5c1d4613ef91fca4e95ddb94a6c8954b9d7832486c7e65aea592bac9085544bb97493ffc5611f5d017eb2b35259d5850a5c542aa250f6faf639c6b9617ce8aa01ef05a3e4346155f919780da2b3858a90a38b68b09db514a45c4b8dceb57db594ec6662109c50c444afe591a4a6dab0e6d0fc7ccb47c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62bc963f3cd266fefb5f92f65232631b0ccc416a5abb39cf688d18d585f94e5e71c136635538e529156b089c97ba9b198d26469037b7934161cfddd5fcb2d70d64277a78e87a71405f0375f75c521a553604913200eaea0f27c491ec07d46fec36b7f54527eed728fccd9c4c601c23c864971f1fe717f5e862bc4b8b6d779494;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5804530e0a255c23215e7f10cc8ed74d675eb86796055a95dc12633b51823d586b83bfb3da3f7d26116df476391004af1a089c4d04e9a5df91c5ccba2d60dfce546d6df125ee85fd959018dbd61abfa14a04e77bcef474ff4af9940ca87f342f59cd0e3b8467a0b85e44022c639fc8173a631c9139559d2f425efdeb6de898e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dcc2f2936e95be381cdd204c9b81770d2f9446843fefbc9a4470f9f607adef896da62634c3ff025111cda085e100fec2bde533da366d1d00bcd9671e93aba6d1442307403933022971032b4eae990bcbde96b7c1c98039c8694b646c9816d9f74772c8afdc554b5dc0ca3353d0128c74ba597dc2bf4939d57a8c73b3c15d4e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4303ba6438c263cbc5fee497ab0e3e2db24d3e7421aa651b69c9d299c00ede27c6a9eebdfc1d8248f0ddccfb8a09f7381c7af1220bb9a034fcc86e2edb25da9d7ff6a88367deda8e959f7fe5795d735f7592515f50efcaac4f2db7c0bbbc10b13264b008993884010a1270e1a90e3f221f25a4d67e3dd6040ef8406b7a3f82a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab500ccc8e87be853d9993a95a228e6c4e0da4509fd30a20fff98c99a1388ccdfadb39f95092246134772454c12050ab2bc676295e4828ef58d757ecc963277bd225dedf274c3dce8b4e9c5d36b28fa0660d28cf5b5a62adee41db729db8e528cc37e9f220f8aacd4a5843c8bcbfe914b2d2cd7033e4ba487bd780fcccb68fe3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b11a8021134b3721dd0de836d1a9d2de704fd3a667d6c9582f5b9b7cf222a35e7de8bdf8ea78a4e29879aee0a3a79ac3bcb00017b3a239e9dd85f42cc6b42c689b98b54d78c8109284d9d3199284f3308645946f0eac211468d79c7a0eee2eba70e07320052056707caa47074f818842f1ceb1e76c688ae8630945d068d9ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6453b4b7d7f20fed3a2af735f6ae83077e922c679b4d1d54fb66e291e7955a4ad4c19da02e560b8522c3d41040b746c2c5700cbfd157793f9ac1ea6527eaf79abe6dae20124ebe675d8ee993c8b404766c4fa80cc1ba8f18719362ef069bfa878ef6983e2596a992e8fd0ec53e3a37aadeca9acdbaf32e267d7a7f13dbd68c92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d7b47df9109c091642500c5769168638b4548f6f719ca8bb4112b7b32d1c45f18875d38d32e2de87cbac3cc4dcfec64c705a56ed0e3bf32d72d7f13fe75a0e023eb7bb5b9b97be724e15e7f26ffb6bb3b90ee4599abf4fc21a623c5b175a0a90dd961ba1ed1ffcb414172e0c7f7840226f4ce4adaedef3b6f5b6f49e46cafeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h609e59d962e63ce80614cd71e847005e4170e338b518a0d23ad0034cec983fd793bf6f9569408bb0be3f1ef724030b85fa47f4a66f06a93f7b8dd1acc24601b0050568ab49d0d7d7f005cc0c19156696ad48fd4a90932af601245d07cc53fc63f86c04757ea14b5746450f68407093d5f53eb11dabf0c6746679676987df9f73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5da7209b3a72683d7fd3a6cbaf0f86e2c75df1c79cbe086444334a10e599af1bfe218e45b3a6b4540e4c0d9f68dcbcf14d44de0b6a4c70b8c67bdfe7b99e49458907d6a300b423afa790043fb28e869f984f3fece1b8a54eb0c4148fc1a211d50bfe4195883e73f40ae4384edc3fcb4d6b0099d4bda0391d9c2ee8ea80995ee7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h773dd0ffce9b3a1196242608f03fd7fa3f3204cedd59ad5fa85c77688c1fe56602aa9381b7a5f6a9bc15269cd1ddba54cbad123748ec38f5668321db719b88807e0a5c4f018c2652baad9abdaea52aef7215e35ef13a86b9538f0b287cc4598f28fbb18925a61e4301e9a2a9ec470672fca0b7360108d263ff1a41bdb44c0acb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h971b8f523cb152d0a38a497b405f56862adb529a85715ae3e1aee55c3b002c08f45cdadb3c11c0522ecbbf0a9a25b49191c0dc8a49c9b244695f985210523a7e519709e61065469ed79395fdb4870fc463d4fd41d0161d26056501a648e079bf99a2b003fe0416835ba42e744555bad7e09852a82a87e3756a223fa3e5165eb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34face61eccd1d4a4b69c6c54350b9213c958fee95dc3ea7026b896b5b81a9e3031754b71819a237e5644fac50e7ee4e5367dbca9091c567d459063454dab3a678b2f92a185a774ac1fe98e40179897d1b5e0ca7d9d6cc71abf2a54b6265b8c3a904ed666b900736ee8807b1dc15f7741cfbc1f3fbbd7ccf9bb72bace8a33609;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he00835ab766e84d1de0be83919a1d03e3bc4721798fdbef6cdf868f0bd855ec4762f4a7df7cdff7c44f4138df7aaff8f4bab72a5a08beb802c058848e5519e7b4f6ad6dcea73e8fca7daf26c3e1d53357874ffe30cc6837e6f02665c39c1ec85a4af6ac9175a0e58d838ffa98a2d63595a790fa802d4d84bddc5ef404841b27c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93e9e6c6c8c89725d4a220e322b5e2a9a3005116af3f62d22af6625f33584f253e398130525130827a02b8ace3810b647cae88efe0f18a0159836e6d34939db057354db295279d581fdafc0f4e253821a4257cca9a6a69e9134384607455a7a793396c7693e8e0ddf0a1dd9a5526828cf8f3289763117c68fde59296cbd67c78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5849d8d279b1308a30f0ce895b4f2933ac06ba2f9440757e669891f47ad9fc9fad67df3e2ac7d8fbe894a0c882f3ffcc4f08ddef2cae9c25a6937be6fd539380b6c39de2f8dd961de61721a9b5910b4f3f35eeb48ffabe3d2a88550a7ccf0604f50db64a0c7e79a25d9753da279375f38a3e9b9344179c8606574af71bb1186e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66f0c1eb7ad4f500ac6f25206bdf256f8da4b00b4a8c9958f3086347a834d9be70c4874d0bc518b580c0d361996a6857a48cc92bb2c4dadf2b98694b2d4cf6022fdf9994287f1e298d8b96e0a1234b055b4c42b55c4f7ddac28989b9135486e32db8928cc29d3c7759e8e5b717f1a10f4a0f14679365b0e162bcd61a66df7d61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27071709da13d72bffc808c88668c9e205997959158be7db94060860102df1796d4f534363207d5eb92399780a965a04d4c514a3edacea32b19b34991d44acabf2b4ea03833b9441b91527762e3e98b0460a479db9f42ae641f175a099dce928ae162f0b3cb16620504abc3d6e95e98691e65058b7bf14bd0138f6de74d76d72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3099568011276fb36d0ecb90714d8fc2000cc96f135964a3543b0b3fdbfb42c139cdf7eed1989f6a4aa59eba097ffbccbbf0ae9ccde581064b0f53d778822c8e4491ee5e53a3aea326227192058def82eefd3a5fb7b5a2095c033478d8c355d0eedd243bede9ce3fafb7e7773cdd129a659538ddc14021f03cc72465e026d8a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d1991b22dd25cc40ebd0969590e8235e6099561668b4d84716cb976803c413be1e69a80931336ea7947187bfc03bc373a7cb2fecdf3e3e1afdc085b9701ce91601a58dc4b0ec991658416fd3a17054637ad3c2d6047818e6543fe571d694a126d47563cb0359887e01144703df8f4f6a316d908db8015e0e0bb2fc5c5547d98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb749724b9dfdab0988c6703a2793b31de28b924e2550b1501577a102be41ce4093f24886eb96aa8fd00b2968eddcbb6571eae7014e78dff0d4544f5ac041048f1fc1122489fb98d32819ab5020693d01a02fcc39707fd39efcc8662d4c6f75c8621a06bc756ceeee684b719c45c806915563ac68803e540221d508a8c8ba4f8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h427ce3c53b5209c5bd5141f35e48658a9424496f07e93e4ff3682ba5010053b2b1a2e6ef102c8f87d52e6601b9d530dca06780d9c831457779c1fd56857bb8f1fb3eb61c8dbc53496de59a4f481f89060edb91704fdb029acdc19b9940fd990fc2c09e6d7653724291049d3634f0989a3bd2193c396b2763861dae5771a42e29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6165dbb4956e0ef6428aa6e9c18bfc0540cee7f088339a0d7168a3f557850058f7022e9098385a46ee936cf5f6b03ad2fdab662b1bd5c007f484ba0c5f2904bd35b2fd5c78dd652d584c852a14c4759cb2d81a12e8c0f59328033cfdcdccca66f7fb5357585ae2d3e23ffeff9ffee4d7b8a0e01d63d7e54ddcecdcd2be44d0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7137fdcefee886a3e7940ad02a30d15f8c3f1b4c3ac76aa095529246b614e3f93318d98b6ef6b7fddc956add5594208cb63209c65dc6fcf67f3223b6d318915607ed6d57c14dfe2fd9fff211fae716bfa0a6da070fca01eb7a6f533231023267032a7a11f1decedb1bf509267620d15d824f1011fea6aa039a6775ca30c5e2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30b4476ffb1b6738740c1bf9a24f259358442ea8070cedfec02aee5963039435303650f96a35e3604f669e6c6ef0129bd3c70d1666f2fec480fd080070a9db4df890dc72f7bda9a94834a31fed058a3e0ddfce54ff9c99f1f7ad0ff182bdb5e5e46724303164560004fadb53d33c8584f357351b8efe56615b072f6483a25679;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8ff91ee3f5f7615f2dbe8fcf4c8ce93103d1ab22c8a6a975973752b4d4e97cdc848754b7eaee507efadb96426e8beb78c85321d202e07a500f13a2bf5f18a273d27cd29fc07adc40cb14b9aa088ba531026ee1e25ed8224105efad3e4e2d710671e46e77bb76e3a165b6d19ce863ab40723c8f42edf56cef9ab56bf27889a2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30b1cbec5e3dbbe1fe85c6da7b75a4b45926b687ef8ab9a7f6a732965d970e10b992faab8e8f929c186c3fa7ca273a94fd11490d131ead9ff33eb206f3e5a41ef14bd1818dbdbba0970bd453a773a47d1b4d1b6fbdcb6f22f85d0a2e466d5ea902343337b1392dd8d1119a580fe9e450eb33f1314c50a89eb4a3f64be5270e7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h383f61de47c628cecffd24262bf0cac0c4d56060cb9167f51ea0c89336e3224187e5e4922e4ad7a99a80d42ddb567dc4fe8fd083720ce0d5d8507e0065558d6bfffb79f8303c317767e5e7d49a7f4a9bcc130876a077aaa2d992b949f98fbdb537d0c250a65a3dada5248f69498adabdd34d637dadc7371223df667faf2af30b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcff0dc8daed141a91fa1f09486a397c34f10a08a5fddba6151d12af70acd5a56bde86cb113943795ff92c989ca14f30b437ec81c593494dd927c79105b893cf949f306d8d7f43055a011e8eabcc60b552648ab278476296237469f10ba1f6c62812756c0523759e69fc826daca86de612c86ab1f00fcde998e49bc2f5f03ec4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h806bee3e4398edbc741b5db5ec0de990c8f86e43978de266492f7fef4e001e445e442d94b56e803a8a6d9088a1c630d0176baf152b92035a2c844fe9db705b911ed74691d1565de74cdf4f97aea6e92b56f0601afe506defa6ae53b5be2edb4ac14d8a69f61e43231dc28f900182e4aecd3654bc81713b2df1b8b25e74c3a85b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h321317b31c556f697b0e4361506ae5f217b7b163d33555875af8932912cd61a65a4f562d859e337ed9e2ebe3d8d75665c059ce074f50f3ac25f0aa509de11dd118d23bc173d002f6ff3063ba3c1555584522ca3c8508d2953c40d44c73831abf8fc5df870edc9b827a59d19fcd8f1aab449b5ffd283882b7dd19e2e64db9c0a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c03e5c203f61ad6b7d4888267afffb916c98f76ae083b01219bc5765f4d89305eeea04d576fea761718443c08f16ba2ef1b60eebb4386364724d6630842746bdf09edb59d6349d17d89e18ed99a32edda72d38c2cb3edfb3898a4c90f21b64ddaea4137c0306d7da1d4d20cbd8baa7e0393033a9fe5181248656328498fb48e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c3e47d0cdf5e3d3191871abfdf5a28f3ab710ba199e6a73f9fbb1ac19dc8096546d514f1308d015bd89096a4418ada87ddb8282fa7b3f996607e79ce67c6de150cf5de14c29d715e58c8a583be82125a6d87c79232d40fea58f6e4ee27ca30b8a57a911b2405cf1e8d8fb2fc7dd649351bad5ebdef30872b2d8075470828ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82a7ad0f242306df3d763142d50064878e07154798ff80a8d01d3c2c484c720a125e71bcd51cf7f09b749f1a80d68702bba53e542e3bd30a8c5b1ebcf5f302c553bd7d05a28fbf7feba14f572e883844fd20749dc6698fb3c9189fb9d623374fd3bbcba918f7724f1791d8985059487bdd2a5e784e41458000a5029ecc888b72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h172c9305565a8308631ff23774ecd8aab190cebee7df0276a07b66f41aebb807948a88933a3e380ea571b4edb2d6954ccb38bfcaffb93f8beff8b82f7b6c76f9cdf796a26bf440ed8c3bb69c0005d29dae0f3ce647877924dc69b1063e6f35111e254116b4e63db20fc11cb02f1066d8a3c1ad787b21634fedc008eb3077fd21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd99272fe8d0c4e9d34ae04009101ae2b6c8895dee3347323a196d478eb5847ff550e6d166d3a445c67f04521b7d02e0f5d1aa8f565fad082169deb2b9aaacc27f34f8350f6aa068725c25dd71ff25f80898ba70f689c798a1ef295641d5d7d3bfcd3285c5b55af5148a452b336ee5c278817f49c360c8a98216cba5bf5aea28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9abfb07f50fbc11f1173c862bd8c09ab43a416bdd0d73613b93aa76013c9149540d0fb5dd69840137eb757c63e78758ac6eb0b201ece5603a4748764a048b8d279a55a7ca43e4d7b5d81b1505e35b5290272da475485d319d6771b125510b984c99d2b1c32ca56ecc6b644392ecaa16c727d7a8a30a866f8f5b1e407da197f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfae70b11707f5ca56c180a3f2532d30e5a3085fb7a2b0e86304c19dc8bd11c1d07d6e396d171fbb3a351f49e2186daf9cfda99fab56728b5e125633119a37073ef03575f6a8c355053e614bf659e1d86209a228515e771ea210a51c205d99e2a4c1cd36513b38d61c77d332607a1c5921cfd0fbca4ad2bfa0f9ffaaf35c0c2cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6982e510d5efcf5f5fc7f3764378a684091ab634280bb618e3b17747f52f6440568ea7673a4a1ffab2b29bcf79396413fcce0adf8486b319925e788716c2fedc2c74ad57fdd7991676c057b6ba33787d0062a21e108386bebef4c5b692c9eaf86787e3b2c00acff476a92f329ae698e85cf05afda06642eca2bb4e6c2dcc83c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab01fa29ae98ba2e68da4d3aeaf1766d8f2ef45075fa98af489b57d64b0d65fb43f638fce61fc05261f9f8c82ef0c17c2ab33fb841cd62e7c09b8f83364cfbfc7da11c2158456b8da0c815e955b1351daa1315b973d4fd0749e2d581f2e7a8ed28c9e0e235b92636f133463093d1b9f1c656db0fd43a3c502ed80833df4e39f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4be0175d1d4eaca96becea5367809ba3c2d34741c22793e49e6be235a82314526dea3e531d2ead4b7a756a99b07c025dbabc5574df35b9ea9a1af27b7a6b6582510564aa4daa5721eba8664792015eb71f77ce7a49972717f8a7a98ade7e5db033e5a31c52464d7eb7881f0bbde461b31511c5ef688be55f787c381e97b225d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6283d75abc30fef977dfa95015248187692481eb8f97dacb8b61b7bd4e01aebad14ea17efd340923208ad0c173141c8cbbe59a93bc8a3339d09f8598f196f6b5ee244858adb80b6caa07df265806e00f470e3c407bc726f5420d5688dcb13199f06c156e6942a02dac1b18d1674ce49954e59ae58aed6621b1b9a7f1bc204a46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9165bdd4428bcbdd8c4ce99ef98190563846f1bdc66b67062a910ebdff82ac71ab0cbf0adb427d34f99dd8dfdb310896faa2585b4960574bf70c14b8a6f3f3786a59fbc9e44bd544ce6b3f8433b6aa4f6901239e117f6db87934e41fa8a69f2833b7f73e41d13c7619f04872e1a7df2b03edbce5c5c6229de6f3e818b8dba937;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ed18926c19f05cd0d54bc9335ee5a1dc83e5a6477b2dbb58ef90923c2a411767bd0467cd4f8f2ac0e2a358cdb110cc0096c5c4d73b55e67a48bc86b41681ce883a4dd27b360610b269a2b236b16621f21446007e4fcd6038cb001b313c0e004285a97a999092f152ea690db4f6a5637c4d25ac1452f50beabee701a4f2ba3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b23f37e62b06a57368e88c1abc5b114b28939d188b3ed5bc8583ea61e0b5b6db276fce08988c9c078a8c7ab87512f7ba54b80b3c4a360f01f5e91a2cea32f8316428b28d369ac94109b50a675d2948fdfaa7b0115eddddedb5df3f4cab20e50265254f9ae70f876ddeaf53df405e4544ed817252e285a35d736ee2f17f5a609;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h493d6718c56c81184901727b01590934d33eb3c6c6b5e870ab452e5df68940a5d6407145230f753724ba09a132a03f018531d94bd801bc3b9c5e51742691d11bd45443b6db6db37b7fe1b9abe7f971d3adacb8103597ea86c41747d0a68a973b5ecfd2ca6700608ad3de8ffb5a1f48865b08c25f341c2b69e418e4df676e3308;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadba12c847e8481a70cafbe4a665f3c7370b3681a35956a0eb93cf09b20598b5f77b0230c539e780935befc85a069fbbaf773f4867a9837351756531d00b10e0c9eedf6d9b82f62c0f567d4bdda5f137f3c4ee11491c2601a8c1155a0a3ab7c22600bf00cc1ebf4e8a89ad84a02b0bae4356c557beedc2edb97ae0a9267a6bec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaf3dab8ac869f17e55fe4373d669b21ef33a941086e836f6fbc2adaa2a5e40cbc3963763e8da019e3d35ffdb2b31091ee060a8b19a838ab39eb83f5125288eb6fa59c7c77dba451b1f45d1dc3c420272933bf25565730113a0dcc8e22adbe25cba0d48f27e2ffdf58a5f1d6669791b9a12442a9946c404231b0a4d63e704247;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h255acdc11fd4a5fa3d4a86b9ccbf8eeedc68d56fc9bc4b10218ac64c306f5d9aecf0924872f3c9a01b603f22988b59965fa74b500d7b098b3f50c590975ee581b6d4820b2bb319db12e7058ca53e9a25c855804ecbef97cdfe25d66db4b5f5b47c1d799f01e5cc3d420e683c1d72db758186f2b0a682b3413a016c2c6315761b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a6b96a515cc1faa997448a0b8773416981e845439e62bc8370a48ae46c55c2500d3f69e868332e833b57f64831aa8a7cc767724c25a0bfdfeaeb4e4c7d696d7ba8c4c20265c8f3b9dce8b4f35a903235a4dff89b45dc8bb0fa7974f0fb9b647bb25fceba9c34592a40ef1535921dc6eec8985900457764c1d3a2ac2f793d6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d052c70d746e071c1c4b94a97d227acb8d8c5de9e2cc7a93cfdb85058721cae249eb5a22817c3df0e61ceea432d0c839f37dd79fe68d2d66db02ce3b8262f33e41c99db4666cf8d596474a6735f7e7d28d593f5b1273ca461e38f9e88df10493abf121c477cdc1e93746293c9a66455a61baa2bc26c6561ba53bc46f334764d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he383be3a2fe75b2c3ce5186fe0155a1ce7deccb47e58ab8392f621a005826cb7efcb7ddbf1ca6faf4d7e14064e0ed6c4083ced69599dff4f8012d548908d86932ada51e1cf00a38e34cdbe1f9fa190b7b3a16c0e7a0444efb16cfa610770a24e0490096fe5ef2c55b886de6b124d6fa238ca49741aaa81e2b122752cc6afd43e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1f0504062b128041a4851aeaa4310f00699d9e7ca12d7d15eb55f67d0f7d0cba2800b98cc4bd4922808fa56bc06ea9956df2cc4afc567923802bc614cc3bc545709f2c83f05fa437f0bfc71bccc131ce23a3c7283db0a0929f253493d308dcb25147a289beb953d7e7f31f20c015e1982c1e8b24fc0f6d4e9a566ee0a5b05e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55aa59164c9d7b5b5ac2175329c606e0e3170e00c8f677ef7ca215c1c4bf4f5d76be2c15730ee0d62fb3fcbfeb295b9b39833fae80f5a0b28f6e5ef69f78c1bc856a76a0ced9c649073ab5077e186cdf2fe954bdf1bf17ae8a2667c5cbce308ff55306aae7012ea96289f108318744b2fc20024a07368db266ebdab834b9bead;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3c274056f54989818f80381c642e1e95dd500f4d9c34318ca423ff79dfcd1d42851dc67c7e61f978f7bd9d2fae3319138551d42dc4c799feaa7c4398fcd6823bb1b4d1068f7fab0d600b6b6770619a45bfaf3bcbed7625c82b7cc884d86bc03ae11809ee6e186c4b9a27203309e8ccbc5adbb9f0b9f06bcdc92978dd460c7c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bf58384c9f80d0d4fdb637133f187d215eb1ab0ef2d8c5e46bb1cf5e556cded79ecf985d4b3995b22e3c2593b12b21d28a3ea41d7c568a6172b88ce8fff6958368238be1ce460a8855923b4879e75bed62a3b750659e82bd5e27efbcdf47fe5e8a5ceeddb66d9fd7f4355e36707bcb6ab81928a1da9c35be270a3c3f79e70a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69104bc9b2811d6a857781432a1cf2167316b1c246a9ba9cd04a059b0e1df313e3e7f6ae852aafa05bbf254af289e9f5df10a711d8696b78fd204feddb29e617de492ad15b95ded51b403b492ae65e5c9788f25fb27cdbe932b59772f6b3ab76ec9da8d49f2a37076bddb09f36f1b5541d6d54aa403c4588d5fbeebb6f31df6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc35811d46d8c31ded3d041143a8d611c6ab4f3b43f3db2c96a305326b58228bcaca62ef575fe6ddd4be3635dcf63a74d506f37fa6a5007b76ec44fa7dfbca6149bd0aadd6222475d7e3f2c5777a080609870387dad54a97e852cbd9baad4ed13ea5653247958d0bf4698659af41ea770bcc0f7f137a7e71057bf93e24e26e6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef79fbeb0f53f36c93d742adc42e37102c549ea5e015aa5e2742d33abe6e43b62e1134f8f89d7e4e6820a6ba100f13e559223c643680ffb51bba78671d59009539688d344f001cae00852af38daf988eb9816bc5e9d8f112bd01872484fc737cd201a5302bdd6c12284e0ca308c5f352385612cda076fe84893e75d711771c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f25fad59a2f4031dd8e5c1ee43222ec240df5c30103358c4354bfc0dc5b34faf5c8971ff604d7a3a10b192de7b936774a6de835539714666bf553fe392bf0729ce5ea6ec4818750866b5c976565fc49656824a9763d2f0613e4ead6b3e1f4630997d6b7ff155d840f0bcc0c855641ce1def9194545692b94dc9323a012901da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29ba065be2c57fefae46504828759a1f74da5c1fff60fea15e38cc0b95ba54f7dc65d0d410dddd4d2cf007a109bbe0fc8e5ecbc052fa73e3e0da60ccf8287d93628105ccd6a39efdbe5578f5c51bc930dfc5c8c53b6ad1bbee91452a15e020a3be4c5ec4fba6f2466ca216d41484d46aa4ace3a616c7f8a5499bf061714ddd36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2836f43ac6d065fe6084dd72581de8c8418edaaaef53a22fddebfc2d641964b5e1c75c8c365e8793727b7eb72f9dc657ed9690f040f293fb17e334140d5bb94ae3e1db447a2752f441e92d4b4588767c674d58a53134208a78cf2c40bebc9b8731d87bc0dfc59e156cff438103fa4b71a43e76463a192245170af79b3fe28dbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e43c2fed327f33e3f74642a1e362223dc9b615b6ac9c138eb851069412dd4404d5e37bb85d4d9ef7ee837f3d4c755d940f6ad072e8d6ef54b723228c901f28ee4f2c3780c43198dec031d3e3de77e398cbe6676dfb1e215e3d1d8ebe4aea1d3bc5e6ee331da62b7b2e3ffdc93630893230a20983ec14071713641670c3afa36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2b815622028de41c5e61daf7dd19607f38469b3d76429fbb65595e741192b3f5f7e15e5364f92567810dd006d1be301fea9846f4599251d3e5bda0f7d51d8611f90c448292cfb684849adf0350af2a015ccebcfdcbb791d05d350479b00557b63d3969de646b25c85faf6d204c226256f2d4d0a2e8a2d0f87d6594f16507e88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9d4c00a6cb83fffa190426a37ac265ae46e6e7de253f22cbaa2fd563107fd8f188bb6e70cb09605478954021014489070ba643ed2d9b6694047778796af595d9c1364d7eeb98bf19ae39db7e17ba57d1f284cefbe0f4ebddb24913ba3e64e2526fa93f37a97cea0324d51353f61b9952921bad3ef1556090a4577b7be82870;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cae43fbc6ee81b7897f8d8743bc713d6268d597894b46feb10273453090a69776dbc9b61cb5a92b798e7f0e0e20d8e77f83ace4066e8528bd7db1705ee1e09548e945c487687112ea3ed02b0c0cbdbea41edb99a85242260e8c32898b05abe452d7a2abd5e5e70a6337f5ec00026e5036213e7a5e923cfe68e45472bdbbc8de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26213d858ed9334293f015ffec0f4ba047856273b81a5fc13ef7088071adb5d204037d51a25a6d966406c1e42d0a991543ed3a682e7a18ff3403d879a757d6587d98bf6113bf6f9bddd3454b1a0d6ade927681d64392a8b8e6d7a67a5e33ade947db9b59a28244c778d29b2aebed7506759242bb36da5de5361382707f824999;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdc42d4b02d19c3ee6ac045d8c61bed3b1774ef525668f67a216682b844141b08542b8bb45b62e8b2146e97c2e43571e3e1cc2be0c41d2be436ac2dcf1076c4c69d9519040c828d75af3eda792ecc4358042a1e231c80206c0866c34085532844b28d51e0cd84de70031224d6640964b09afb236d45a11547415bce0a6cae313;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he009a856ae89040d15adff947b6d110103d7563b574d924fad343b17324e6042216de827b33cdbc41c6de4094079ab3d0def42a18008e1b9b0d62dbc0664185b0fed714f65e8892e2f64dfbf41954a0986b802fb6d80ae6b10f444585532d0aac0af40bbe34e46c5b4e499d21900620429a8bcc65545d5620953d34d7d5c0aeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80a3cb5659e8a6bb3f2fe805137b0af31d05423446bbeb3285394d1e041f5019d0ea473e7904cad0972ab8a1efdeaec456159d942efb38852dc49a721ba2f91507e04d7c7fdc9caba478a72d5cf5ef5be9a579322d42d07fea614d10f4f2ec27e2cb2bfaf20c0191a0dfecef3fae6937d26cd616d0e78095c21472a5f688ac58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ce819aedf6e83d36cf5e01daa296aee79214bde2e96cb72f30a028dcd28f6584c05209fa06e81432e4ca01b8bff9494077431eda800b4d871f84f0719acda768c3c96ddc6af097cd77656135cb4d9e4064ff87d2baecefdbc7ce022efa232f33b7b19f4d0745d9abb1c36c4d6c1b52d28c739ec00cce85c5e702c7c66b4b167;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b03d970f49897280e23c13537b80186b4638aac7bb5c8f3bfe45af143caf8c96773b5146cc1a3a1871486e8c3d5a8a3d50a15965a5181aaac85fe32d7267f82faf6f21a70624d376845d91f0bb374b4b35b2112a0acd7f6cfdac262f1fdbf301390c72f96f6b2cdf888e9a981f3f860fcb8f35a58c50cc92d77bf7b40807e3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b5ca6c6286f43ca5790aba926a2e133b7d30a97aec7ba253a609c5cf0109dc00a8017596cfcc4af41ccb56d7a2765d48773ead6560f6f0c0b9c10d8fcb20c7b1672565b221b2e1615da2985153218203e2f111d6766018394a86fd34661761d02fca04f294409e66a718f36befb9a24a1250523a8197330bbbbfffe3efc1857;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a20e0f1b8ead04e4583c1249f5eedbc609b284ab60e8853ecba4197fb4e996c2479dc0e0d38e3c9e9d32834556ef66079593b97dc77d2a9c0c77a17ca915b405d508af80c9d1cf63e3e80ae6d5dde0efa6be0bf4681442235f31b9ab1f51940bc23cc2356a3ccffc841b71a80503a107c4d8713bd4e320e9fea01ddf1137f6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfbde849f3c2900e148c986f08b11445fc12853fac851185326e01191720289c79b735d21166c21f7a46e067c9ba16808fe1c8b2d3ca0308a275a397ec9940aeb7bc4434b107c12d63d630490729530d1a626ed517cef83cae973a5321fbc1c6e9394cb7163d4a4018510d7049566e532ab737ba0edc7e964e60094d2e3dfdd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10ba2fb6be8a022ce6c7aa046ad27d668d2305cd0bf84093d1488ab79caf7166d22471f97996355a97371c1ffe8f4e323e2a7caeaf97feebfa8cd1d6655c171abf52cf1e4bd84c00c32213ef53d88443a3d0b708e01635368cb3e3eb0c63586875f36b61692269b7726962696073c3f89ab4b8f596e6152ec842dd9408efe1ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23a5b463b9d8bcd907e5c465cebd5ab86c0095d2d6705c166baa794df220cba3bc44a4a29e938e0f387b2d29655a482fb7c4d6823641e85f658d308c754b1bbf566f2a787a95d76be126efe1d87bf52df090de26876866af50e3c7f8781623c45800a50371c79de47caea7e98dc064951999981090b8d78308d67cbb11025992;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69a6693861eb69b1d78ed7b5b48f8cf9e83b91b821eb681480b8826b0d4eba441fbe6f52373183e34199bd75a9c9cdc1ce82b41f3641321ef02d86cfd9dda4b6a33a4c679a99a8d8e21b8581495269e003b4025236210e6da583f68d1d53ed2efaf318171403afc1859ce50f56935d1b334cbae9e736a2d3bfafd2286e379cc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h105c90ed2ffffcaa963a0e4f5ee99068778125490b46f452e3e7ba0a1f29eace216bfe5b161633c18bc3d35d07897a349ddcc2364f8a80695a0fdbbb4372f7321455c3746776cf606cc4a0be48c8884b3b2890e4c25e06f11bf14b6e9c07a30d30f1ee47cf4dd34aa0091427cc1ded2e29fe3efdf25ee1a4785d2b80f1ef0f75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50329a46071bf63fe339232844f7a20beee0060e5b613600a9acb1c414b12cfcbfa0e3f4bfa8a6ea9d6ecfb04db56d6ee70a3fa773aae4f15325885eda5839723f265109adc03845943375958731b87d253ea8ec34855abc4bfc03128d5d0ceb5223b3fb63e66411f3705b67d834c842d70e1f6ce8d6cb0b11dcfc687a318d3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61a1bf4810529a4607ac07328aaf36db0cf79610e556148c9e2061a65cf962502eb597daece0104f09d71e87a2b0f176ef34a1d8f1a1da66d2eb7d029ac3c0f40eb532abffc2ea528e68730c9c6a8b4a7ed15f3a76ee380ff5d0bfd6ca41a857e2c98e8f2204ed85585ec8f8b8e50ac0f606eef84f229e811c2b31a3062294fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h360e4f39e6e2cc1bd80600823c60fdcaa94e3cf170d2d92f5d24315b093bb5eac2dab63d6357fc180ee1432227fa343a5550eb4c7ef01666f0e3c8d6e7205e936b9c536f70407a41b833c5b45fdac611d2923d3f8cdf0e3ad6e1642171bfe16870a8bc0775a098f1d3ac936be0afcc1514d890b630969cf6d15e2e4be0d3613e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc631a361606b8b6c4d12d6bb62f63426d8ea3224a103c7163479885a438a4b190fba6931a89c51033ef53968bcf1796bf4955e86b7648613171d5ef6d71e8221d235e21562a5e46f338f5d1175102d15171c7be541397b27afa53a2147b5d6c5cb377a5ec635d195978685f1655b3dcd159f2539ef4ed259eef27b47d99071b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h117b8b12336a8f6ce0172f36957ea8db5b11f6b91d07a02814097f7afe1b929d6eeee68ca3159a23ece77e7e133a313d9f99d319ba94ffdaac5a9c9012332a69c2a0b20225f652ad4f004969e987688e4dfa698a06e576c6cfb476a25b4ec868c1442f6108bb3b4419b4a1832da27e8c5250abe0f577f5c360f8b8c81ce7abb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedf148e86f79149a04382f1e3cf880d47de6215d7cb6524c9546627d0e2a843334b587fc5a96229e65d2917c526caf034d6e51d26324090cd7608894b32d3126b31b3a071d99090f5aa2a44924988165068883d62637a25e6adaac2d7e1932bc4154112706a658a93b8f93c4beabaa2daf2c1412ab171bee87f0491bf6787028;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h372348433b1efbe5bbd92e4c9f87cb575032c55c80ba69613ac3dfb93720d8c35a1f5aecd510a1cee8f6129a06b1be9f040bc04884750ff74c1d6c5e0206803c0080a360bbbbb188f37d254d8036f22d3f19e462fc6f56d1d2f88830ccd41227121b750a0ab17a1619dd37a891b95647e78b39ad3d1c50c1405bab1f3644cc5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd2dbe652de275a29896265d5aef5ac58cb94f06415916fefce57d087de7e2a935bc7a98c8ce5c69ad55d602b965b3be71d67fb323803a985c15dd8b67d01b5fb3869b72e782e4446e2758c69e8ddf3a1be0175136ac640ad90bb12dbfc992fa372c0268a8801fb33d54877df783612137d0a96f27ccb9283d03c3b1a31da3a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45f37538b951556cb03392f3554c414b68efd4fc8b0ebf0d380acf84d5ed1f290c6186fa7a6cf026d66b10b0c4de1a0b5e0d276a62c30859ec545cd9c4f28da5edf827364aded6576b145c7bbe8b93b9d1908f248e9f55b10c822ccdebc875502b8d82717710162f0b06e14ce1f90f8c22c00b7b04c76226ae513c151e94cb50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55ff97bf41c1d0112df65817fe177be801032d70ce547522f8323a4fdf12e0b3edd6a7accc1e38949c7514e823f03c3507b475a740e28b997e8583d4e498594360cb4969d7d9d9024b399a08b3db0eae11ffd150484734f109afb47f5a7f7eb6730447f4198acb8f1acc4f77a8a6497324dfe02cb7699a215ed90f011ccd57df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb37ebf73435c3bff74d29d65f8a048c2983122644a2e62534e521d79efbb53a919f247f922ee6b013d0dc8d47b86d763a44df1940cfdbc376c3aab4c4c4d9241e5d5252ac858d589abe14cddfa14cc7a24ff04fe1ed07c04e8832a80a75081fa40406968af365ffd92adf5c97535e30731e2ca1138804c874697fdde7e147828;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37ebf067215ecbf06353e55e92c332a1633f8369876396452fab5f10dea055d71afe3a9f91d0e5f0c8b317896364e3c0db1f15e263a1fc7bb67c0e7074c7a6fb55332097d65416c1f22a318667bab7cb64e25b7852b0a8d9298367920f4384e44c2546a59359e9abcf657e5e2772018f0dd625f93686239000042d2d66c76470;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4ceba72d347afd66f07a7a5a567c3b3620d4877e7ba8515414576d5c3e826eb7fafa6d57a7afe95983506609eed7270b26410344711cb0a2d146784d6065a9497155ed77ad34e1f09c9e14f0d3c4499993fb294a07ea3c77b058d27f215611296e6eed61a9ab10cc26f4433f4d3d1c2d3fbc7181a6109a1c1bf69c2d99b5fbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce72b037928d212c876ec5d189ae34e161e3583758e7bc01a3a5fa6f49e4f4ce5bb4e8165b01d8c3a0355b958f18d9cf47caee35b4a42ef79225c4667d369cef8276fbad6362c7a188f47b24acd56c72846baa8b31950ee9108f0ec4b6d4451b7d951375856493468f58bcc2a593e194615c53735482a2d43a6c3763ea2905ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h173b935bd7551481fdab57996b641477b6251e5b66035fdd5d0f6baece66a2ac3a04189bae46f154d627f7f566a904c596c605803f8c70b01b8269172e548cbe331fd3c3e812c7a0f091ff07f48cb4fa177aaf98d8d754f6db6e2df37d201dd9ac7e183bb2128b3bcfcc5ffade9f693a0a4d6226f42d4796fd2a195b3dc7aeee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d2516917b4ab4c9b3d8d981cb935ebd0657fef913d36cc87db638fd9fe4ef938a7be7f51f8b0786b89c44d1bf9f71e30f556df45280cb220965b30da0cd2fe9cc542cd8adc84d1a87ea1bae5b5c0625624ee62c462c9629a59b2385f8172a3f0d018270d4f916398740552dcc6dbff8f19409e2919e46c4c4bdd2c15ab35ae1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2aef9ed759b7a034a75402480f99c0905d92acc40aa59cda9f3764be12b37c3badbe03a8108fc52d84f81308f2df0771a0bd98ba7676398a1c82110468e641392d4dff53e4e8fe67f284649223ac835e11703ac31ec04f46e2f74c09904b7f3f241b9a8136b28c091abe0e8459d9832c1edf72f6e66ad1d7b6765c84bc5e47c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1b3b3a75529ac1e22068d6dc384da99de9b98456b5c4a76c7f6bcea52f849b2de5f1fac5103c5006e18a658b89c8b1ffb3c3822510c45b0e10a284f06062150fedecf9968f4183f0f3e9c7e389eb522671f75a4811ab26d90fe516695f3bfed84a4a0415e0dbecb09488a099190665ab1dd3300d26737d1d17536f0470e7f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h744235f997218242ed800b8927fbfc97071e6da54dff23f3483ef8b8665b6b5d44879582fc0856566fe7fc05db6f1414117099c36e181a5f03dea160580df448322d696fe33188359abb5781e483ec69305163999dc0fc5a8e5a75f4a7d71328cbb33a01dd5fab8af830a77fdeb9ee45c453e87b647f88ce8b810d7cf80afd5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h424b4969112b6d7b9b6a843707471dd770887df4dad31165d1b21f1f30165a5320cbd44bdd8312664d0a548350a67463d8f4c9d057d317e245f2cd7d244b478348069b33ad3563c5aac8c9c9d233b985395def74f63ddcb52387b87bb0cf7748fe5c54fd775536a671be99b7a1b0d880e16365c4c10b30bef81294fe96e741e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f54e24baf9eb30f3074aa9da2ee5a835c4fb545e4ab6e6b82249ef2566ed68ac5136a7bc3701327191062601b6e1707598ec518a36a297c626ca9ffd994a4e431d44fcf6d04324a88a50e03c7e34e0ed721e4280b78f55566e3b123653a77ee6230025aa84bceca94b4e5b7718c538ab1a5bbc6cde55ec9508187de3a9567e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce9f7d06e4ec5dcef695efa6b83f6052e7dd1f3707d9a6ee04119d82b4f09e67751bc3185680f48847b29f15fc396d7d37d1cce285a7ba2636af0072b912d462edace545e8b24e471cb6c4a03b8bf81cb323345afa18aa834bf4d35912a7d015621fa49f26d736e5b16f32c9e326aaddef22ceb85301b713de8e54062f3de982;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6c420c2ec15e435cc41a985ff772ff782c429ad5095eaba2b9748c0e3de5aec5b55c8180b39443051fcf6ec92c7a6294542af85b3c57120367dfa7d0218c5b96baaf19208d313cc623f4ae6e1ec34bc02aec3e9008111dc5f325ee936ed5d2934222d630b275f4e2343bebf4abd0d44824d95bb1dea3ff24b03241188281c9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8060abaff1d4b3ae3e6f54b537cc005c799613c316d1af2ffd2d3988cdd6dbb73cc66d4e6bc7b0769ee81c029fa25a4f950b00cb373b10cb9ccc29ea2bece1e916dd48ba8882340adc3522dc1e3077b097285b4766da845d8e74fafc95e16669c3ae43bb873d2678f540b2eb595028ece76894df1fa626315d3f9f358b5be667;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15f873c704a2928354458b2630f8412dfe92f6c4214cd4c9a246015288fa97ace4df9dacac1378311301fccd5cda1fdaf31a77211294cefec63153ce084ba881d9232b546f7295f3fd98c554d78d7dcf79446228a070db4f50627e67b76583e4a6a40a6e9b9e4ee378207858103faf1b80a8588c9b4092c8ed411407118a4c9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1254515a839df43702917e730d444456e9e60cd5c5ef244f7497948f7d40a103a854b5d5a2b3886dda211b3c0d61ed798079417e4d70cb1ebdb133793cc495680e4f91246e991b2b4dd75708988c3faeec4715ab36c9edf4a1b0d01b5d1e50f8b56e8982f12cf9ac76eb7c58288ba3a7b59ab1642362a757ba7b2e481da68eee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h449c0e1c2ea6933699944c352648368abd4f98c4a25dd5a8ff5c498f321d77c923515b1c6868c1978342e5733584b17421bc1c6c2810a7ca25236394fc0661f53bd96629e4d312ba4dc61a76342f6babc01bfb3d151327e92802ad11833cf2e9af8a15f038565f545071df01a59530ce3039d702fe34860b530582edcda579a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc626e54c75e284ba0d271e978f24cd42b3b3978b1995ad763329b4ce0a316633015ff8fcff8225228e54851b73bc05e2f072e62a91e292cea4d6e3a92ad7d6f874ee4ba26caf19f0bd5a57eab357f6bf94bf49e256c7517f875d9cb63f8a5bef42251dbdfa357349d4969a8a16ce2472b5c8b8168d776ca8d9dd14d21e2fadf6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0411027def644269f5b4f87b07c1428e8868f2f0bc8c3f0475f18ff7402aa06bf7f0f636c4b2df343ac468c8bddff24ed8eef2792991b29d33a7ef21541c28fc1880980da5de74bcc741f3b5e2bdce60f24284019a50649466488ddaad6019f820d0df313f9e75a92a55d21cd71d9791417197fe6e5d78693d4ed1fa791e00b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69c7a37feb27d828d5b44ae29332a8bba4b159ea96528c1a6cc0d5890d49f27a69c9e6c22e6024fb6e8e3a50b2c3f5e05a7462ec96a5d79b33a735363bd93f303c4199fd767ae00e48f9726e9eaae0b9bc221d5d342395c9129cfe4c4ecb864d3993689248e82ddb7abce38a235cb775c4689ade724e7d0574a557ac3920ee38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4046f67f418ce27be6d1711586c40ff7e5ad15149c740ed5b8b572d0cc28a4ea792a5376a660ffd4a846702a1b96c567e1c06bb37323d7b46e98b63e59b042595320f8810bc28ed4094e6770a70cd2c0a480bcc3be06e3a8e800f7ba0b7c8316fdacf4ff5ddce436d3673486e909e138b67ef2972343bfabc68140d187cb0903;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1018b13e5af53d0e9fe8368e7157caffaad7734e0fc2b12c657167bffd19fab58024ed5defa1979ae0c01c48e50afbfdddd76224973731ef9d57841f1ca8bce5a886404e8750ad3aef0ce794bc3da1fa48ef9e378c05e7b005dc41146ffa4ddecc54eb295c5bd245d2d22a3bcb52fd45f083d08654040bc8618d49f81712cd3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae6819977857711b55a9823d9d94c819f3000aa130c88d765446cbdb9f748348df5c5f5d304fa31ba836ffa647ba8b1b2cb984d3fb2c1c74d2346d7c6848005967f863259835ef9a845c97bd93d8e5d1acbb5ca0d3888ffbd224b31fd2086629de510b9ac524d621301f2916731a017342c732d188756f10bc7109bcaf773a81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82aec105fa5696490a910f2a8e2c3bb127728ee07010104e86cc62f92fe3628f894b41a0e2df150ce25e196fb0a660c95c04f94ad62353e0cce61781cdbc20037efe6a47454a0e7cfd5133bdde3d4c5d56f9b406351ded8e770c5db51713bfb7f1b8919ae9f6d282eecbaaf6ca7470520fbb916358f282adc8b0489d323583d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had8acfddf65b0f81c608c4dd7647920d2dae281396ab22454e79088f5708cda069dbbe9abf8ae04941337a997e91ad6aaf39cb2d1200aa15153568386cdfbb0a873235bc63d54e296bb2842b2e83857fa90e5efcc18d95faf9fb5984b0aaf074322b62badbd6d8997bd3573d91e91000ee6a2e011650205c6024f005e21a785e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b9b489033acf2b2e666df299fb5f6bb74adde7c74f305ae830943c552a20ab1906ff7bd160deec83d9b2e1c6245c4d4732ccf9dfe1028736f46b4576e0c8263d976326eff8571b46bc924c8c034a011e3731defed7411712633495a3c3ddbaaf445a78d77893b28446fe222fb82b90879ad77d8eb0dce8a9e6aa43fd36ac772;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b1be0040d14033af0fdbb59e84834acebf9390509cfabba8c5b190ac981bd5a9d164980096f9195b7052aaa454a466c4d7f73693cc43319b5fdd1c128e7aee676ed5a8a040f36867fa69af04057d2f048777922de9f9317247ca1261a77051017ca737f4141fdf0e565a4996f098ea6d78bd835c43d39bb44cfa75f54531218;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56a4e45b53644c101bf3c7061ba5d85c551bd35a6bac2a00f3dcbc04a87cc844442345aa8ef4c114a125221007b7e2adf0df8458df2b0318bc36224628002ec4d62e3e31e3710d4872f9e0533c6f9fab3931d7a31ded91f3fa39c566e21dd911e290ec81a5680f5edc102d629cedb2c305c46b4a41330b58f8a8e113f92efd06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha08f3c470339754fcaf50142b48ecb48101b7fc37b17f78a0fcb2fdaa82e5f4e855f7e0614aa4ced2a255b895e8afd45ce635a4c97920c12f7ae76b93195e3f323416e9eece2f289e75ed90f157248e09b5b66983a2bf68ea551dd2c057911bba86cb807a59384bd14ff1dfaee407a6b71793161821f8a9762189294ea624de4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haafa22fca3f39c561af1bf05a0b95052f720e4ead029a1f1de92996f595fbfe7630a6514d64facf5cf1b21e850892eef5928957266734564750c46784f58a538be7b3af941585086d29e8afb44ce578b12db1f2750846dc1d18cb0555b922606de52839feb03ec5ea27738a75a2464a3a607e4d06c32125ed41b9f4f073ab0d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha002e6e8676f9c18004b861dfbd9cf7daeb90fa3b514c20af35d9c7e128e5b2afb8c47a0a8ab1f2c097995c5397713f76201abf1c5f3ed82952668c2b2024a0840c02fc7a3d6483597e4e8e869d17f6093c800f688110e0e6582561fdc034cd1fd900c052533a690f8987dbeb784c72b4df802f8ca358ecd49f81fa60fbc19d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2abc47e51563ac900825ee978ac67d1c2bbc0b64b3a5904fedadb85740bf6e1f2133ca23227bc446026d94e065e49211814ef4244502b5e846b9632a7b0267087acb87dc8394bcd1d18e55b8bc09d2b89ca79988d1021ca6f7e2cbaa81fa35119129d6507abc2e7ec08c8a9c8c3e2fd07f39cb9219d629ed8cbe481ca86404d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c9f0a672ce56218c2375933b8fce9ea2b6c6ed8dddf45046f8faaecd79a81b4316f6f16f07387fe86007d4433f8349f28a5349a46e1b6668a03c78a1698c0f9839d32ff96110971aacf524392826fa76371907603e7ff87e99ae216e85499e13e7e7d690b667fe9454461e0f7b58817195c7855ae2954e153d8fb926640fecd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7b3217d1861af8dfb934a55477d71bdc4db26acaea8685086f7222ff8e9e395f3026613f39271fcd4c741bfcfbf4465846c833cdc1a96a92c30c44ef1076b1db2095b8eace55fa785f4f910c41e7aacef0f45e29ec93854cfaffd9c6c5cde9a50078e26d322a933ab86d806fe482f89bec6a8fc648d169bca7a3adb1310d3a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62b17fdf9ee6fb6a528f2dd48d42a31d9c7bfe6c51739cd26ec43e75d1e37b574c182c2a779f88a996af02904d0dff1efb6c1495b1ba1955949f866522ea93d7c82b818c658d3e3b06cd2cedf5f67db8a692559e98dd992d3df95614db6594395c876ccede62a53c4a9a1364f94e4eb385ac037b5921079dfba3ef28b846eac7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h743297edef1dd768b0f56be4cbb600fe4d34c752331bd6121313fee5c3536c5d899d8ba41ad78b016ccd01a705be5d97a52888a1f71e99ea6e426fd6b16caa6030f6265bbca5a5c614d7463cac1c1401d5d5c353d0510e087a23a1ecc9dc87cf203d76c39b5b0cba1edc9bf9fd6252b9106b66b505b6d0b6d7559f6e2d582a6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h299d7e8c64914a74148459d8ac9d0867c76784159c9085b5058fbe23aeae4ff818589c21faa2727bdb86ef2a4c17c6fa6bf538f4a887c7948d20db90391472b58dfd3f4c38c159e7f2b43ad0a5cac4b88514e1b8f141d46b8d2f6152235a0e9afa5ec27c031165c35166ae81c86a74d28064d5a3ace83079dc4dccff7b1f1a17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fd749059239d4dbaddf25fbcef1ce05504af36fcf38b89ec302507c22f46f78856498edfcc6d9559d68e0d8538f5d1c448acbf68ee21f710d91e911c5498e55fd47efa4df7a34c471a6f4b7f56c1ceab33d5cc7cd0a7c881d45b002157f83fc21395706dc9010b577ce732c998056404d00614a13ea5d07b8a105af487b6220;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ae588fd7cd95e8c583ebb8cb1a8260ed50c349647aa67422816f3e1a7a83247c331cbf299e47c0a7d0b34416a7b9162bdfa5cffeba82bb021b8ae1888e0df6d6d324a1aa1254f7e945c498645327ccafc03e23f55fcc99c65c462337bbc1e5d88b8b923fe81edfb38cf535e6914ba5a3e26b0542d81f6fe0b12b4f015104a9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h531aba5789e6a328afd9c69525738bd5c960b772c3b157db1fa1caf3acf4d70e13345465c76adfb385a7308855d34f33949cfe105f032dc7e0292fde52ac19b393aed8fbe80bdcefcbeb949eef9fbf53e835c30e5165c32e5f5dc254c2b88e5f0a8a9f1ab37693e53b8b095d5e56a144281602da6b5ddb98330764bfb9169e64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dce83f4e6d33dbe3d9108cc326cbd44b7c2eac14066bd42b939343a1da0b6212327d2ea7550b7b21ba6169aec69e1a20f1349a06acdc35a4eaf77f417472cf85f3a13bc40982652ac33ea82265e0dd3f20ac47a33a655beecc760d857246acc6177d3d97ac2e8b4d779f72aba560e041ab1cc6f724a6a9bcea83f9977e89608;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56c46b0a7f825d48dcd2dcb206d0d6bf9a09bf87d39d0ea5372e24aee4078e1474c44a8e7f6dc019a985d8ec0c23ef4a417ce9e04a375b4e93a60367f63236bc0e7ccd9462f1e4d5432b531fbf9ea37a48fe659681a9169c9cd52c6f09ea1b3067d5c36341dc0a6147c2fa46020207378d6620aff2ee70019e5bd64592bdf9c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8d580f11ba533b9b1866b0b2639ef93051a09ac1b2e37d77c83def6c92c24818c47f64b4f4a78dd7e0f311be3cfa36ebfaf8a2b4dad28d66c3a02e13335311092a8304cbe768db58ee7934fe8b5125a84810a0cdaea73a42fdeb423d86d87596a43d8784375a72a406615d4354a41f537789e62034043c16f8cd859920551cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9b705f8e604f099c03a64d6d96bc0b37e602226da70f4448c4e860d795aa43671ac77c0930a4d317a243001099ad931194192cfe3e8235b6bdf063f82ad5c9694877aea0f05048896b96ebcca667ada74a6c4a7abee1091e689d43c920c49b7228b503d14bfe805c45158285b96384da520863be738ad84eb0f21ab8724b2ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2614a0f19c9e5786a39f31810ca24e9e7699491d079985fc72fa3135044fd4d552def4dc628ef47ee15c1dcd7fbf6a0d497fbc38cf5f54d523597372a03df5365d48489b755ca7bfe0ece32770158684c83893ddcc901a71224cd330d1562503a362672777935a9d917c0515b39dc2374d967659dc066713d08b00b381ba98b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha658a1a1524577ea481dc503646f979ab3a6fa352518cc6348902ba940cb825ed0c7e2d0ede0ec7d00d25377f25a08bde6f316281d6764cd061b805048c3a1259eeb2c7af07e987a122488e57c5d5eba60bcc610366378855d6556ebba71a6765d71658fae0148ccdce6874dcc17fb1c6d72c8cd85d40ce0efa972e2e9a20564;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd77294cec2e33a9569556c920b167331596fee1c058d4a32c3da5ca8da9fd8590f25a680a0452ec67b0a65f9a30005df5c6c9e0906e09c7d877444274e3fb772d4d41989e286c51f9b663b683554ef1c331eb3adcf42e76cdb6cba43ac0330ef797879224809fdb190aee74b76d587f9b57a54f3d420ee89a4d7c3fc5804491a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6fbbd58ca370a3e6c1c0d4dd84d1a4fe4139996002314942a064c917ce08c609b59b9f239bcc3b644e29ebf3089cad80576e82c0e478857558bd77b844784a36480cff8a07eace9c0547f020cf355d327b83f699781e4d11a971fa2c8e0e4172f5cc3de88f24b91dfa66592c3b209582b7b03215f84ff996aba43c51c1a470b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91dad67768c72a59db969f9cce455c56467635c1b7033523a2929eae7bdb588501d6da1d3d7a1c043013d3348792d03c71db3fac43cd95b61e4405b6a4fddb2d4243f79ced0a04af6889824e6b884712b3af587845d02096abac5b13c911e9cb1e2bbf6607cf3d651524cc3c997136c9effb18fa756baade2667f39f1f611d37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf73ff44cfd644cf12195baf5cfda03486c2c0914ec524ee8c6b404f6875d1c553bea4700a00235d205988b1d0970b2440bf9bc92c34776096b65d5fdefcb3d67fb68321847ce30bbfe8817ba3c97dc945faf0c6edf02eb7b8724ec78dd4ca1b0b4f7502b0bbf0e664a1b90ad19682f4e0e7b724e60132934d46a93d4a89a45cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc84efdcd12423a6162df43742c51acbfd1d4e33fe8ae69a7f8f4d82b9fad90c496f799ffe7f96da2f09862ec2bea7755635dc6fbd7b5441b787418e3ed8a89075a962ee58665bb9a53ec2844f3b70ae51c5de346982154b222769d8c9cf26184b78bb1013e5096660530e1860e09a8e35b00741b2593a3abde440f42a789a5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e623dccffdb0a77250ddb3320c4f27569349e7ef4be4cbe9f93fda5cb22f0442393c626c8ef771b4089ab4f486821ec97bde2903f2b014f5825518404613f3d53e04a5047435d719fb298e112b33d90a05279f91cdab8fe19c912ba3be1dec96fa2ea6e8297bf54251712f4708e9685aea5743bfeef08b3b17ec7d8e746ada0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5301acd8397556a710de05e189272e67142fdc3528e99ad8fa14cb4980afbf19796f0f4046e4d2d5b90ef875d675d0ead65c0d96f4c5f4adc8810170aa534434d0a71117957a7716991f41832ae2118af543b7e355414b644a9fd9be92fc4ab89f98db1cef6d3393057947b1bc871d18ed54e92b1a47bbad0f5979856fba6e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff5aae813379cb755ac45cd0b37e9cf693d8d2513a240b18209eda2dc77a80c11304266ff21e8b9b4c049f4570c445de0a1c84b006a0f2ef9c53ea342ec82f7cd96eca9e09c32abdc835741be15984afc5761051c068cc8608fb95bdc22411fcb00a79c6dd85e943bab51f7490107c5746ec9a02ba4dbbd7e176b6806d46529f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf01aa342d891c193b4226abdf3868014b9d1c7bcd9fee783fdac41d9a208362232576cf556f3dd7970c68579726991e491edecedd7b7a83b12534a9a29a7989b9ecc975a636b972860e81028db3adf2a719579fee4b0a48aed1987f0fe8f8a9ac67a89e2703d6263e99cf3f480a4395d18392dbaaa669c4f2a13b308f53485ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2beb736fb38c53c7ad18fe3ed5d1a7e0982c9a511b12132cfcbb5190a49b8a51e75523175c65142fc236fe8e91f0778c3e0ee714147a60dc2f59c1a3ae5de6351932a5edb3f5b26996ab7dda00b12b08b01372a0829c283ed5bfe13183b1349a675863d79c0d0e0b433d9fb95b5a32d857cd644dc2f42ac353aab15931d08521;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c69349c38be7c716a9dc7de648ab64fc0bef049a96806b9d1ee6e2739d03b7f1539efa5b9bdfead831c713ce541e3d164c872fd6f49bdd581e529fa9743a7288d7138f3efdf39261b06418806273f667484c1862657dc90c20be9876b13fb7710a98379dfc21c163265678ca52ac3b1df3ff2aa44ba546303cbc558bdeca56e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c03b132e86697ac4d8c3d62375cdeb37f1fd7d0690d889556b9773364274f035cf933fec6d875dfbe37a602705b32f0de5d600de9f005049d2cdddea81eaa4d9705469bd87f76bac028d5f98d552f5b2b6991d07372a7ee88cd645afdb3d16d53558b50c2f0ac51039e06d1ba6876a16d8cabd16a0aaa220c002b23a21a2896;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57506d221ebb5d251c3030d4fcdda5aab02b1ec52d6965a414dccdda82bbd42db15048cbad53c96f80fca336a23eee0075a442f02797087ce90ec3203c91b829c35d68bb47552b1fb660e03291baebd918fb1ddb639a1a4b95c2b554087ce1bea6acdc3f86947be8209b7b76a8bcf7e024ea205559680a956b73d2885944eb87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c71c9fabe4ee8c7bff01cd5f4476aa7c36127e5c22d76a0688e258554e4e18855259cdd09f93080a86afb983ba835f38f00d8307f5d49bd36251fff7d4553cfe7efea72a669a3e0016997af058c50504c570528cad52087e9f474e406c1e4904bd913ee0a85ff36648bc93157d2bcddc28d0b8cfaefcf2ae68af0250f2bed74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7213d50758bc0cf40389e96c17f10de142e68fe5972e6bf12ed9ba483f9634814e820c6e687e7b7e6f6645d8572d77b54218b0d0569e744f036b647962498eb67abe959b7bd3676f44d7982d6d763ffe6d43a5724ef2d8abadc46a11db9eff2b9a94d11fd640eba77864674f2ad94b9db728befd53aeb0cca5c7f4f3d2d87d41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cde78efaa0d73f7d059a93d52cebab977d55f72c3b8a4e7711991b941b08a3eb59bb8b5f63102d98beab0e2bd1720acc74ac0da4fd7fd5856f97411f2a981caa9a71a73976f4d3dca8f92f1a40af8d301b4b4e288acfb7393e328d7e9375e34a800aba31c055ce2814a67f2a44501a9d5730d691b4ffc039111bf6b9279e62e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf5c6c66755d6944c725eeb8208d30a35bb80098ef728f91dc6798fd097232f10e3fc77d5b8361e0de0411af20f868fd1c70c5c899588025bcedddddfce1f9091390e647465c72c774e1281316ad774538261cdc24f0c7ecc6ce779e37e51bd009ac792880a79e4bbef3f31e819142e01eb9b5836ce24a1686d6bfd4df791c84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed4f0f5d51ec9fadcb90d91ae2ac17e635a5f3d634ac96b50ab781f585d3155b608d5046c55d6d42ca1279e3ea517556eccb513818fda475cc6c68430613f1bc59f6627aeea3f1d542dfc35d0722b843d93817720b70d9c26522ded94675ca0988474b8755c00094e3aabad8c001d130540e07fb328f5e9f93f6f565541536dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b7e6d921082a3248c1a04d58d53e8c8f9366f07738efd3f20203ac8e3cfef463e0c719f271595b121898e7ba4daf5220e72c7d3a89660dfb7c47781c9c615ad963fc550cf9ba14bf9adf15b89fcc2e73668560e3bd3e2fd9ebf91c03050a7e744167afb383a9128fe1951b7e98334dcbc235e9528b2855939a4a2884d7d0125;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a1c29fbe9bda58321c513acb867521546b09da4e3dde1b226cd17811a24e7457d5a1ed1563d9e9710623c3b7a62cabce32316ae06e8b76f37eec6fc1f3ac58a4049b7f4ed967cb325a3b55466222d5d42bc020c27e0333942097205faf1ef9ab99b3ef185664e22eee82f410b5a3c1629d33f168b0cc19f2c27bbdd8d9c4232;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf10b26c98914d67923b931d5bdede32392bd119def624e683e085c3beec9f694168a323bd188307344d865c03bb4e38ba05af53948bc61919e0a9a38bb5457e0fc4f63503f39e27ab83dbc35ac2d4e8f9143c32d6e5f58bfe2b1440825e6990614163f34769c8e4cd6a99a0973878b9c443fd0cd02d0b1bbd0b5a0079b3bf1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9299f06320d7a73fee3b28888ccf181690f1ded975099934c9111ed97667846ea9d867b5b691dd4304acab173ae744f0d11e97a07c598e7a002d68663d2ba0d4fe69deb18016d56c4df0753881d5b294b9976cae2e87302ca7e3bbfd75c3ae22e76aa67c61b733b5ca6fcb68998a200472328299281d324aacea315a2cbfe07b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc86988935ff4939858b62c958a60e5ae0d8bbf02326d7bdd57b24848c5a9e61cf9215b4458139e8ab5e31acffde97a2aa85d95762b7da3a29f791b60c7a0c94edf768e9da002720c302fd10e43ba323edaf98db8df61fdd163d3acbb73d49f9403fe70a62c9f418733c2cd5e9c61063548cc0a12cc02572852e7a7c5540b90d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c46eea7337d2c6fae76ba7ea6d485f314a70c24d4178ec6f7061b0848a7ba2e6b4e22f13f8ca03c342fba868fb87126dba8cff53a6207e62d4cf72300fc90af0defe53758396e8e952f99775376232408ee6fe4456c3dcdd979a193828992777b464e69a2144ec1988585b595d53a1075b42bbdd6dcf0557e1ae34b66d092b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha463539a5262c3f5ad95fe08d7b0ab94140a718194855c32e5a29ed6f4d0ea7f259cb381e22bb41048e1a85443af654dde407041f4c3ae08fc4d0d8b9f0e5ae0637471ec44ffb93c0f706bd406658766211f9c5a73f65d92dccdea86c7d8a3bcbc27f20d386cfdac5544308f5e445baaa5829ae06d4f299394f651ec36b46ced;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he02082e64ed040e767b4947b0b6954221794121dccf0063faf42b67db885c9d189ecb674e5fe8ef5d6092edc3fe6068ce13b8d091e78204515e31334a05b5eaaa0f64a1a4a21a295d7017c56f93734339f452bf7f31c13b867bce5d0b08022f5629d060845b1f8b3c02c39774519bee45c4e3fa5af1cc3fe58205750e265d5c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d2b03136bd52689b857fa17bfd66b4ad87f74d0579d6d6fc445504285a9d697af4146a41c7df4c7cd3382da7fbffaa1e9d788c3efa413ae0aedd3064dbaf8a686fd60648f92b4ade78cd04adbceb11869022ce962c496b31e476992ff94fd433556e2b301ffe4cbf3bcff9dc5729739adb431dfc62056d87f77d05261ea501c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b0a752e6e213e1ca944bd31aa7e1d229905206bed274c228b3c07201b34231572d0a2aac0be8a853a03673a47e0b590b4156b254afefbb949cabe140c3a97cbfa2437879801171681b07380d8d433e9f2a4e9ea95a4e58f67ecd6786e17dc4e31aca1b07498a62780256ddba9a4aff22e06ab76595de9c82a73aaf3b39cb4d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82741facaca959561c9bcb8994b3507ce49dda95b89a3500cbe15e10475ef645cb57e8ea4fb3aadf8bf7c6a8640a5957cf4d20c00406505cc3aff0d1eb4df24e14a9caafb776056bd25104f30c18aca47c5e10aeda83d7d056e8532772c80fdeca2cd98bd7b35ac8095aa7721fff310dc8afa0355ad146cfb424d209c28c80cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha75c3a55e3f1a5a785bf2f11c122f487fb3dc3a03ee10635beec472d14d9b250008a3362ed56155caf9093c01aab406e005e96361d02d70ca57b352c3a2958fd9d78f828114d6679846c3ebd8157bfea99e92d8a4b29613f055d2bc1972395ad68f8e63d46a53cbde2ee6e939304a56c7ccf4ba6f30cbfe740c81f309ec2d5bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd58d22d59a119738bbc956d3422affe6f9b9af07d88a7b522eddb087cc544bbcf95bc20aa18d7d7d24cefd9ab6c6b3c3b21a1979f1c44236662fbcf66bdd4c88de602f1bfd0766ec9166736b52e14ef33fb7b68ce0363a01bc258d7469bd521bdced00e10762d25969053f3a7756a494667ee345b2a9caa8bab5a9ef74d15991;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h300ebf3c704b733f15d6c5011533174f1a4133a57d4e59331b89d8caae5a8a102e5159ab5116d0bac7f5ada5f4595d01d565a479ac728fd7629b0f752725921dacce37f8500d60df25df110e95b0f71936d0512a9b6f68edd46c774aed67937c74b84d5cf5b41362063b06439d875afbb35d7ebe87ae7b93dc3e4b06d73520cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9301344ddfd704184148e529e36e7a2c3a25408d9b1863e17b4309716c5eddb98b05faaa749da911c0dc0e1c78078c3ebae62e4fa6e025f512ac2dd8cfc5cbc24ba698f46b3e8fa81f056c22dbd9d7d3a1901627e0d7b61c47c1fb9949f7bdafd9679c9262bdb3dfca059470287bc6a8ed37fd9fefd86e580bfa5828dff43f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd19a4df344274a93ae6196680eaad75ca1b3be9e23a159ab5bb0d5dd828b0284b7c0aaedabd8ba96906846abcc1a4d10e10b156f79c183980b4d534bfdcef170df7e521bc9ad48b496c175f1e6df8362c704c11a2384b58e26cecbd588b9c01edbf2b770a862129bddaa9240f25d3df0927fb0ffc3ce488ff3faa68eb78ebcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c6233a773e3b97ddef74dfea847fbb83406f3fdc70606e9376f3d6d4c9eda77eca0b10824cf04c42f8856c504f175285843de7230b0b4170923a90a5bd4d53a9d833b46c86b37301464076ed3b07defefa3d56b10366aef59d5983d4995b21f9d2f44ed547d1b379a8615b36fbe0a316cc6851a3c573b42333a2ef26984e874;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0a1c03e878b0e8641a55a750bb8ae01b3dd3dfc2668a234e31953ea2cfb75ed8df79ac870aab9b68e0b63d628e4e8fdbf24f0bfe9262b932751ee8c71195b22ef6949c027d6fa4b19ae1504fe104f373e865bd4b50668eda111ef8d931ee7873ef748e13c4c6357cea83aa72791a6e13b3b99362e66d0b95444bf6b623ab5c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he55ff478e33300ebbd099cc6cfec08f4d2bf8b8e4aa32bebc3becd48cd7bea803fe97fb1b3120b50a5365a48d2e0fcdaa0c89c0e355f707139029e87bff1772483f2465af24e11ff6ae05223a55c3a6768f29286552055720bdfef02e1053400239f62ac7baaba2a8b88f9a994436f55d847655eeed967728137736cb34f7235;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a1849fca180570e32d0691b3f0f6a646a32fdcd28bda0e2955a4a49698e6205e1c93c6db75abb67394e09d02cbea6f39e23312502a8a63a3ea94b819691815f7b00beaa4f05baee2ac910d3f7f6c9f600927814735581fba4330c24cd25ec3e7fa98b92f9b68f021f39231624366ca76859b06df9fab33a78be1ec2ed125c82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a8125ef724b36efd46844df741f9d10259ca4f56ed5881a473ff2f0d07b3a93d8d7cf0216e2fbb10c890f89d33709a1ff725f8d9885c26bd0a0df9ae8ed2ade422c27221357c93cd7424e43156922bfc29b8c076d86dd9040a8af18d5724d3c251b89a2d8a2a1b6146bddd58a6a0f27b70bd8f22cb033b8f4fb392bf9492521;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e9bcd4e19744a786a4c9506bdd2a0361986841f12224196e0f1f17d1c85e9e39af3e93dcc8deb78f2897800d9c21d4e02076702c300b4a6c6a4cc4180cde27854b937e934bbcc5ed99d9d46e1896b5e08a4a74113c1ac22c77eda546bdf4350ea87b877e4154b3aca6527858f74e1f5270b8b382fee3cd80f818638f9498e3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc66eff8c36e2a8a3192dc14296dc02802060f688bf5bc11bc14f22ad676b88fef42e2adab16fbe7ab301ff848aa8ed2193ce8810e7068e0b9edee6654f2f7165f5f64b09cc30509d2657de540b48eeae43fc1e34e954335b4610d7f1145e9cd61a1cb0ce485af8dccea88c969c28acd40153259724353f9bbbfd4c3c1f49a60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdce1a8d50443a887458aa7d7e8392ded94e4f7601c7a26fc29a9d3dc42c1ec2f92a97ee2e375450ba25ef9f52d8f34adc8ba4fc6f2bcbd193655db126156b0f25a7f231735eb7edc1f01335b836888d55da93e66c3e3a736e2a4260f3b0ba814b30b4ee526e665d32792a3be47e541820313b499eb239b916cd7115ced47cca1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff9ca2a1921859f3f569c10c4339e898554e551bb63cc45fd8bac02a1bf1d10eb84d092dffdc18c1f664d293bd241729ac9984e05ff8a059cd3f332c681a52ef909b11f0effa2c6cabc86b165cd2b86450ada317ed2380c0ae7160ffdd8bceae430333f56eb246780d23a1ee31eee6a07101027877cb8f7d51e763bbb058a07d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h229b0de4b43bc3bb3c2fe6ac64a19efebd796eecccae98b6353850f1f7b305e569ed452291514f2a92bd364c8ac8ba7cd63f3835195deb5cb4914e007bab2ac462fbfc9e522e5c1e7a2458798d1a77a813325e6d41c3aca7809c1229fe1945a914ad66348ab20db31b86cee24dad5e41d6328b7d7b106247e5802d54e60b2413;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c635a9a132ddcbdda2864eaff203a0621b3f87675c1a0568e0ccb04a0212f56418553ceff91fc27cd8f32d7daadfe0935bff07632525d1598765f31bb72ea4fa60cdbc080b0dfedb04bd1f601264f769bfc8fdaa66755275f40aeea9a210dc4e72efb2a659f14d9924d88ddb9293acbba6b8c30c4f59c6c1ab51eabc8437c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb838e37cbf8698c074a22b11678dfccd34fa33949010111e8e562bbe25099bcd2bba88038fdc7cefabca2dfcb2d64a2c03fcd6c0da8fe1dacedb26914c9ffd23d7edae83c8d1d35132fb1b865f9e06fb51525b42fb505a63a785a1a3422afc6ea30c74c768102e2cc744257b89d6ee0a064f24aafb87f8ee06112e71d05fc66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf07f79d60f68b0a41d663ef88212bcfcd508721d6e66e07712c68754dc21c52d6cbbd711db22a976825ba24f0ef10d463a1d6ed4792473f695c6d763869c46339fbc7b0e9840dd29fbee09cde60b7da1a28783096af7cfbe5bdc327c9058f8796c96a1fd4c70b2b5a69ec1c7a2ce2f797d6ccca9d10c47df239d01f0854cf6bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5717cfa0fc8dfdbc60410933d5d37d4d961d1deba516bac71cbd5263a1cc9f2757e966012112f68756dd011e1925b846d5fe2e34aa15cbf6fe0c76bc784f9422ef023212c5673ef7f587471c3e6b7fcf3dc5b8c5a01fde26687b25e759185d5353624d203a94cd4ab331d89255324b53a426662dada9ff73096037fc623f0e3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfea5bf3bd65dcf3e2cd8f76e8c8fbb04eddf7fcf4bde7da169bca31e2929c4c65d950ed506b50cc34fd819cec16f7d87c109acf8c444a155d5eb263a4427b1951ccfe5ca54c173bc9535fdfc1b2e77fe7a52d644f3576d096a0a00c1302f1d95d634d803c4273f2e594e77352994a5ebb5b74c421a51714937e9fe603c596753;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42bf81904db6a4ae6097f9a1eaf39b2d5416116f783107cca177650eb07c22b3516e68d597508e76efe7c8a12e66e4c53e11ccb1ccf7ed53000a33f9f7b61254d5c82808f6ec9528318695f4bfad2e04417b66bda2c450697bda5b69ea1337a631eaa76d2f4c9b46100596b9531a8e6808c21c52c4ee40ada32f80bd318f816f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h202159b9f9700d58a2cda3c6238fb280a045eb6f1e3fe2d741b0736aaba9add0aca3692000192f101fe32898b7e8b2d43978c815c6a6767b901e4740a198035da63380c683d83c0edff299cc307d2002ecbb5616e01a0ab7b1eb0c169127c632e4c135a21b878f26c45a5eefd2c0708019bb5613754e0ce22bea22f9fc31ef1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h411bb5fa5e0e4a1a2718988a1448ae59cade014ecade6de8df137a5d225d985fd136f9ef5c10cfd539af8ad945fce1534f221b40bb59917979cecb307632610a31c02ac45a031381491525199982ed2853d288660fb54588bbc3e0782285c768931b4a18320e8081d7b5b895196a9cb2a077227790bcb2996525f0102f3d9c52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4555d4dbc3c4c180b462461d6039018d50e87f6a6086648abc50741088cbe270d605d2b634fa55309d6fa29568fc5687880ef134d1ac335530d9283080263fd26bc0e043065c8c9c8caedcaf812091ff4b7c7e5b4de40bc0fe8d4ea725a04e7d3552782e2e1472250d8c44dfdca6803a2d9bf8e06e68b2af4cc454d01744d08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37abc56bcbb98d6073bb54f34ce1606c2f8d50b6f1b5c8545d541d7a628f85d04ebef2a8c72928e2519b2337c7c8a827cd9244bce9641aa9fdaffb36ca690cbf1f0e6295b7dd34c351da4a35b596eba1d1ef132327edce211c4bc775e6623bdf4500f13d2ecfceaf3d3742eae45db9d30669831e75bad611f6da82949a33dd8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2abb690093f0e5f39de5e10be9af8387064abe0cbbe4fe28a26ac9b01fd31ece687932bf32d15a79ef75c525c15d5734d82a9a0aee1c9aa830c437383bd136580c8d94234dad9c0e8b87f7d5f210d78a3cfabecc1352002b01d34e30a113e3368cc640b95936f8e6457d7cd28b2cfcccd6fd0d8546d6c6b5c5ff784225f4ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ddb4b02adaf697ff919c5a16a2fed6dd47c657c57ef778a697676d4fab5bd761d39911afea425aba3ff00164fa2fe96cd4603b6d6f462ea25406d7681977df5a44de1892a687c0402277bf05cbbed7dee2e31d12af06822cb6ac57e4db4c815eebf7522415f1dda94480ba203e701b79922c938ca369cb36ee84ba6bb0f3c77;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ff05acc5acb50203da77dbd6dec149703eda5ea249fc5f80f033881176882b77614bdad42cad6f6792f05dbbd7742dc330bca5b4e07a1d236405d53a5eda5924bbe5c392e970be3f1197e3800c65b5ebe642fd80963993e789544b4cfe8a31ee3e206a8761ce08917cd2af14f88a6e292888f3f8b3830a7b7903309f9c9bf4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8959daf7acb8224560e064287196e744da327ce41ce3c309d26ef4a5f518fb7e8321db96fcb0c17ae8528553a2d454ce58a61b992dcea778ec53887714fe51f0a807e80b50c99de4c8460f221834c28665d0dddb8ecab0bf8790c46c43742d625f37fa3fca0a7180a2f527b2319cb7d34dfb233e75efd4ab94ead12c7546ee05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62a1ab5d1e0b167276d06a8ed99befec6e99d9e8e0c5c9a2b1f6340c508c4a3138c17a96f4d58ae2d268d488c97f64cf4f09cf747b8044ca21eb73ec24ec0dcbccaa4ff849a967aacb0d5b7d596dc2497f43dfcaac0ab3a8a620e35d23df202acfcf909d8860e98cd5bd3c92469b278138810cbb7f7ea0e3222571dbba0797f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b0587e57f0e4462ed8eacc21f88edc1e6648366dc686fcc075364f595d008c46e707814d0c2437a5c3560b800f743f7d89d295d943b0c8dc142885ec188b6e516c76dd3a2970023596d0fdc696cefdde0fc15793abfe289c999aab3ed19af105448a91331a74b63db465908d21b97736768f64bf2cd21a0e64320f3c9157c64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e847eb845e5feb2e25b33a4959dcd3524f78a823867a8094d4b5d47c88ef9ef5dde07280de1fb8d57ae71f8373a530fc5e484b9709016c9188e5b431f6e1a7738511497d0d10ec28cda324a11fd11eddb302fd8ce8f1aaf826141366d04cd876c4ac05dfbc75c5a9a9ca7c21da5cb164bd4240b7f85d107db79674ca1cadd83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ac2de9316e09928eb722675288147614591eff71c51454c64ac817689d2a1e464786dacbaba9f5b3e4a56573934b3250fe62410ce1e5bc5734df9181745cfaed947056b39a28dd20e453e685765a2188ab4543e99e43e205672d9830dc68b3e6d89b517885f30547a1a53c0dcae9ae41128451a78616b4a5b8d5386cc4ec046;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb00f84c312cf530cd59a95d8ea8fddafed1b355fd641e2a245d436acbc653cb7c6acd06bb7d96240d4ef52618e2b997e64744560db7d2c4f4ac32c88d236eb6d8b8256cbc464b7145aafd3a5371d1a537b37baac0e24d58946e6d4493304745f44fca6853c1c98f15bb94dee2ee56941a3ed2d4919c7100b880ae75c4f2e44ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb32cda9afa89ee8501f851e7a8a9f2267c27bc20e70e5244d9a7029a90bbe673dfb80bafacf4d6e7125b72e24e39296d832c75c0402c29e22e5485b02bfedc7b94d181e814d43b8491c6b2eebaac6679404eb05ef83ff55d451a051953e36ea59930f62db5ce01d631c594208b235bf5b7041ee424be739e93bdeb03af3638a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1de15e51376b1f0b6f825783d20a3c1137795042e93eb36cf50e7c6f37f30bfe04d502b3ab828c00d4101cd1c5d2d52b9c345f46e0ca84bb9e6ba6e6eb700eb5b009694c99b8c4c55136e3e68890d5ff9f4521982855faed7b9a2a4510445cb053afd7c120caef7e472bc69dc652f47e94805bc20d906d62838f3ddd70d9e00d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcecf0858f98439bb22de59a03d19274fa2ca6bc400d17ee72e8a286db283974a8706fff5a4d8de6f105d7509ec69501770be06eef001ab39a3048e483ae64c967c5a3cf95bb4003a4a033c552f3f74dd9e13ceb57a82bc5efa64e08eac17771ffbb3d9c1e45bd98dfd3959833d3e26064055bd88966f079fca1b92356b57ef47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2367ba3f293a1832117021db789de2502f002268a806041d7686c0608b0d70a5a3ddace7bc751271a51dae66bd57884364b511b92e27e38caad06861a74fed998dbd03223808ffd58f56e02343d1c9947822a8450877806dca1a8a28ac1cab24b0578dd6ef6980b2170eacb746b0052fce26f21a55491fcf92054a411a061b11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4c3c9f369e32f13fc07178042c3c6d70657acac096d6cff92e452d2166b18d9fe6d8a7ae7e37e83e45bc0ecda4b5f8ccbad4c0b7e3a068ce95de8a86d6128b380d932a513401bd55cba37238769fb5d74fab9f5a61caf0eb55c7dec04da9468446ba98d9e81ff9eafcdd8ddda993d18d8fa7f6d33178a881d9de33e2283fd90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf02587732d31094c2189270e3bd3f5bc5c79930f2049e41111396204956ecf9873efb4f63b28ac7a57b7d6148714f5ad6069cb8794c8838cc86c1460cce115b884152accc443f9f84bd771379f7a793f2c4f8df9f26b9a7df59e61118d9a3a853c45ccb5980a76ee0be92bf28b8c480ff765e6dc950ee64d228e4f70d6e59334;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97925a0a2e74a4f2993b888f9b457c9744548b20b7443f2295eb7d85243a9d29fa49d91390fcabb2cb249829413bb8c56ea29f441ab58e206575afc14a0b1eef4d2f8d79d4c83cd7e56c889eb5275b51b6e23e3b0d1785266cf128f6cf01de6b8df4d889da49ceb695dc8443bfd5c01b3838933ec39057dd775578eb55be99d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h496f7215ceefaf845ed329bf682daed37f2919a1518e2f44d156b0ef4c431d546993b4233d940a0afce67045311da4c9f472b0b8323035f953acf3900da76198d008c71b4f044ed6bfae248809f618c50dc5f2f2e1cb2d432ab3a519344b80c917c9e1e4cdf77ef8a97e079312aa187a13951b1a096386015a2feff49b46971d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbccba28bb40b478d4884377db541a603eeefd8c99c38b0de06b1b89d5df1fe03e0908ea57a55b90cbef96542d707cf2498580a811ad3cbd4783eb63ba705a773f7199b5e56520b41fb932575b15df39e14518482f9a0225af5a2a9cf1f4bbf4740494c5e3045794595b387e499332e9c1ac7bd232960e2cab4f21cd65bbdf83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1700b038653f8b169b7ecd75679be446a561e36eae63c8473889cf54d3d77ae304c0266bea6335decb5dfa3a820d71cc0a45061f1f76414146fce8548c19b540c0fbbd42b2d6fc852b2554fa8f80e25a647fc9e61436513071482cfd54dd457304e97e1f23ed1062fa345ab503f989ece41bc5a07453add899ce9805dcf91b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42de894471c9101fead3a5452b9ac15e44083059f88328baacd6bd9c4123d34f3245e41d43aa5da32e0eeb703e09e4661921802566836434e49089ae89f5a6edaf28675b7d63281bb7e2b0988c974fe78d60cfff0007dbf17d66e75d0e424d981ed1e0388c1de180e2518e449e7b635ad26a72070e464c6ff1a23841749aa614;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9392c5a771d8013e6b26dbb0877dd1ded457915ccea6b349c6f329121e24c313290b511885c9120cae0aa44d3deea0f18f7bc431b78f2c1d8f9f884696f341d1077f03ac98544c002ac221c7b02654314700fdd8a6aaa0f9f5535008af591e04fc83a6e4b98537807036063d5683d2091087fd69d0c9f08dd4caaa4289c5ccaf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86467a805a9c2585d6e4c87346630d24451dd385e8f9bc52a3b1a8082f2e885da72f608fa6144f4f23f126e134023386e60cc8da741878960cca66998ba509d71f3dbbb375ed5ea66ce2f9a2e374dcfea831dd0355a20e4adc686e2e87e2153fdb39d55202807788366e915c24e085d572f1e62acd7a7388133e21769bc19b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c7775bfec0c6451fb8fa9315277293fb6091af9912a041ab98d4743274156608f2186836d2714d2b7f202ef7247b05626d864b96c6b5f87a6d523ff017aaee1f80e6c0764c1b72a3bfcc567b6828b27c54f0e718fadfb87415eac91a46e29f0f9f0dcd0768140a62405d1fde080af872a5cfb248f9a500e30d7f8a9b97692f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45eaaeefdac1409f7e8f93c377c8d5f685c29c20869ecf588eb29439c25a11726b05a4a1a132088170af6acc5e67c6ac3fafd0e49c99e73d3358f3824c23af5c2d57ba5ee3edfb6009843dbdf663c701de0ebd88bb3159c6815375c3c6f43435c068b5f582f404c40242b0819b1ab8f810b8d39873d177f2b352e9c3ff3e1b8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4001b802921767596badfca74833314be98f0ba6573957fcd73675ee0f3d93a0fa5914f23b56813bf5f78ed61a9fab3fc6a9d131877ef3a2b570be0148f247e013d6aa27a670f91a96aeb40c36f2c84fb44cea393162dd5832cdfbfbfa304ffef074e098b2391ec6b1416731efc6a1c554903fcfd913fd097c98026e86ab1512;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f5c836a1661381d961f71fe9f67219d13e43dffd35878863a86876a513d2326ce0001fa4ff4c9e7700ea064c4a6d8f7f41553cfa3913be9db9e9ad7eb65a96cfed39af0c8e51166d3c72670dfce70a0eefcbd3e90e56073da17a87a2b9572b789569ef289a5ed59a99aafb6eda2ebc7c2c9660fc44cb4d7733fc9e625eb02de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50b29a2d860b171ae165bc7e786255e6f4df1f38cb29dd857d5153a5b3f20a4464937a8493eb7a1d9fc34e904541de6bb92d50b45bf3821b605b39db1996f8f5181ab22db2cac1c474513f96b7ad74a8be8e8ed3bb5055780d041e45b60f12faabf9a190191d5f43d3a40d438203f6a67fe9c8b4f50c22af542252e0d9e830db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6bd1840d975a9a2d3e88cdd80c8438faea97a23bd1d381a923c536f11395db775243dd42a15a5f9a2f6cde3c7def04d9926dd14bfeb8ac8399691e149b8101d12e00cd924d21135951e7d5aedf52f8e0f9e11d9db242ff554bbd8910b13f91a07acca24ccf55120d87e8eb07f9202d6b265065c510d06b67320ebfde4655420;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had4c008a1fb1cc9a3ed0f8bffd62ba1cede9280393b91adc0508fa0e3c36a2e55ced527b3c45122f040f037c90edd5210b864b757da5ec26ce13740355f38255454e02f7303bf6af55f865ba583cbdcf12db6534977e0de3f75e7248f173c0abe269501a1efb41c6f593c88769e10fbc0a82f8aa1e9ea6b936ee70d549fa440d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c4a2be816caf22329de336522ebc24bc4c62580b7c53e8d8362aa4ad86392e348f77858e1457b730ab7d30e2a492dd0f773d16db7917a9550612c73efadaa7656dfa554f0e995b49c625aba6cb0cddc27577be8f487d7be97be4357b5238fcd84cde36412ab0673414427038b13fa956a3b251eb20f8bd181e811b4206a1ef9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cae2258bb6e4f4e6248616c6bda1ccdf52cb375a9dd18917c672a99bd1902de8eba9d31602e05ac42e8eeddae79ef72ce905673533e1f85b1d49352e946901f0e33f61b44ea822dda9ee28e091937ac6c5f741c40459c077ce974732736ae9fde53ea1254e8a3166c9ec49142a7b7d14a5ef14d8938ce23dad14eb425d1ece8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd3b7ce440fe83cd48fad63199c871976fd8d797316efb1f05b91ffbe2ef9c5ee66ae4ab219fce7b8b0464eb414b4a5a6b62d5d630ea2d9b30513fba99ec2668a5666bc05dc1d673674ab866feb54156c047f7ad27d1db03706e22de6329ced56b77d74abd248504ae49de5e2dce06bd0552bfe41c3238a3bc0345479f5dcb1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h846414bab6088fa2188b06c49832c2f510e84079db8bf87b1e1389449094aefbec43c9fcd0dfd476ba34fe8c108d94a0034606b48cb8fc943fc1b4aa948219755d14de5835d3f86caa3300c5aeb6fd640111e84cef157b2d76d2ac7c137b270c5f03d37bf17d08e1957245334861c2220b89d71e5aba8508ec289a87a18b3b21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29b977c0ac6aa6b62aaa59528a72c35e7a97a4ad297e6f49025c9dbc823c86d32d262a045ba02cf2db43e445e62782f0c09a024a87a72a931eb7a3d2a9051cf80c36c89724b288240033d22edb81fb5668d82190d8351f210797a5a41fbcfeac4abea43c75041502adb5de5891331547419820b0287f762d6c9e3fba69e80dad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h427a2af657147d93b791917075bdc08b0101cf6b5018a7ac006c9ec8bbee9e63680a0ccee5eee568a46b333d24a4fb68aa5be282711da634ec8717b84656583dfce121befc512084adb60440eb660abe236eeac2d488edf52f0e6a578bf18fbd5e58b39985e2f7fae4bdae8b02bdd830fd9f97cea7b5fcb28e2a503271c170b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d1eeda62c452232ad789442a45b30a6f70349382016b308fdfe348ade38fdd13ba576826c3982c0967b07d4d84838502db5fc41c2aec2e832cedb69e445501b6c0df053d2e583d9b3443f39edfe807064b81f81257dc961bb12c485fe898454b144d3be81a729f22977f6747f50f30a73f076821b2dfa4004a37516b89f8d63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dca01b6d3b09ecc7fabd664f2ba0d8e967d904aa5bb15c73e2f2963bd4e5e28a743feddee00f38c28bb659cdf337039a214c94c90b8656374449842f7a11a9f02c94adab407c18436c88236021f2f0512abb6c0d088830de833abc0da888a2e0e14ee1583c3d8f17fccf65c0b383b2c305c29169ae0c32c7e8b7d163f14fc54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd0e79b55c079d842bf01f6b37db96300521afa8a44c5380961ba73343361f85a211c47fa89ddd3e1c21f6352718d9c0b582f020da68fc0f73003e99e76c2f063ec5d615c001a80f3a48c79ed4056a1b15440531e20adbb366b6e793c1d1ed0503323120721a97bdd8109eaa52d33f46321326c73062c497d159e25c0cbe3aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5565d46d72b0e142bb6b3493c67bee30923e4439c6c1ab082917ae8b1ea677db55f1651a408abc210bafdec920532a880af5c8584be33c5c306c47f5f6292f5ee9ab707b10208bdd343b497509a43c7c59d809fedd14f423c7843900f2922087339ea7d9d967fdf72f0378b15449fbc83b549ad75784f8422124c8486c626ec8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h249edb772bcd121eff56cec2b9b81883ce01ee121aae80c2a8966375f99652e19f0aee7d153ce311b19920cda7515ed4c646626553eccbd28149a750cb8abd8aed7fec93d2f5baa571c553e8dba55e0ab5d47d1774b070a27ae02d30eb8bd5222c72f3449523aabd4d8fba957e05de54df38d43b53d82969b2f88854bd0aed95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd121b117f189c5fb1634a5c71fbab4556279ec6c050343504cbe3fce07a450c0c7ef458b113400da2e2652ba027aecce1796fee43660e1e0c27ffe7dfb60267130adb8b582e1c519959a688e2290b549c550c712c17bfb9a5e8f26c19119d525449dbcfe6e42ac2f13a575fb9c809ad8749a966168893a7f265b28d1c0e0604;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91f156c9b5acfcf78a9646fa1f9e99297bd669fb3cc34159f62be6eae585b81c3238268cf3570a1e7ccfd6a7eae9cb77b38e74c44c4083745e9d6e98092378efff7c4e2066e23ee24f24cf727dd29887345a2b6cdb119f7943ebdacc07b1993f4865d0c2f35ef54accd6c6b219c94a0704ea38fb91b76f275ceb3f0d1c5a1c65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cfffd0038879ce39b97a16c2ee703b116c6efad3d711e8df9eb0b762f78bbf5a6e89abaa388cef111b353291def9e0e707629b68512105df275f7c4e3147d9267904650d5de63d29507540bca73c2866f0cac684773be35a1dffc3f738b5d670c9b29be827bbf78317d21fc4c4e819deda6b20ec39ddd26662ad3570831774d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h423c6907d5a1b53c0a091e9d3c95f53c4cb8c995fd137941ae8a302f905990f25712e78c7de969f13f1b6afd599a000e70f3d1f4ea6fa449fc24e36dffe206fa16d3b28c48d9932928a438021f3ba31f597181762b4d771553ff2c79106f949dddc04533dc88728507ced7c914e042758b7ba65f52586a329a943ac80d88bf8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fe47b7fc167aff123bc933e9bf2fe953c7cd6847ac5b03e24eca4e641d69ee97836c982c0d1313d1a1f3d1294e63a6209fdadddb213c80483c126640021e2f23157183b6f27ab1abe29740e3fcc2eda4fc441912257be0fa41c5b621d97dc98aa2778026cc1a509f2bff54960d0a2d55c34ca7bea004daaf4d2445b2d4ee7c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90e8e47f592d5ec8068871e01f74499055f03946fddbd940a9bf6b3d7b2773e19a4be6fcfc961d7d0fab9523eedf10d7d976c392b6c106cada8a65951ca884fe617948350d5ce635884699f23ed03fcbb805eec4492f7381b8ac7ed3cf03ea6b7ce8fa4494b1b8a6f2692c03b00b40d95faf8163eb618cd63e9d3d89d08712f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4944aed594920cc2f1b331c5e1f68f0584747c7120346ed37230b41d93e614b3630748d09a2f58a7e81146d2324b05df34ecb27a23fb12c2d8f442f37e91862f18a9a76623c74b053d562b1b40df20ba04431ff50887d6a8b2a3c4d9bb111b5cf2fcfca18df61151d16a6ca9baa3ba8ad72c3588c9cbae46495586ec2f719b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49faf7213d6c9f866e844caa5c7d33bba77de0f899b663081e16204c66c16830b3f21047bd775f3ee4a823a96eca56a03c908b176ab3e0ae7c576ebc982804331bc7a5430b159d8ec43588a89552a55329c7f7bc3e9928effa0768bde15cd0d2da3baa943411b2b207a0fabdc43e003fbc967628e77b9deaa1b8cb6e6d9887c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h529e52b5689b65b0baca419ccb4d82ee211fdcdbd1735d884acf0018e9037ba145bd330ce27c1af6fc4f3e1f3cb8b810c44af9b9c436b5e0d919382b2e2124a37797b7d1201d2477e773ac8dc6649f8bffbd44bdd418702131b5272f3000a3cf5f6b279a5c71c36d5245c4a71abed314a25c4e58f2c641f591cc2e2dee1b6a8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba5dfc29e917f7331329f2dd0a58cf140c61076c1fd8a8ab74f522337f21cc595432e8a086bc7705513aec921463c3ca044c23f0694af63e774e0ac5a1da29be0767f675e1f49db0c0705fa7f42a942f669c6f8226494c4d1b462b725a7dfe7d559e0e30fdad92e551c513e2d9e609b67a730f8f1f9cb2a23cd4d1ae998576ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85b2e1bc87f5083e7bcf56893153ef887727694d1cffba9739c6642def9cea85352e885e32c8702266c6792a6a10c11f738cbe646af20578b5e882c4175760921994eab1f2668eb447f44ed6e11b58067c48b6c65064c63777d78e179e19446d514dfe7c906b2c7303c45c8198cf1f0eeea81edf3402128ef0332a627732683;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4381c3d8ea8a9ec46acd6e2eb84188c06f72405a49d4e0810e38cf81aab1638dab07443be90e145b7479697a9e8d6511d3bab8730110ff40cb930c7179501da36fa9e3be4bd8fad1b8e5f93f72c2b059e796a2d48d0832a538b8abbc89ed76accc1cc861eefde2dfa9c68dc1b27220a79b272a0f9d95d63d608f1a8327124726;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he71fe7df8d589f9b1909b607de538462e3bf3c886c81e895691434ebbbb30952cb9e656cdb21abdc215a9620000e93b4d9d10fb5676c1bb064181b997de2e57882c00da1a5cb645c8db73d1c3c4bce7babc19746a715d41fd547ba6630664b0796ed4b60d38b35814708e5fc0fd8e88f9a3973321f550c4193d7ec0c6c70f6e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8860d3c69d45fc301a2161a9660b2d31be280db7d0cd8e9aa9353865982a25b22ef987457ceee7880095fa421dadd78466930c18f112cb8fb3f1f26d097f5bf137e32ea52b379347a4bacb7739db7dacdb6fefee2465ddf34fc16459945820fc40216e4247fb7e9c482764f2a3e0f1c6a06b8db68f97732f0f707921d7c045e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8ddd0794dfe86bafd4bdbc2fb2a82a91c2ec840f6367ad39b34046e06e38c52374717a43e09a0904fb52b16d54127e384c4243ffc6cfaf49d2109396c989636af674c34fbccd52625e33f10e89a9c7f9b85e1e15ca39990bcc7f0c38f0f5659af512a12ee3b7ed08d0b2bfeed40c5ef639d07351884711c7955ba892d494ba2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffd6234299ed6b74829d49095fe2eee1af5c56183a30ec4387397ba49d1f33227e16304083896b85fb7267d50adaf260bd38ebd3df23714eea8d544fadc3dc4da8ed95a41b1c2cb69bcdce0b1fe104ec28f8e5c7cde98233242582aae1a830a5d0055565c0f16fc4fd4dc5fce5c21db3497dd4e98081f1bc88c85f881fbae9ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f475fc0b7652a24511481e41ff8895442f52d011ec7c593e9914b9b7ce6327c1d8336a9ecde10397cf0267931ed9084d4ef06a6ab893cb342c51d4eb12a66915fb644bade19341ff6ff425ed708d593ce537aa396665e468ae442ef37bc6cf37e01518bec025bf9878f1610bcd4cbcce8d265191ae5071e2d448f86ba38e090;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee84b85f5fb7380371a244bba2cd837dcc9a4a24686e39f37146ab000ac861c96a033ef738fe8b8812e82ecc8d26388d74e71f124babc35bafca938527650dd3660e33a0dd22ca4f41b6b6a8f03b00b0a2191c58148e9dc45d4ff24b5e6bbc9b803f230521659f3e0b36b44e9c44abe6edb335855619b57bb50069725f9fe57a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb034fae57b980b2f211ee2fc4f566e27ed3e7da6f7b8bb76417dcb6ff1511c55d0de1263069ab0ec12b6e802cf96c74142b65f58e13bf1bdf14beae24812db062e00bd38051c36b7f650f60700418ef74f2ed973dfc93c75f5f85cd3419e5948e7f9876028d13678e54d7ddbefa42826603fd2a5995d5a22b59649822b863a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f7199e25d617a4da3a8db762f55f6b539c5f75063d2055602d67a29982d213a9564b208bbfbe71b609f79208fab76c0a45821fee57a16bdd61cd5b447fa6144a46797876850f733a12523e5910741448b50f860d53461fd016d76e8f2c2fb2a7cfd77999a689e8f97515c3865ba19f6fe3d218dcb6cc5debbfc2ea926dba391;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h260fe4c3990b9b30633b7cfabac5876bf67da273d0da6f2ea6e38a0d4aa765c88659cf2ab7d881cbd943d5560a860bb47de8076416d5a1104bc29dff6a4cb4125765b1f9d2c84a6799719cb1c395f1d9f30394a341840db3c3cd56d63ee8d85452e4d687f859d1b28566c107256b91941ccab5607f0ecebc2ceee857207129d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9238c4a777d0feb73780233c75690a3d1381037bb94e77ef30c0af23fd580df40000abcc74cd47c7784cd6a5c829526be2a683a27388592bbfecb0cd8e04694de8cbed7f2fbd3b1280a68963f8fe10a584568534057d927379d6e83e7c7188e8770c65d3fd328876ab1c79ea2ea2bac1be67f117afb1cf64f169e34dfc8569f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca9fc4e33b2c98b9249749967d98b542fb214cc1e6ccecae3adcb8486dbd57e94a49af2404b143fecfee5294af983424eb65b126adc840544be485f0c03fe275fb455e9898b3343fc7551f191ca71b991f1721dfea8438ac2a29823f15ff81d1a2a26f511b906e8efa6eca4f618509a14d8d506bd03c28741b154d31291b26e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1667804e49df2990ad30dfb68d2397747e86d905f45c53493dac136fed4d8cd3eb6963bd19bff764ecb1329967e3dafa8f7bac1da0c3bf458a8939d60334cbd0edf0885d16944521fa37cf417550d7bb169211661880253d5b3a877b99ffa4547e2837fb9072585df35ab2f8f68241d46ec44d3c62027a2f998dbeaa4f881bfb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58ec89d761aab4f02593b9ba70a6c7eb92727e8f6ddde90a5a753aa2bff849b4254549bd7a451b8730e5d4b965a4568b22d1d0d2eacec70a02982e5619514ad9717b46c2dbf2b7071656fc3c4b1bd907dd6275b6c6f4382990a848d404e2b19933c39a84a23db247a465e7f36cb240ac0c0d52450b8b41169633d12da251e985;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h157c4bf5dd25d563a586e6ebc579a7a842e33307ec235526f048459936996867377021d00d5fb98ae76ab7a63288993d0d7d0660cba1ca68ae4a497bb20e647ec3b3ca8293ae8ab6f804bc06a077dd9220d83e66ee6db789180296d116a04dfb046b9e4c65a3bde4edefc0e297a1791cabc955f92bf91a9e9a693f05f8feb203;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55a19ab4a05d7f134daea332af4c67b2afef95b888ddcc12cd7093c35d6f49f0daf06d97eee0fdaff4537b7d76a4b7186290b03f60068003fd82a1765f6fdfeb7250083478513c79f68d43543ec4451f62b14497a8847c54b0ffc8d350c25138df450191abeb1bf50ff82084959880ea74463a4b903a31882ed420f9c38441b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce10c05341c44277cd0ea6943cdeb1cd62a2550bb4273c08cc8e5a54c5625bb02ca908e63b875d3607e9622851e5bad398bff34df72922bfbc643eccbdc2527f2c9891485808a82222c0468866027da3309895d3f7daedb5b7accc9bad4c412d46a1b0eb2bca2a9c715bd834c447350ff2ebe981d293acfd2b110d7f31c7e6c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9c7b3f650708974797b549bfa95ff87b721805ae1530b60ddc3663b9036d4a929e0b5dc01d8027f0daa814c36ef29b8e6756e4aa4cb6fe75c9a50432a1f73096b316f154397f39ac668231f6fba3462f95315bd3eb70229555fbdabd3ff1180c454d627a7839761577c61e553a87482177e161f64ddae541fe0767f59583648;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha30649281784c40077af2538ffde25c4770aa92689102004f39217a27bb080d05ddd4e0d6049f39320e553c5966ad3de3d5255d003641e591d3fac2b8e8ce60c916315e0df137c678f309ec747d24a3b42aa229df4ec727927cbd955a2572ba588e0e89d826bc13259ee0c1a5d64be813b6fc3db7cd75a67350fd3791ff57952;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadcffec3a28dfe100c43672fcaf733e5f5bec7e601b15426261d2fd824ce3b57b4aacbe0a0a569d35af04d2fd6cb0f1c1b0f3d34832dae65f4c29e3b5417612b1ab970cc5e5dd3c75b64967de48b7c14513ead82d27778540a753a6fa1f3d85a6e40a269997be9ddfcc529bb8aa5ec17fcd20e0e1ae5bd47ed4560d24080d03e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9ed2f66fafbdb12f50b85d8d4bb68e3beee364e513611f25eb92ee075a62ac87aad1f0525641796ef32c14db5d7c05e1a45634f8d2c303cc0df1a923f5bde1dc4427c4d4c967043aba610f8052189fad53a2f442e1acd263ace33a43ee7c9c2b1d7220d38162b490b28ffe9276a8873ba44f06e0ecfda215be99df2352a24fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a1a19d26c82ab6e982c5af963484fb2b30873749a6ba29a0bf7de6acd89e7e9c30594a2e6842752c224dd2b47351604133db65c61ad6981a78fd2f25b2274e032fe600ec82e1986f654c59134bc70638be37ae4afdde92a43e9547eee5f27f34c1807ca7882b629920d96650f3eefb3b39d7e1f51dbf63b31718727d3e5f846;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f61012934b7993f9db544871947cd5a73ae8b39e4812ba02708fe4943cbc6b473eb79683ec87957c65fcd83fb70b77854c2f3c0ea05367763105f843f554133b770810a69f12228261eaf7f26aa7d4a507953acaea93bf13e69d3910070399d3a1858e3cfb5dea3d36d09b37df4068ed64aa41328571ebf918b7c7f5ce42ff4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a298d750fc043042eb8d7c5d083a06641449ae7eae39d73a35a7c1ac583e183b12decc17f2c8a247302cd6ed16ed2fbb4938bac8b957d0bfb46e2e44e29a9bac9b31cfd0575d1ad76e44750cddebc0856e4b069dad0bb243acb936c1cec005a14de9c2978ca60b89e5303829e7085789a4aa0ecabd19f4b71ae0cbbac3182cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2db0a036768a8dd58331207b753479c00809b110e724c0c45737f634d68dceb5bd9fa274fc51ac5345dc035f5df5aa7b1d69e1872009e49cba467e57dc8f1748f9535fef410edbb05d237e3fef5da008138da327d25f6d8852092f6eff95621ade6e57ad95b64910d626e63c6a214c8bd89a485e5e904be7407ccfc85fea60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6226205ddc7cfcd403888659898b0f4b47e496c552c13fb3750d42eab235216eae7c1ebd20498dec41b84a3b789f25f1708f29ed29ff816d684d58cec492fa7bdfa5d3398c03751dd4ee9b7ca50c13192766259335623331101ea1a344fd716cb99dce2a3f4d63f13c810ebb2e3ff2b40ad11c50a8d6bce68c000f10fd9f1be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc41f669b541538fc721ef3c942ed03961686fefd7a076c7981527d7993582b057c8bb61d49f42bd6331032d05c5d19e54446514cba83f3abc8897a04841e6ea025841249776725655261570c2cbf4057988d2f31fe5223306b1f2d03d404e854cb563fb9877643dfd73ca281f033cfe735b136bf24d46641104cf1e366a5129c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8629b972f28e3cfb1126ede6dfca54622e4595c6d6e55819d0a038307d4811d30f2b2e815aa35be5589c559e00a75fae41b8e6605ebacef4a2a7b36c832107759f2f87a2170002bbce8cd3cf68c513a5235ccc8f8110097ecd8f5de78f27444594ccc791652399f5850adcb5ac801bca6da278c877a631893fbb0e9299129fe9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7388a3f292bdee6a384eab7309c7d7457707e531dc7ecb5f689497171bd9b7764e319cf5bb8d256f39fe9dcdefc63f66a521d8fcd9060ec2e0d1e9dcde8017c11f6e50dd5b4ddef106ee37b4f29978ba94407184e81e4eaa42ef13adae7e9a03c48080a7ef39de90787a8f363419c39b61ea1b084885f7c3bed027d7f24c4b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52c0559e99d77bf001bc985b51e0af9b4f5316ba1833dd669acfe00050c5a832cb609a7a95c44c9a747b4aca234ce50211869686843b7a0e06398ab3cf796c3516bd47cf5c8c2971b9a1815a92f32622891679bb8741cdae7525a7ea186ab66a0156a4aa6f14a74c27fa2683e421c39b58ebd928282452964e389896e6a962f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1992f71024db48201a5b335982b3eab706af63b7552b46227d4065921b1072b9a20de576a5a141f7e71e340baa54c514fdb267ec1a42cffef40f040c61c7a473e0a77a0d9545b87f2fb78c45e15e9fbb38d3cf07a8ddcd511edbb183d7de26555bafd4fd1bc05d92395cf0973fe4d4650906898505cbe1545aac2b4609d3d44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dff00e48c8fe0d66a5b27c37db393f1fb776de1ad7d1541e99f1768441474312dfac7c0c7ec388d2b9c917c9379321d55d083069037798447db6543b2acc72811f6123ccf84b8dcabc6da7ee1b2f7cadeef245a1b253bfdbcfa7caf86b8c1c9c3cf9c835b1e4bcf93ca3d0a15d8c0ea134ae27bf073d34d7963466fe5540a16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b1e5ccbdb21041042d542776256a316e07076375b0a95afc55de275e5e83e5ca6ca3bee7518ade57efcc34c80c010c13b9f6ed840e163180487461c827a26d42d57aec44cea23fb4da494f9152ae449deb663e915ff49ce8e2da64df5f6d770f9c8165452f7d22a75629e03937c19b9cbaddbd3e045deef74d0306cec90f18d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h480a1f61fcfd5ac3f606740de50de11b240915dc2e685935c80405bb19e83cb12af221c53ecb2b175e239be58ca1c886b91a68c992877b7812d40c33ffc6ba0828fc4f0e5fe06f17107ab91a35edce5c1d0d486da0d622da027911f7997c85e8f012fb556144bf289040c675fe767ffc84ea83e926187cd3c936dbe4bafc2b11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa578c897be7e339a1649c9f702b3f38143e7aea189e7a451c2ecf21cd609049ae27582f0ac6bbafb5cc23e1d4495a0b67f7c046629d1f881eafe69807b022a96662b2193b3a70bbbb6857a1a547c6420f25018d1ba8817eceb5b1b7b981406d4fb0ffd35e1f767bfa1b08e8f0b3608588475cb65fdb67a4ab8598d3681f4d21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fa019f683236ec94ea54dcfaa91ccbfa4e374db1f607332005cffaec0ea6c2080c82e6adfab53d4d24efbb591665594fd20f74834cdea65f88969fe436c68d86a066aeb583c2207ae11481f7839b3af71ff34da149de60f6dc1d943f7bc1ecc200f03f1a598a62377fc956474b1f4a71c6a054aa42c8522a8f3dbdf166709bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21cc66465991e6cb1f43f3c2ab6488d454d6e1c3d14b17c008daaa0e19daecbd05d92466bc2c02f18fa03ea616cc5c85a42979c94261741a7a041beb0746b0284fd1e8de8aae9a798b7151c8bddecade714820b906529f7385eeb02212905458db092e6d043edb39f1e115b2f3f0630c5f35e08faea14840856e3276cf4fd2bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdf232ec811b0ebd74f0d300e071c3da6b4661c0523555f71d498d3762e22dcd758f5351156fe3b6833a1fa39277f816908ac912137fe4faedd3e9a26b023b3169e44132f3ab00089f68a4ba0e23c08571018ca139cf58d88ecdf6063655ecd5f56d3be646a290ef98e31ce35023e6bfb8f90839789dc41625d79aae8f5278b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6be648075938f820702709df1522d786d0c9dcd5c62afb9f86af40652bcc3712dc15f1cfd88be86938ae6626166077ddfb86faf01916b841fc85628959c8890bfe6e7e7990c3952ef03b452cdddb39bb89d18d8355130b0049909348c9e7064ac6ae81e24573f8e5b5bd2adfd1f224754b21fc1b1f1f0e820597ad8de4e2fc42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha599045c0e50786312e4eeae9d1243508f4d9dd58ac85c45f601d9133389f293e88ee9a3300454941375d9ce5e2d43d1334a93bc00457e8d36e98cf4f20cba729228f87701da8e45ab4f6335b206034e506df4d78e5ebdd2e2500d01fc243d6f5e6c794741e39db193ab49ed0cb565a39071747135adfa027136aefa837fee86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd76b56b4bfea9f7f65e4f421c4c5af3a168519cdde8cae6c260fb1a250af90e075f52d2c9c12db1f15bfc28f3433ba786b1f1ffe7e4287636a3775efd405236112609b9deeef2682e56d4b82d85208127ea8ea07fbae889336e9487c72eba43a80475430728afe09f618438494c6a57db84ff3d6981f10ced38e08d451578924;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb02a861350ba605748c088d7c21f5df81d3ec137d217a3db66702d67ad2d7ceb2e6be5731a87ddc7ae120083b5df3d243dac7ef73d5d7a9a13e637d505f64e5b78b3c8910c96e0a0068e2945ee8c854e954c7fbc68efde8b7de1a004a97d928979e3184bdc09699e5a291c303fe77de86bc76d4fe2c8796d2ff23af9332b11ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cba4907c44be19867c97fcd8b5a8f98fd79d381832076168efa7463fb90d82323aba9672c96a7e0a600d7bd9ac08c9f47f096a935a3bb14e41a74d26ea41653ad1f8ee1a180ec9ca18ae1234f68f4c7aa54321fafe9ca71f4394cef04c1073505cbaab12586f5d2cc1d8098bb924eab50ca0f1c8693932159a619dfafd69e71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cf8c2cc5e940a465133e834543a02eaec4e68580603b589c8449dc00e3d4afec73e3426741a962f92e8623d3f17fc1173f673c8dd5f219976df3fd2f23ef482a83e97e65a2f46f28167519d9bf46bf921529a713a51a5101ad950d24d91b4f8d52feed9d5deb7851874c37ce548f266a65e85ea8175826819aa231f780660ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59bfdabe43986a287227279ce37af0c6edc933db319c277f9c16c705336cbdd41bb45b51f62cd06fd031279efb77e9a032ff80cf7ce3db7dd2df3e1ba50d54e0fbdf5f167201e295d3128112e280ef7a9dcde5b3fdd7dfe3c5c6702192e238582b4e0bff0c1b9f6edf12d6091ccbb9c0247c278554f2faf96f6a82ddae692299;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5cf6c2c160c9028cabb518e1ec78defa7baba01545842dc225f0d527be9b130d2fa2e50d9f8625537c269b1d933fa06ffc18d515896057fabd4fadb5e5d0157d2cd02afb427e81709e4440a79cfda0188cca720419ece9f1dfe3b3374e1b1fcde00b2189d977f7ac6bd8d972cd0a129ef3269765871dc4d36a5febb130f05c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ac9aa8956ccc2b3af265b049c3d9041f53a561c8b33d85bdab6d28022e354b08c5ce29e7c51597d2ec5f848ff44aa2fc754d45799a2c04e48771879635eda865aaba25d948f343b6a41251e517a71d33fbec76d52b52239ecb9bf5d882bf838deb7200370a6bac7422024b4ad45fdf90269e01ed2f9d10ed030e0049c3c7f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a29cf9618e1cb6d3c0e532b1bb6509695aa339e0d6b2e98b6a788652979d79faf5e5fec4d74d2c77dd3cffd0815efb40ef3ddf62222cb7b7ce5e3a5e33bd007aca64a130c4a99057ef2e47cd24134d998fca07af3e252084ded7835c32131805c04cf10dbc0ee1ae9ff3b63f78a74560c4d3f1feb0683503bcd8e7aa26c87fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb4ece358e5d424c7b45cd76df1f823cc3495ab24fc94b584ca2a57cf2d7bfb47515949c311540815736a4ac82e5f8dabc4158f6f8cf4a3269403fe0044435fdde7610f8007257bf2ceec8461429131b94ecaa35fb9144c2840c5964c3f8294b8211014e73b10837d2e00339f354a1584c7eae3c924e87be6f7bc4565f45af82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1f1213c9c4be5df958552c7affb72c5dfb1947ba53ba005c778df5099dfda09809e5c115ca03a3a88ff96f40ec4f50923951874856ff17e01af3454febee85d9f3b43a1da084be77a051249b037bb105a3613b570c467b0a57f1e9d336801ecc9c4139f3420c14abd5119d06dd98a66896da4063f79ff14463cd98fba702478;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59880f9592a5dde222edb501d057f9778feac7c4c991b9371d019b81ae9f48209df22da3ca0730023b9b323a7a81c8dd597db1cf9aa5a5a46710d3aa7221ae1c7ba0c2eef2fc88ad32dbcda599959f69e7fc8d64270761bf8bb2210d05f2b9c0cff3accf82c0277414420a1d0ee849ff89b3afaa180e31978d85a991582995d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3463bca8c64ba1ef708dc0b60d0a67246dcad2336778dc6175138bf3ab9f1e20fd70531f567dfa7645f79784f2ff450ef3a4c6faa4b0cfc7738432480dbb870317039300dcaa22f8ad7db125f8675a12994b9a0188895ccad6876edfcaed018b3f454aa6f019f290b60becaf71abbd9c1866b33bed286cb27cc30421d1a9238;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h835389183640047be0d0f4ad16e96f1e44a4d513c9de8dc1b3d2505cb165c1bb6df6d06c0f3f81c97963a0a7d2220951a2dd96eecc4d7295fb04b4a0fea641ab004e3daa8bd0bf13bba696d2616ceecbb2a346908547b05d0f5e165b06d64d15f0699c3baec9a2dc88e5744c82f62dfde7a7afc516863552954c765d1e445e3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2fe242f52e3660b0594097eaf3634fc48b124af0eccc21461830d89ada6b92cc0eb2c575208bef1de4253aef93e6d7537cfe0bd7f5f5d62cfb78b48c7dede0c5a835b331d9604d5cdeae681e472bdccb56ff8c3a0d867c1ece85dac8cb6fd17c29584662783cfdf8984d3bde5f12142fa0ddf2271d5711126ae15ddc8efde6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ca29f104b478a1ff0b1397630f2baf0c273cdfdb40e83068a6fd833dc72f733765220334741ec5b3074c0fa6de7753031bfd712908cb13e059e40ec2eaab6e397bcea1adc17351f7c535a2d842fbdd06040fc15601d8712bd883d11d4af3863ee511c80e206f43fd72dac5963a2d0f87d4f837df1c69282392293191bd2ab4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f0f1711336ae2dd8e8c4f0168f3069f19982a1ca9cbbf92628c01a011dbda3c30123c84f9203ad680e26d531b76c0d6a52a6c502e72e690c6ac69c41c3176696cebb6a31c9bf22a25732ea986b89ab0c3b8387be9ed416c6d1418c0b9158621387a6cbb3dae494ede80cbf6c2f23cb6e84dde9bd939b1dac178adea0236b022;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1a131fc5b288f9ac9728234b96a7ac2b0ec8bd10b06093fb9151b4c86659b92a8b8fe231a92e27777cb67b114549adb34ef2794a483a9f3e20a841d58de0802afa291e80cca1f9910003abf98b8e34c0db27592633622257618ba44ace8f65a47b15d9de80ef87394223fa2c7224f4352ea471ef5cd3dd218025720f036944a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h668965d83f3a36f767d95ac51ec1e8a0f8d35b4da9c1ca068a5e19b38ffc708b18093cd1aa0ac25a971b75690d8e7203a318cd57113c6795d3f4d2215239d4235585cf26f38a84c21b133b148f81814c0a252c922c58ff93ef9632dcee9414e338a851e94c3615cf5bb087cd5de3a9e493eafa722048496d33a9146323718b35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf07a6623a8699b353cfa9910c47b8f77107cb75e1341446a437c9d77bf4db2bef1a934e586b774070410e9ebe3e5c8d77f95361129471789351aa398b801e296ce5ddd958fe0ca5764aa185244b79e52f7b04d65317b12a5ab0e7c66316db4f42c70bdf7b78c0fe81b41177ba6190b5182a48fe1f95d7a78e18d0b03748defa8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd814ac7ecfc1e25ddad34560f9efbc5f58743260c57d09ea6bb4123803554b4a24cee82d154106f77073c0315b5ddfd92420789c23ca8f8abfb5a3878eccc422c6869ba188657b3b49d80add0330956f85986b12639440e05d206424a96c9a18d386ddc32bd3e8be38c6ed5a5f944a3731efffba26e592924df27e40ee97238;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3af082daa7fc7e0794c6c02dd06c7c797bcf5a9452edbc8f7f16daf76229ca2f54521fce401f4a651be17ddbcebe286453ab85024e33603d877fae2527d397821aaeee77916c3ec83a96cce25acd2bf0b700fd32829c8a542cda2977ea2785ea74a76dd0f93a657ca65d8ba6ac3bb7f449566b0888b27ef12de59f1a1d8b766f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d6df1a7697dfbae89a6c1a0740dcbf3c7b205536342498b9216b74db27598b954753f3e8d31de65b5e91a4f2c8112fd3daef99a31bfd21cafde16bf3f7362012064230265f293fad23dee205017681185359e00550de4d41f79cc6a14de880b4fc2526c0aecc153941b1da07978bfe01373985968cc8fa8ffc2d8a20d78e327;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a05156503a351ff26bbf9bb8064031809bdfa67810a951ea5660d7e5c1046250e4ccc3ce67f6880e543091d334aafa5181f2c7bdee95ee39c61dcd9517c660862b24af5c6c027e540985f04c9abdbc441b970e32b073921629aa13f96f7cfdecd00969f14938d5790e774b05c659c4856303c5fa5675d791b9d2449eb0b4575;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbac95bb970bf8fb20e36e3135d5883001c98e91fe2bf718aa4669f93a370d81643920da6528ea0f486119f10ecbdddadbbfb9413acc1b26576fe7ca72cae4c08a2b872ca933466eb00e4b912e18f295659736ea1bcb0e36dd912822f3aeca0e4547b6d3538f1f5f9c8cd078d71d4bf83cf5a599f9b04defe479f5ac566fe88ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd98537e7a36044b0471418b068a90a3211a67f0e6ee62c919152e185616133e2c1f7ef9bde4d63fd72770b1b85d45efb102b6cefae651802c382a11546f56f6b6fbf2d2018be0ccd86b0ae0db3e299b36e86c43d94848723db2817f9626053b39b3b78f0ed87eba942c3243a011509f242adaaf3018940c6f80d449548840f44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fc77098776975020ae93e6cf28e5d1ee26dbc2a13447d68b1af0a535b845f8637b1a65d11b6c7734544356b71c00486188e9e9ffb8dd1f9e7227636feaccef1796fa4d90a0d915d785685d1e29b641539ecb3d12a0f995b5f3d96312eededf139b03da3393e9765ce9d6a8e2dbde2e1baba88b26057dbb94d2feb8b80951e35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h791a95fab8ab939bbf24ef0f4dce6e791e5c7869d79bfa033c6af05cde31c3a071a1b576d56a8616b74f14bbdbae94b09171699f3369a39158d3967c13350f5ff074401e66abbdb38e1ca3db60a541937d24915e2a6383cdff87c22fe50875a09acf5e9d8c520e7f25ea8cbaa749478ae0e6276494a40936926ac2a7c9b56fa6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ce3d572506ab4c664e047a686ee8fcd90252aa2d87e26080112fe0b68cb08f56c852aec98cadde73572d797a76726b67fb4efa687f4672c123d312721e6ad3e9cb2fbcc93438a034aeb665528285992b84be6fa24c0f0904867b0c1762bc1f9d71f9979dc9ef6645ab1e2455ad2a090ae60bee84d3037928865a945c06f9568;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae033638b64010208ab53b2701ceaabc69f064e38583ed458902ea105f75d8f6559459c09d43184156d8b7f307323d93517022f0e9a0b9346bd5092b31673aa7924a7a2489d204675d9b76cab8bad29195550e39ad45ad3a40d509f3d0298340fa81c6fbcd7481de4709be7372c9dda45e26372411b541a8afb9feb255057a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7f08a833a977ae933382854461dd64844006772d46b29ae96b4e18148ffb1af4c4ba68940ec1fe12af69bfeb51da70e600a9b048fce37f1ba039891348b121c29bb54037800bdbf7875c9862af89d7edb16dce99046afaa3a876be811a49c3d64c275612426054089756bb24bf6cabcd482c17668f32c5c75bcdc7c1de421c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b84e551ae13fc8f28bfb3730ccecfa4b689956a746957fce6c2288622ecbad98bbaadc6d7e04769d1d1d295a5b59757e25b66f6f35ce4b3c5efb01ba3cedfbcef652f979d7d03a1312895e1ee128840a6397b26adce3518e6fed59663dc0ed0aa0b2fd8499c0a87a15a03ecc220e2e73d1d74183d04772be55eabb4a040ba6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc77475b80eb45ae76a998204882000699e28406dc24ee8679eab5723c965ca5df639a898b88d7864f9cce4245863ab96799e299489ac6243b889226b6d4119d137b75987c07dfbe2978274fe1eb0aeb543b580d73a6b220e18fff1b2d37ed81890ca7ed3a5c0ef20d0ba0aeb9101d991457a026523f6929d8ca7a476edc7692;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84d5f32febecc83d5973d3a9af0d3be3803e89e9880e1cf68d78da0faa6cf649b25cdd8ad9ff85d61b1b99cf1017463561a3f63edb134e5c07ab0daad57a5f4da7c411fe5a08c832ddc73eda63674637ba684bc93193317d2b003cd996e56367ce4368145e555800f3345a51cc6786305d356caade0d8afa81798305c58abc94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29ae9573ad79646b64c00bbc6681f218845da788a3ce05f4c68534a6cdf120b31165e1630b277f365be8ed9c2f9fd7636042dac9a18049c829fb44da21a319b15099ff4eb8c8899a4b298fc647b207f853c2db99977f1c462611e195d351bf9aa3323c093a63cdc9704ef713063fa47e86a5661fa7d8fe739969f07dcc0c955c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf22b9f820228f3c6d95f66d87398f51885b8015ca31db9605e80476c6d4a9710d88fa405df003216509c98fbe6634fcabff0cc65fa5582fd183138f420f3dd3f8e70170195abef7d2f409bc2fdca9c7e7aba9d762ccf09faeefe7b64e26118b6a35f6b0b4dcd59e32617c5c5fa94680d764f1eb953f8988051055f720af178d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9acd0619427b3022ea9ee9decb1170230a8aa9b0bad34fb52f5560a315d962c2b845ecfd92aa8f704a2ff46d6ba0253377c2bbf010cf1f320122116dac817caa937b9e7ca44140fcf2b767b36c21557333a76d2628659040c5ec76aeadbb171f410ed5e494554d0d1f4646d0bebc3cfd04ef622838b7c051dedf6672084dbbb0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha533552a0f34fb0fd3bec64e2de20c6cef443164ba954ac26ce495c75734ad8b8f07525146f27fd954460fb8c641f0351c66361e97b05d87fc7480c57bec720462be223d05e60e50a4ca8916c87e14fbd4b17c4bc4cca3d36f799f4a21773079dfcdbc91e4ffc4a78000b6cd5de7f9b2a320cb7e7a73f50a4e124f1b7d016dd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e4d49f2be0deb9e736cad04defdeaae0ac80615ea04097dca5be7f19fff649f8be150b01d2e983cdbbe40830984be711b1653ba2ecc7855db6c67ff07d22d6bec8cf9eec06f9fc6dbe02c5dfc38eb764d5150cdbe9a08f0513d7723ab95700affea4bec6db67d35caa2473f495331ed8cbb5253ecec0934c173350d65da89d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe447a2cae88f87e2f295354660ccf6ef54a9543299ffb476e1a3f6bb2c6078882973e77a77bb0e18a9a05e49e1574cab8b6ef3189e0c83b6ec6e12fcc2b8fd745c15be3d4013dbd5f658c8496135ba306b9713a5f498d5ef9c1119a5da5e233d71bace4cde26bc2f5f222bc3363636eb9e71a382386fa4207c611b585fe50f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf09a238b399a64b2c5449e5d3192927de6cc5f169ab2aa5219dfdd5b4e7b4e9f3a042755843bc58155561d936a10d644fcea50bc25c6d2db7289c50a941b340e02a762340fe3e852e9a428241e3eef905aa23cebec65d79c56e9c30a2eff9c79302909facac5ef2bb336a5a43e8ac3a295ff48e2b4a3a9fac38a867217d09499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h688f474e90f4ff93254da011f52819a026f2556523200a4290e88ff9154045d9f2e2d47da9335151bec907cd140b4bd1c5cd5d1b845120be22f5646e20220bb3f2f40f2f75e599b2b73e5adae5a0ce5286891b6442c471a8ca7f26636196a7f6ee858b0965e63e99963e91edefe423138596815cfa5d3312b98f0de225e7d6e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c02f78678743d1ba37b1d09a6967ac5b67c233d000faea58da7eb789b1150b335645ff2d40c0bb6756ba976801b90be538b728054055ed9a8581c3b975b1d8cc79fadc6f7c4d4f2b66ea6f282d5bdc449efbb47feff363b768ffd63d55579abfce2c99729ba3e36a9c6fda5b572ee832a05e1672c5d85ef6a6cde5f695d9948;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2b49da353ea31a8e5fcc6460bea967beebc2301ab9137dae5e3e4b22c27bef79d40b1c74f8d18f66d552fc33305c482ea00a681955e9c897478c75ce25001d33651a20e5f7fc903f8517a787178bec75f17cbb3b8c43290d2f99e656cdc7eb1099f0b48542d7bd21d00866c290c877e61294e38d434d69a0af694a4645d597c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8104c2640b2e0460ed9c4e78f7906b9e44e23c1fd4b4f9cc13b2b2135acc77bc379e085c6869f74c92e2f11ee2ddc835345a2b74d7f0441360f77fbd2eb9718123be79c5cdb831ed4097de510eb6c603a0a680da6cdf5f79dd48764f8f0a2a5968ded0b74f4c5567661a19bf55902cdb34de922f36e3c668e03cb8d039015ba7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc23c780860e6c57ed31a57d6f9c102b791dab8eb216baf41c8aea9bd0e0b4551e196675d5445099eed8da380cd83a28bcf9d504685bf53288cd72e683ae1b68b8510d28b39ea99ba1e8ab04882eea2ba156444b8560b6ae3231c9404cb00c94c1e0ad4cb92e63bf585194337e60cebd6fa3bafb43a64fc955fc4a893f8740249;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72576736c79736f73cf9d10639c8e33a115a2bc1112c9304030ad890afcb9cdb517f409c13bc58df555a1123c226e8ea2652e8d0775ebdf15540383bbba51ce1f02729221bc303af434682a78aab0aae9d5d2d0cfe1301d2436deb95002edd43579af2532bba1a8739defdc12da621e8790933db92804cc58937cc0990cddb7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21635a1c5119330a92f06576344da041078a70535b5b69298b2957a450d006d208c2271fcace06e9ce703389a8edefda7d9d3313825d630a0d67b92a50c4368869c424f22693f838919e61a48e617a745a192f48cfbf9c333e4714a0b016d9ecb4726a12b2ce95696d52492c5031ce71620d80d93d2292e0ddb32fad092300ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h981d21803f7e4080486c5663fd33906af36b71cc4637dcc271247248ae7fa2af902a6a2eaef3a318cbbd6cbe5e3e93bd83881c7fb5cef90d3cc8a40b866206b7e39d71738ffaab8730ae4667d8e232dcec9eb8b826e993c3e263f28e94004207845d2e8845a77b58379d6d3f6efedd98e5ed902e8098c1458eeaa21ae5cc4d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h882fb00d680b40701b431ff8f70c8d513345913ea9888e9b7e36b9d9f20b4cacace89cbfd536fe46f1c399ef2c7c867a787af05348e60fede8c32660f81ef8e139cbd152ea74a7b7ec4703881ad4474bb475a9b6a771dfcc32bb9b7ef7050b69eb7bcb3ef2e81df3c207287e0fcfdf17cf1e9ca1939e1c6c446f7f7621dfea5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had84eb6bc8451f2f16ddbf52b39b63a8d33c2b16d13cd8bab4075bf7f2f5da0af330816344eebc95834ff62ff24525fa00f52d4316507a97ced84401fcd1fa5984ee98b42e5322e2204b5fd6ac550c3507c70fe25bc7947a144b2cd923b23ca6e8f1ae4929e42fd7f6f4ad5ab272e737ff6f67ac1ea5bce4b6d40630b7cdafdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb29dec951bf3bf4c4fa88b0a329024f85fc8cddc28c588f1559dbfc55470b07a51e41d474105c6ad73029362743ba4e6657f6d8421b2d8c93c9b996a2b0620d40562002ebf2630a3be471ead7a79db640a8412358379d42b339f352b255ab74c275157282af0919171ee79260ac3d1f51d0e58c2bc7bd0feccfbf0403c29742f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ffa0b9932e60eb177bd05e194a0a095264648bc1d3e0e61830f393196006574bb353d9e73e11aae9d68ecbb3aac0018793b0fe30ef58572d916b696b827cbdc9a9ee9d2e856b32d4245a606ba232b6d64e44c7ea1d698d8da1200b5841a63202bcde878e5f920266d6416fe8345f0198684b2a07e0b186c71554a18cf17e850;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6f7c694cf6352f59368de1df3612f78358d9e4ff31a522157bd484f3eea30fb23b691f79b4fb121c4f1ebbbd861b104f13759937f86e9a444c469df2def7f3b0526ddf96d633c4b3e8d72a3ae5923d48c8c307bd0211a270d965f1e89c193169411016a7e40a645580cc170b543c7ec37ac9ccaabed2f7fbc7a12b68160a63e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h521381321d201153dc8de997dfc3b70347d2c24040e5ea6bf41489682ac88631d53acdca599b9821464ded4cdf40adbf237b22ec035b23573a675c8007d5d0a4cdfa73f42a658eb4ad86317431201af02180bb6bb1c3436f88b3e74278b42c567e883c79ac9b71dd11d9a96aa2b329ead0cd9228245d74bbf1147427dd12c965;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed64323d93e18a5d03db6697f2a8f698ee57f7276e57ad6cc37a40e67fa3338db76b6c75b357366ffa5b3e7bec20326444bfb29e46ea717cc508ea233bd176a08fe53428f2934f1c508cf4d93e9ad039fe660a35a4e2ceeafab9e1d34e30b49d88abf17306907b88a8a1b6b4c7690fea5a7180431215cdde38c47308c92844fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h237630bf2f9c19195f0cc7ebdb40649ecb7d25b8acbc6f3ab2610665c4dc19493cd4d4199c819c322c1f719d3545757719b366a12aa8c61111e9c235a6f0163cb1735a614fa64b0e595d495176d9e2d478bf3e15346237485345d29739722504751613e17f657ca61529a8c81798a0faf2e688d16acbcb554c5ac1e992cca2e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1835f68134b0de9a8c4ddfd077114fc5395919925c557fbb2f64171827e3de18d00fd40156b263e03aaba129f1776c76fd06535d691b146484aed23f895ffd5f868bfb4d00e238c87b972a008ef344b495645966f70b254420c2b28ff3ddce1058bbaa590817a23c1e1d8935d7c045aa769466443bb3fe31fd1918aa0adc304e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h323d3c8a4272f9af1166f9feed9708ce53ef66964c53930dc2744ab678d23833b7550455914683ece833abd3e41c1650bdb061321a0be16ecb4161405c1972dbb8b06a5651b715c0825f51e2948b2d227aa45aeb6fe25b3a26c8d0221e24db9b0370c6af85e963ba83bc092d2c3e4076ae4d014d3583d754ef41690a72aae7a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h887dafe5d4971db3f9d9bbf3f7c65f30de213e2ae964b3e6bce6f17d2566b6b959d57005138df62aa9abb3877dfd30f74f8cfbab9634f26c3399595b732f0b30e00daf4bf4cc3218633a7020250d374a2cd059f32845046dc52c655398c460827e3445e86713f34f9a6cf2bde271065ec756215afdf007bce8f7c452a45f86da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25f8f4d1d7ae216c9d464e865d5d68dffe8cf70b4b9bca324e1db627a4cbf4df41174c2cc5f5c225e0e93a8c0f259c1ec51e5cbeb1c818e7be0454e3ee44d382d345ad8c8729b0db568af54a9e613d8854aa4b307fcb7cf55b5fbfed241e9725f3aab129a8edd79ba01665ab36f93a20bd24ed404d952ebcfb36cb7e812c0c74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h253b2f8191b82891484e7ca76b855216cac7dfcecdfac0f7b0b46d9a2e474a3e720e9bc4797229909b97ab137bde8ac52699ad8862b6007af48972b1471a1f727eb13cdb08c15fd9161ff368626694948bb1a8a31222c298cfb681e136b03d7c0372249bbbf1344c2de39b454edd5fa11071a9035d9886ba16c8556e8d9a30b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a0aa044b527143d07683e33c2a7881522dcceeb64c2d9fa1d443648620868940f2682b79a58661c336c59025d7902804b4e669a9cdf978d934f1bd5fe8a7ea5ca2a9ee5c06403620d432c9b11ca4bcbe0adbb8c42ac8926447afa34b9d9efd44991171dd936d11502554bbe76caab03828389afe41f1c0bf4cf3f8ee953d5ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea9895bb436303fc80739d78b8ad69245dc55b310c1af360282a7e9e3320b73f6e1c017834cddbcf5ee7325dbe042fdc152eff325add79454b79f5119938aa2a0eb4a2a1032036bbbd443cef4a30cc20656158dc718eda01bf9e1841b34d179d3d39c8c9efa97692c8489b1db08066e79377431286e915250e13dfb1f8d766a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28bbff8893a7d5c35dc972cf3138bc411928cfde594562ae6eadd7c1225c9e3fb722c7773ce3dc08157cdb40afa74c2e4de37a6441ceb98a27efc7787548d579bb3055b3b6dc2d905474368ec7f7ad5db52fb8dd0b04e5e3e4b4c031341ac680b2b37969629aebb70fa469549c0ac1000b0cf36047a59fd228857966137480d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f604a21a0b99d2aca4d9179fa8a10fc9722cb4cb178c026edba4eb707ef0df7df875adc0fcc8fe5fa7f0c687207185563005e5232c76bd9b5b7528c88991020f5cca2769445a366edf3eebd1164217b795784dcf041e737c6d45b18b6ce5f18f44107c004cfb14c9446ab8a4966e21e7a845d6df315e93a7c3e046fdff9c97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80054c3b343c02b2332c8e179a46781c7c8b1a9ceed903304b916a042ce2366dd4842a3291307f221c90a497c395c5c3bfc578e28770cf45eb75abee37ee5039fb614653a28914edd6c1ac3defdea74b9c68ee3205877b41dcddf7f1d2e1341f3b24ff192b30dd32de327f0570d3892ba880bbdc8af368014e69620320ce555e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d75ea770e6a13ffe7fd59b82934401c4e25a532c38fdaae465d1a1c301f962c647daf7495a24f0f483ec4df5c8e6bc58c3bd2e5d399891668b90bfb9720e157db22e1c4125560ade3eb1a2653dafd4bdac75663d1a67212f7bb926d6242f2b135f3da08ce0494b6385d508ff571365a01ae148058cdbdf5fef9c1d3caf9f8d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70d943a27d45d69a1f0f0dab114b399bc9f498e7667ef0fe2b8d110aa41a8458da0e58a98ed61796557974675f15056a6d21923088677b761baa63b8de2c30f936f9119a489da3e817b1a1afeefc9f9e81f349d3d014ea87274609985bf13bc96f915009cc525e440cab83db90029de401aad5d0c97ebefe6212c2352c8e8410;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb0933416db2c874f5287e4494d0a680193c5060c2a8bbaae6c60c06ee874eb51b328ae325a93032a6a4999271bb96f5fe08a6764a659cd108cc00859f62488f489e6872ade7f0c1c79ab6244ea1532c5688d8a09e351a965b289f820a49d6c69728da5b87b82e53183363edcc76421f9d344924adeb7f86716c3eb70b2f89ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h923c1aab46ed9fbb3e03c70c9f575d35621fb9ccea9697422dec64b6a760c6047b977656093726a35ff2ec2e62b7c9454e484b8245828d754b4fbf912468fdb565bdd07a14cd514b8fbab41242bbeecc7830acf5ea70c305689a1378605a5d327ed72913b7b6bb15d9cb5da0836162fed66aec070ad9f3ccd34bc1f041b2b8dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ea110fa851941feb9998a29451706bcd192dc5afbc6e3c93a914378ef87f776ea3033718ddf9af35d337069cf43a30531787f4b509a20c0c86cf8c71ed4ea758c06a01d4edcbe052eceb0e2ed3fa837131f77145ef3c30e35f26e1ad4a7fa9400ece1873ade08faed89063e3755a8b158da766ed2757e6114549df8d97c0dea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8b53dc48773eaee9640c62702f3a887018d4f25a32c3c2ca5ab9bca32be24b423cd7c8da150ebb868ab96dc0f4ce697250e0b4a0e4358027b0a280c2277a20bc60c25a251c4e708bc46f63084f7d994196381ef38ca59a03538acd2f46df5970fd1eb206299bed98a7d0422b10a56e0895b2b8fe0b076cd94eec3914481bf1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h873f520f7c4a70427efb956b8d4d2d94903d519fedb3092f422dc2ef8d7c696424a02c36ad87f402230781a4f5786ad91ff3dd26268b8b23fbb527d4a26814e93d8ccd924659935b578c8ecda208f48616f2e240254bd585fa1abe8ff72194eb4c9d26bc2d436120f1e2ab4c05853b29f8bb3f4ac73a66a1631ec6a724d0479a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha02c7ae126437b5a62c53368ebb7dfe64520d24199f294d2ef337d5f8b1a675ec28a3f4da19b0c6417e7427292179642cfd5c702557497681579ad9745d4131de951a999f2516c846c593b87772284153292224af4652514f61f16997203744e37bf59441a2a76cf56674ef9972ce8d6c745b6f588a7b47290a9e8ebec92479c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26f6dfe9acc0a19aef8427d4d94c540b81d61cfed69d349c7709179fc34d6ef32ce9439b144f1f669abcb23a6abc764c05ef8a2a9b000185ca25633fb140c807ea760ef7bf14b63a53ef58970fc2310c1e4f3b2e1662f542db1c7fa655f38b05009c690087754dee90e936b15162791f554bb02f8b142a7011a815dfc3a27eac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef07ece5a69683df6094e4f0d917046d4bd7db8b2717c2d42071ce952545c26bacab1b7f6d12bbc6ea49257d91f11cfd3c349700629163a494498c7b2b21cb8b77d155d19d3ecc5f0aff93ef7c53ef1dbc0dbfcb40b1031bed2e9bf36e7b63c06131498f5586cf92ed8e9eaf1147dd163bd232b029e42d273dd2d195dcf1a306;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcea8cae3add29575044c6c8fc61ddc8353aa98b6fb0d1e92ae429dfed1987693c8614665cb502885df99d493c8f0cd7d9475019c2ba69f147bcfb7f2b9240ebe7f0715a1a9f74b70633a404873d81ed7c6dc0ed348a3201c1ea8773a9d498ef021e71b07942c73be7a77e94da245de26a75140741720c230f123471fa32ea9d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3850fa0abe85a79e3295563b14db620cc30bafd8482fe51084b6bab5773fefd7ba5bc08c261b3c2d4c121a984b3616f364701b5e49d94713417810773391cd7007734a9e8568f2ca7afbb6a69fbd98c9ea299d12a0d874462e639981a220c01f5a145124e4f9eda9d62507759d61d6d2f6fa39f170853372ab7c8755fae9d600;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he76653b0bef3a46b5c60d3b82f70d119795056ecb29e55b942e64fd4ed9d01e475390490300be8b00f0570ca86393373ba578bb0b1cfbe47e2a59410dca9ced05b06e014311470fe612f59ad59fc348119fdbb4508714a0b3474f4e82f50e880d1a3adf9ecd35d24808af5d5d44f01de0102df6d351a9a1ed07b8a54abc1122c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfede5db8167e0b7d66688f34f0596be294ef13dbbdea109d6c3e9db6c615b08c36ee86c1db823552e93df6290c10855eb040b8031e44758238b0533824d67777629f59851f8e9a9a42d7772c771531b76cdc959bed2ec5331a6add694c08730d1bf8fbaf2cef62a67a60f3b91b8fa6aa6ab0d182c7f19f6565d9bbf70b5f9fe5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38f4a8b4b5679b1c7e6bafe13c7bbd1d3eb813f8810f04dbeea261e9e5e247fde0a9ed0ca9ed310dff8d849879006cfce881897717825b67fa885539ecbdae44e46f6b8adcf2e05db4a35dd6651a41ec804d0c5276a3e7b7ee21f40ef48a350f63c90f6bdc5335dcb320685d5c62f4fe652f5f7adc439556dc5bd67a8997eb87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41d85db593b7e949377d8a0b0e6168329e547a822e9476e91f58e577ac32a8260fbe7d5c45fb45f95b06f0e4f64515ce5011aed65904be2af5f8f2e2f98e83339d5f708da61c1004b38c64469b8ec69a316a7ab571da6d62e556df9d24aa94805b32cbe55b3d5a688d49e8d1e79ebdb009d07be170d8c83dbb28f0a6db75b23e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h777aeb62de5249d8991ed75150ab65994ecc1193246173bd6fe06e55f38b3c9707c3c0c21469a25cc2f23564813169ae6e4b0de94f2b8380e64412de5bf6472923b47c472486e053fc2f38de1e2888cf52b62082f50a7293d0df13a75bea295bf223787ad044bb31f1b6d9e926adba9f24a708954e3518611b0ca1134c484a7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dccfc3f73d035b266e78582af199bc615bc665b05b500170446753c516895abfd9f76bbd5db1e6264d2f095098b12794e18646ee869599e93af78c2901124fa3413410499be6eb71361b008340be2982eb5ad2034e622b1d3aeaebee20c703651823f731bb5f619b4481d8b9a1c9cf42f71a9507997f905625911270fc3499d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd61dad0d1c7fd7ff0fcb49484e803b650a165b97f7db2b5d80af297dc974ea7126235bb3263428e64ec220cce1538e4e3ae7df827dadb8c6eb8d715a58ee6a1860a815ee30848b54236e9b926b016ae4c9b0fba9f737b58e39a1188c642f44c9fba60d7417f6de1bbcf88ab063194de828f0cf55de96777ed9dc61871d85bb02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h672a65f13cdc0398f8d30c5dfe5a6f487140487e7660ff2017dc4a82b4a0cd8f86d09aab454cea3e145746f58057897dad9c927644af13e55dbdc48082e3f55af76a46e77beea67866cd4b410c9917daa5c005c16c3016bf7c63512ceba96debae3f328d8d905da7c643bf15aa00bc8eecc387e38ece08638b7f31f4fe72c482;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b76e1cb5513f6fe18a2d8f94c4bd545bfb551c32aec47a90814fadb7858d5f407503b0be8724bea751700f7797d567c6921b49a2a4bcd09ca3562256cf9dcb921052f016eccb5a888e78407f7c27adf5b0b6b2dad9086489e50dcb0dc6a611724a97d88ffc57eb110c2412c236dea04d2e8178f33bd35a929d6bc37bf245498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfee965600afff188be467a51e8b93a6058bb5699ecc97bf9f3f33c16022b546d9c0fa304ebdc801a76c097591d4f97b7e2c093e4ca62186349972d15bf6a0dfe58757cf4ce78856079465abd12f4f8e308be61c15def77dac487ae52c58a6db9382055d08ad7fe74d584023fab2586e8dc665945d19c8dc0146097ad77001681;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f1d21f361825c6a240c45bfdb81682c4f830e66189ca4d79dfd53574272141015def41f754aa2d4eee92d3220a62a0d9ccfc6f86372d637ce9ad67c9a2158553dc340b0a4e23afbb8c03dac6232ed9f797d96c1be65bd475ef5c2e8750238491b8984c65b7c996c6b1e6b02b833d3de77b2625e45c8a98f88f952da96b4f027;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7ea01569cd5ed881125e369603e8ed94f7faaac6405ec6b5c87ed5b8b61cd78e76d97843d2240b5e78d16e20c7060b84d25215d4f4f029b63bd67762ec3f17cf06114268f036a7a68522e13bd1af06841e0839c5f731620d91f070a6f82b8c6ffdf10f966481f41dfb2fd885af87d922a693f5bfb0349b627d7f89ea22f359d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hece7e1a96bbe291fe9e8e781c81571cd7be8e441ecc92f59c662abd7da3c6318267f10fc3e5dc427a5d0120ddfb0ade6feece61e103aa424935a65bbd5db8ce429be3d042bd06eb653630076af6e02e7544b1d2aece028702e05cd8387ddcb8df6edbf95b15947d004b87107a3357c81156d7c3319b76a7775842b41541da22a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f3cbbd96ad63665e7212900910f7f881fd420e7ce671a47263afa2295286223276ae00d5fff8098a35adba088f86278de832bd1549a3380d0b34176b221592c56d850e456515ffa995d6ea566145a52aa2686f89c4027c9038258620646586e618a0079f14160d316ce165020554320a2aa46a3e110ecdc96e47c90bb2aab18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65438929be308a1800c23cd7a14216b10a9489742ee18db630474bc11651b2c59cc7c8eb1ad5e4a7037a20d0ef27f44009e38ec6771a0e54d005178df3ec8c81111c2081a4ab271ad5517e95a51cd7d0f263595a066ec1e4ac025a2f8f7a9c23c40471de0f9d2f14ca50048f88dcc6548cfd00fa70231c5ccf4f630a4babc3b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1b6e634193f0a1fb42c6633515f787ebfc1be8a03b495cf3641a4a27e647ba6031cd14b571ef35b18db8eff6bc83793829276c0096207553b36af67092f03ea96b55c8c3badaca31838b468e2f814239b718f72be2668ef6b2949ce6626c77af4cc503862498160f40a3c9126212fa810149c1b6bbf157f6bb1f3c9e65fa86f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80a7c01c03260e18359a6e45ea94085c091703d7eb0cd9f51e2f7fb63758b8ce710be4894de733922241c556d533fde7095c1f297302cbbc94d1756b250dac546c244b0d3d6496dbf8c308c156a3ca25496bdbb69aa7544f4f8f5a9e7c4f1ab9e938a9b5364799a3dcd376269bdb2a3bc7e0003b9b54fec220e2fe3263a85efb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6c59096a5ab47901ee0247232c3bb5635b40da79d6f72e1ad0cc849ced7fb714ae9ed4d6a85f18e9ac1544c33ed7a15fea7732738fc825314fe1840c2c7c3438ce72b975a40e4c22e094287747fac6b8d19739bb45b8a3e6e7aaa4a167cd2e703b248d16fee717969aa39b61f34289ae5d6ae9fd5d3e97c06ac084a0b68973a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60f48210e5827e74ff78d776acb328250ccc6aee10625c9da76bfdf0cdd5b15975a0e2abb8afa32ffc03c0eb5a35defdc9b55452d04405fd1bdb748401f453cfa537e5a12082d1ffc282cd978bf24d73240fbb817a11a485f182f0231e32363fe3dd0af855cb97bf476e7f7082e0364e93dbce6a2c1b2994408330631d186a61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4f468de1541b4a77012c1c6fcddb29c8fb311a21814f1bebf56689dbd09b90982424baafb6c794d8422fc1dd99ea0cc0f01c7595ae426d0422cba6bee8104f8899856cac90a35b853f5bbaa0af0dab9ac1328d5e8080f51931cb1c9bd1d6b1dd22791328bbe3049b8a006c9fb2b62dba2b59097a146fb4c46e7a55413e58c62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h373090fa94f9adadd8ed7cd72a172b2ef6fc8c6797eb06819ab2e966d46b8e67bbc0dfb828ea93763ebcfb06521f2c94a7ff8527be1814b2455fbbad719fcf6adb6f8f3275f53e9b75fb690e62819f799a1c139ff424e7c65ade444ee60ee410c7969e6bd069f89ef8e7fc56d9292b6ba9443f2734d8072ef3734d4a471b6808;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e18fcedaa2cb9572fcdd8ad8c01f5f7f2460dacc0b27c534bc13a64d1281dca258ee6ea38aae3a19775a18aee5fd01518290c00436410fcac85f2996c3775f1bc8f16c1939fd73e6ce8d561f17fb0ca513b1e495c46692bd35c111c431d6ab38a6f46c0e33c6308a8250437fbf24e094a5792ba201e699cbd9c651922e3ad86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e79e46461fa6fa0033ae2ce26bfa1e7b603366ceaf03da6885ab35ca9bc3b58f03f0ee8fcc058f92cf79a455fad60fa93d64b3d195d155a2ed98dd662743e6397a579917dd636ef9296b4d31bc12904bce5cc156db75bccbed434b03c79137b6f0ea9ddf1c426b655a2b718458db6cb5bcdb1fd07c71b4f98cd009f9be8a498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h835df0367494b77ed7a80b819dd58a432e5afabe28686af246a2a59cc1a1eadf0aeadc2064a3dc236a6ed2b489771ba13dd601c242692d253a5ee54c61e2e0f052c3519a1bc98065d10a7bf2b1ff63e505be4fe674232f664ed087b58a5f04bc21240bcafe5051e7a049887fabd783c0103bce643f75360b3ceacda3eaccf0d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5682e1117a103d9fc345dccf554bdba533010828a0a4c24f422911cda83014ad95972e67b77785e595161bec0801919369fc09289981999ec521213f13e9e2ab806fab3ed280036721ed90b422c9770ff5f0422140fb37cde3b5590f2fab8dfa550111c1356bf515d7a3c61acedf3d6d06740ee72f042f5321bc5dcc5fbcafc3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f95d18cfdf0fcf629a0924078fd3003770532d6f1be4d30aa47fe7cdd02e687f39dc93bb83475bc2c4ef46faa3cace7a6b490004423dc43b3966c7cc2c1a9ff62902c38b08294058229dcbd3f3af0c659efd93338dba3be3f7234275331379b9ceaef5c959c06a24603b055642761c3221859724c0b1735d05925e57efc25bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbc131b541b31516d2244b58fcedaa470e4b68fb236471e7092f0d2726425b4a406ed9c2a6c7f9ebedba576458b82c43ab0de7a8e1980ce1520688c284aa032007df645ccbb32dd4e49bbf48ea6094c47543ad35de908e2243279c7a4ed3041e2cd888d842154f8f5f9c70ad6221094647c519c9d1866da239bf5988565767f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572ec219390145208168d8c8466f91fc58f642799ef916b919466644ea65667541cd313652d110b72984fd4cf84857bcce018d8736e89572ce3bfdd85a3f1828bc3c6ca6b3921e0424793e7e2e0728bebe9be3812cd2f0b63d8bfa134169e9b0b115af78f46ef81456bba6e91eaef3ecedc65eebdb6cda00e07ec9f34692c50a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedfd5f6d0764f9927663141ade3c80d4e46c459570cbb674b1beb995ca1ee1c2a458be952ace85ced828b4d0a0db54f967f650c08d7755a8119fcd29de9cc4dc66077e064cdfaaab16cf6cd32e34c34c17b11f6cc4a5d20d7d6bb48e8dc7be2edb3f13646f73360f055ff80d9cba4af0cebc91bbcd1a78d92c5125dbe17b4bec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9106c996252225ef85f438b4a55e96cee83e541c73f7d3718c9636fe7f776f0dab681bc923849fd998871a253fb1ec371889c8139956aba016f445bcbe1ea073af3aec6e1eb0905403c6522fb8bbe4302e4940494cc25e2f8455808634b8a79bc97e8d58bf090493d24246624bd7e1255ed1bbc6d131ba5b87677fbed30662cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9529ffbc24b8f5129419a40e1c37c5c2154604d1723b97678eaa920769844213819458cda2d0f4cefcdd48474e703ac70182dcc87e07062438c28b099b99f781a6ffa09dfe74228691d5d697e8ce691bf601fa9d2a19d015a0876c30204bbc81d999a4cd670c4baff2c729b56a271c23eb058fbb31cedb77642972ba952837dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a67a0045104aaed0f2426f51ac9d61b5e26a01aae45fa039fe9e655d038aaca509ee5103ed5dd21a706fc178d2885a5d0e99303792c8877eb92c99075835784744564401efff0f508f037755d6f1c21054a09c929ed3f7a57b583b8a39ffea8d193364ed6030660f1f3e992b05f2accb5f8f6daa0be0ca3dc05143d2069a6c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7a26941fb43e9b0e058d0f8130279f77bce8eeefde34d7ae9fb51d998cc5dd7a8a283abe7a62037dc8e2824e3b7f502c6180bbd6d3d3f1009cdd3ffdef5ce7884d1893daee6dc48c719a7de5ae1a072bc5d0a9120d75e35b105e2fe4f9176f87c4b2196d2c42b4493f7ba246beb3b82c161661af312469814a6b20d987e371;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546ba72ff611d3a66a12313971d8bc7dddd899f99fa7617b4c7dedba01dab3d1a346d99129ba1cc4c6b491aa2593912ea3739295fe1300602bfba29d0cdb4ebb4c83a2ac91a3448211361937bfb68a3cd755e8cb8b4f851945e7536c519d31e0f8acd23050c9d8917e89865da89716acb010e014e763cce56503d69afef47d48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8924e6be994155860c9a7feface3494a497d255db280a323227dd99a60f18fa5f51fb4439896c39390f425cfc830f4213839938c1c8289a85e780e2deafd1a0e816316cec4d8e2aae5e46fafd220c6323ce2c95249db172add1c2811acecf083e896e080a00784a94ebb99da7e2f9052c114d4819018694ed1d0acc07e0df97c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ef68f8c19413bf5528a49b5cbf6d28a88bcf87fb02a1739c6521ce9afa8958a2115d01faf2f4a9b586a9368076506f040b230a0257f10bde77c55c68f14fbc092163d02cde35fab955313a6c7bb0e8ebf94f3f7b9a34186f98ea0f9c162d419195a58398a548454c29e2551eb414477dc613e9d3063a6605cf3d8dafb637857;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9312c47b90fa112a2d5760541bcbe30138a05341bbd9d48981632a0d6ad42467ce8da27a9172878b607d363d5912f16942d84e0ea490380974d30ca644c47ab3633853c6efa6fdc490e4f872ccebfaeac0031bffd58ad48480d7c8d211b15d87e26a1d280838eb10db117615d338fd0a23380017e84615130e11c11f54f9ecc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8223e81f24fa065aa5bda8093357343261212c848735856c2fdbab0fce0518f09c7a9afa456776d1d2c6a86e299dbabc14ded9c9e2e2b1e536c8947ab53226ed154fb955e7a7ba91552c2ee99905033e78791c0793d806585c9d8dac7b6236a1d4ccc0abd10e9e389a93b5ada715a4d191d070ac42a0e2e92eebc79f9bc52fde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d836d17f9219b5ccaf39982af90f81cceaf757cbc7303da9b84e91c87e223a4c979b18c8d4a8e3b8383a4124c540df338e760fdb0d17eeecb399d8fd2d204560abdc3e55b83a898afae0f4a0d6b4f4df482da52a353a6da0d722119085bcb57dd25a96a301fc1b7f3e4a19443b8d41e6f4ff0457fddd11f2b942f805b614edb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65f9cc4d84e77d65421ee60ca77abb896d6dd31222cf699d5b0e316c9d22c07036918f4fd6069dea3fe6329e1b6fc2ed96cfb0cbeacea65d2808ef10fabc7eba52389cc98a0c016ecd943e9e5e99afdf584b6bd1ad48b05250b329c79b61ae5d481ec467f9ab045ea971d360076db5a3e6f3bb020aebb89f1ca6b41dc37038dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6f72ae1984413ade2c983121a2206932b2354ecf37a180abc7af8d2061018fdb21480a0fd1e98ddc38daa32404f64705face997023b47f47277144344e943ebd50d4a9359800a94db72949db5b9977940fc35bc34b344a17af66fbeb4c36f11189bbefd105f74bce2ae97411a53ccfe241fcc0309bd0fde4c63bd0841998f7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61433640a09bc2ccfab29f398a7a6782d93dd0b7c487f736fe93f7aa608c499e69b2ce754cbc21cc88dd355cabadc6b7eb379806a699cf0070c175d1f47364c1466e495b60209b9edfb25d2402df02a2c1a6a63e51ab99b7250972034808ecabf86057d62f3c10d73990f3bfa2dce22f01dade7d6e574b37021a1cd00ee0f9b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h173b56144b72aedee61582c977cc30307fadada6fdc7dd5ff84bcef9ba34636d8fd4d1b006b15421155b6c2dec71b01c057f809edf1d74f56fcb4a5331e593cedcd32d4704e96778f258f34d11401bc3947ac2846887a47cd72730718b718a32b1d7b636ce89b45811ef1eb590d224756462627daee2cd7a40831df8b288505b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h980dbd71df01ef8dc1e86c81451b95d49ecaedd03fb89e6bf3b2552dbd2e3976b6c87ccf552034b60e1b711262acd862b3c5b445c8584b71f353a798a8ec2fd8b9ec31c6b23b73db656bc3ce7b1fb396463d79cbc63f15f61da850163a3ad3742fc5749d7befd6087561f675fc2a887cd53a0e50412268a61c8dd43d83e3075;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd91b85459f4ee79fce9ce77a90dd37b588dd7f1dc04458de3d5cabef9def9c4f8f2efe849608376cf0b5696f0c77b755da2a3dae37048379fcedcd438380942afd0cb016f025f8ad4008c0499169f0afce50ae04e2a8ddab0931e3beb3c48f2f4628a33e53c8f6acac95e235ca9c9b1a683652f6f2efe9fe162fa899cd46fb31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff7647273a7d12a0644148a9b41acd202beb2bf23f68149714e9a8f1ba2cd313ba5cdd4181e325fe300d3641ea1b50dd65ab5f757b3612e53472c6b353569b79dfaf65984250150c546b799635162890d2186cfdc7a09e5257d483df6f14a731b75d7047dc728ef78d2db131c27cea996236a0189addd77a3b4c7e22c232d30d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70b0cc60de21f91e8d3e8de05a92625190a842760dacfaf7740cf4c18c33db268f554ea03c843b62640a126d65e6c2991c52a0bd323cd78cc2b63a8277d7b2cfd0d628fc72d4eaed4f2baea6233e767d016b966296a9f7ec3c33d7ca051de6045dc71d59a6fa76cfb9faea5ec159a26de3186c27cd36afd61db552afe3f8479;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha767c783d3a18523f1f0303bf97a6ed774cf3ada1ecb836e4305b42b160affc56c2b6b1c90276c22034ba5bb82ff76bdcbe8bec25b004cf47ef2fbcc642fe822dfdb521fb2b6c18829826eb53cebc1a028454f402f2c972b2294904ed0c88df19c8ecdc6f7657af0a3575b2e5d11288beb18679f3ce88823d65877f1a92047c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe4ecfb3eb12e996c23268f529c874b0a98288345c6a7cfb04a8300a044810b09176760e06683dbdb3559bf8173288a82d6d87df7927f9cb355a3b75c9fcdad561d5e91dc5ffc26a3c21a001d581d2ad17079c5a71a72a8b2d6206b4e0bde531e391e7d703dd9f82456fdf30b3f51959974965a6b03af03949a0af67c1a717da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc2ce726a21c5f7a749efe20252f942636335ba36ff545340baaaa222a7e1f13e4d79ad88d2b34cf5de87c3117a0f4b0114f6b7dd68e2b4071c8aebec4cdee3451d8a02591a2d726dea4103f8e1a0a7d9c7f7d4a6f03ea0925d629db5126a80280c8793de8f5100f326b1ff487918fe870e1c9aa6d267189fba4ba5163233ebb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9fd087ce66eee06a90cd25d7f83299c6bfdbc43114c071dc9ce885f04974f11d2dfd000d98d92c12c434ee5a1cca2712a81573be16547eab9f3cb4612eff360d1cbe0ac697cfbdc4d23945d94926b4bc65bc6882834bda2240a8e479158b347d1048a3cb491ed353b37da0197844367112afcdfbe648e42753575bf442539fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h338b9334575f5a34624ac8547be8f16771be9175651b55e3d9b41f8b256fc26efc4ce087e79ba0491957438c0ccc62a8075740da1e87c8b14eb308f25e43ec931c0f05d880be45f10a64f949fa1db5a9374c0d72e891570b98668e87399d265ce3b03d7ffe705007c8e64e1fe52af0ee2927ad729075e9a5402269defb42be1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1b54f684a9ee7a12b94869c0a72627b20a0e02c55419883288c0bb5344c35f028fa954596ef638451c210ac3378438c95b53f5ca209ff23e1a1927110280cee3ecdc6dee5f533e68e90205eb74947636efd8e67fb44bb2c3d5b9372384fa2d720fe86e9845bfd9a0cd2354d19c1e3d09f1fd05ce55acc17fef4987867041c05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfe447b02a13a5c06770835eadd88c0e93016214993e17974b7465ed48bae641426aea449353ee8da94336f4601c264b99b94ab59976502ba3fb7ee55102421f2dc8cbe8d1008b8a048549b4a98d5fe9849e2ebc0eb97054b7f2297c88162db50662905b1ab54f0b85d06470c836c563d16f2af64421f5046d4ce6da424b15e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57680d812df1e92725136871a09f3d2ab70423f419490a1022409fa9fb38918ff5798307068d663b3fa5e4d15d6f96aac56bfa745ba7ab604337723fa4b0dec883d994518d708da6df202944913f1a5ec1c0eef0941d53a54c0f8046f32e45ac47d43d2719215963980cf5e7050f364c5abbfaf41d0d9b2dbbd860512aee105;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3df0fe5ea2c2eb488b32788f8581f2ca5ea45701b1685009f64fa242ad053dca38af158aea207205ddd8777c59fdb86b2ba773628220aa0b7b5f4599bc2b1f93e1bd8d45dcc696a784e93338b93199e386bc3c8f358faaa6dc92ff75f6aa92d7a1e5bcf2d690c798fa7a4d6c3faec0edd45f93a705f6f69e94577a989c9844d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d84c2554338894d0da41a1efacc1a5fe2c68494d99de5f59dcdbb5a48396622d50f85799aa45dc79f10f1505826931f9eab9b2063c1eacb9ee2b6d2bda4c15c674eef269c1252bbf11dbefe28c26a9b03618661142ee85e1957ac6f6024138124d6ace19ee011f8bb95577b6a998282055ef94b3af39568a8804c8f274f6b08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf034e4071a8522d95701f2458a8f4922b37e97a9498842d528fdd68397741b2bb178db4887c88fe61f02475728f485bbcbcc7f33d8548808a983fbb80072bee330e02dee1e39c969111ed69a64825d65947823f2f688c95032ac5d07db416a83311eb2733b2801ee51728dc74c5e95a4213b1783e62cbbc35cd0c02b2c126b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab81158161ce5e220fc6dfab6f9a47e4f247a0740cdf301c23d6d0395687293de0372bfec274c1f42295d526d400bbb06f72c6d038de337f12a9404572fce8f40119188a01e6f7ebfc3d0712c7573092d601dd33460c171b5a1c9b098153ec82c0ca0aae7c76ad786968f0ed4c5aa861b7090db983eb2f178fdf0e7fa2cb633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd217e600ffefdada1eb8dcc4f6fc06bd457216b640ed247f8b25fde9ce44ee0a41c8936063807113023c670ccdbb6b7426494d23064b0ce27ee64270810f77f6832a4a22086e8a703a2c7be469be2cd2f454c1c714dc9c171f335bed8be464d09a970bc1c6ac1f4c6becf8e5c014b64eef6febd4de995e3466c3598d06b57d02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5315fabc24c4fb65d924723c22f50ceadbd39e0385a45cb140ebdea961b0b61befc71eaf390b7d93b0aaeaf77eb47921467a33375f1d9242dcde18d67c5c92d5c7d248806207e583a05eebe8e0356848177aa8abb3690895295218d4915b36e399ac5ae3803dfb5ea05732cfb8c9dbf55ae389bcf2a0a2267b25a6a9ddaf31e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d6762a9a24e274eebe0181e0274cbe0530bd81b7cd56c5baaef00bf67b921fe3953a9c90f17cf7e7ed386ef1d2328f67e60a100aa8462dac463bfc7e822a40b1286de76d24135798ae50c75472493ba994b5db2a8b1120823337625ad918586d99dff4df8dccfc005bf6ecac402468375bf79d530fce77e74d50610800627b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f9fbe99869f1192b92d0551733c660ea98232efab2b96aeb238e1a2ed9ef45bbafbc87300f5fc8628eb6da664e8ce1add12fe8500ed54a9a8e178b059bcb9026f51bd0de0acc1af2124346ead4e990bd10e6f1517f12c091b25ae7fda8e619a3a8df953e76389123324aebf1e2b97750abb5a1193f3b56c88d6692709c3ff5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc538c09dea9fb24df78eda8678596f3ccbbe8bddfaf00a62f714655f2b2b3d4d20ff64adf93bdf09f543a7567bf5225cab476b7802a542cdd98f98562dc957e576a40269d998dd8dfa854132790dbd329e54b5fda3dda893ce4eb56bc7b60a868421e404c389c231ae359276cdbaafa7bbaa4062d4e5dec1144a4dcb72e2f1eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a0bf3b1c9945368ab95c729cda4cb5356876061bd179f7280185020e1708e826350495751de4b8f408ce3fd9b7706276bd19100b28009950c55cb8d4ca0ef79af9a71421b9185bb0df1d9f99b6cf107fd315d9ef476c74f5194f44c601f546330c2a7a0401bac6fd34a82ddc47eb4931b46c5b6c18175a545ad528bcbf10c09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82af32e288819776ef280a989a86ca86de5c194bb9028858737ba2ef6c037604685a2f2fbdfe0c924667dd32749f13ae5912dbd3fc82e0dedd1079ed1fd51c01f8265c4cd675b538ffc1494673e4c779b91e64461d82624f96cefbcc6ccd61a683b15ee40638616d92e561a8e3fefbc7af38a1debb4961a7ce8f5c9b68fcb488;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69ef6494267ab2e4755c088ad7d9eee73aa110f773070ef679bde78eaac265fe3f59e9fdf31c45073811cca48c5d7242284a7a460b08f301573e845a414372c3a0b424dd60749c81fdf9c49159824c56de6f13246410816539f0837d4efee15071193ceec63606c49d57e2a4cea89a011acae0e17a145ad4d90da9157be5d944;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbeb066e243a54e1598e2a3371e6f1b3b08fcafc847251abb54927e6026b60cd4a4aa1d270f6308b3b66c47989fea1df9e0c83b1ac13da5c64cbf431e92eade7029530ae08121cf2f2f218b40edf9d6c1f84cb3fb88fb85ca8fa65153f9e765ddb3f9320693647d5b0a153ff25f4baef81061692a7da32780f6bf928a68620d98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1c90302ffe1a4a91ef010c042642697d49920175fc3ec2de02435b90a98a79d5fc6194432ffe2e34b271036f30ca010c94fb3907bf7fc756ee29b67d5e36846d45ec5b20a2bfd078c9c951ba99230afeead6c7b3cc325d35c315bb77716dc07adcad6008c32ddcecb8f549a67e55ec9e19d890c49b175ff145e12ded69b1686;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dbcdea7542223ba755bd255858d74d49d82a1b78ac1e9d9ab6b595a941a7bf2468e33149233b918c2b7d02ce7ce1311ffbcf8fae1de06bb4e4f85a771e4b490f7a0451b4d816e94cf8dd5b7d9e423d1326241d787158e2210e0a1f035d69ab88341881c52ce4dd26efc8ba7e61eaa1a2d0faf87172934e26ca5f1429397a741;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h747c8007689db3137543d9c9360bb460ed954433031b984005e1a741c58f820a119e7ec18f53f4c0c32cfef02347189e430d63cc22f099c65f34c882f9ce4493826c8929348efb44746b9e2b13a8642e6c59eec7ac1e4a16789dc13c292cd9d0a2de7ca656e92ae9b9a5f910f6467c2f6c7fdf4dde5f7c96bc055d1f3c501adb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c82bbe241c37de26fdec5f953fcaf75987b66ec457467e6bff9084fe49eb4e5d184328af66c3a3b2a165e8fd5f23c1911621ea29a1878bc69f6eab4af4dc9c019473c34b812b57ad3c1e1adc2c74df1d283acab71f44e95b684bfdea469973d824e8b0a6bd18619334872d32f4459ba06a392722c305381e42ca7612a1e9a9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9bf9349fd827007651daa182210f5f08859b7d3228f0a188a20482ee5c11da36c0d87a3a0f034aa57b1503022313bdf51bdd9883bd6034f3e499d419de5e47aeb0f042f8b2ce452bf1c524d48cf650e1f39f5fced27f0bdda26102ef3e8742ba799e6c1a303987f09b14bc3e1552198173b06fc13220d529a26f6999240b673;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb92e50fde7194074be79708a48e029a184a86f9695e8b30df27367cbe1fb1516bd59f57f9716708411d3f3b8dea74bb238a49894287432b4354885ca422b67dc8ee151cc053d61ccf863972aade632f5827538c0e136086386af50763e21d09bf1e33b187a47f7a1b3febcce660e2caf56735468849535669833115eb84e3e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffcb6d329dd8291995b14783be3519f61447a1479c421b28b79e49992d7f5969826b407b9163d05b2894ac4db7fd38fc3d4bfa471899d3f11233a5e830618746cf3c8befd507241f2cef69b232c0e4122e53baada6766381f06f830447917a0cf8b1b4a6c07a914e4bc2498b4db04460df860bfb2f40d6d706702a5191639354;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h118b484a5b5b85b1227522a7762ea1c5df1c66178b3b63624c908f110190a89ff769cd81149b4f4cc5944cef29cfa09ba752acdba5b4ef48888fa832150825a507834758756b756a2c17bd067db46eed733f360f88e2c770312dfdc3a1ed5c4f6aa77064f39da78a5b089fca5f497dae36cc4a5d140e7b82ac0e41eea6c992ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19539c87a57f134ae64ccfb142b2559bed81218782a29b694a1aca0e550b8b31937a2c92d79378c07c12a3e72743108b420bbde45e00245d162aec06354768f4a69925bb842d8006d1ae01a8e02ab9f4cc233b59f1fe70e63d246a75110866fab2fc1d2387a36506b2c84d9c531c095f366ef586b91e82849576031f23e2c6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hede62684ae8199a7bc2e4173430b24d6f9c68353d80d9f335d7a1e48078ed6ffdfca947c932f2b9e430fab7c250af2470796ae979cf3e5f81941cb1d8d97aaa6a820a3cf651e3ba10caad90f642da55bd891962415a00c14de178aabdd53cce9987cbf76bba5870fd981828cd75834fb4ff92558dde605adb1bddc1e85f7cb36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45e2e5aa2090366a21813f904220ccd8741a95e16806659063efee91b3e41320aa84fd9ec976b5f35da08294e2f55037f81544d83fe3486478b55f46c13504f13d70a7a4b08dded03edc37ea3d96ed5e29f6d88c011e7da64c4963dd49a5114762190f53062c07cefbe050f2b4bafb9ec626a1e8be46674f2dfe5f2beb06819f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6db13d6c69f967fbb94b29f7acd443ee6663f6feb4e79a6b3d466d433fc1b99bef99663662accab24073028c713dbb0d4544e7212ca7cdb84770ac0a65507dbf36b82566931827010531b89f9807bc258bfe6eaca0b82863a041b49ace7ec1b566086c403c623fb7387d666c80f1e6204ae4aec2990283eef5c057776c4a0b12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53180af39f46cb617ad543936185a46c4d6a773c2430798bce88ecb6419ca2687006b3add628ad2b8588f9fe53a25030485ff1d545c29981af4f46ed06fafd3fad66c51c1d9a68365a3640bf12d9da8b51019b4c54b691739de4b8960648b7f8645462d5e1c3503d4de0877031e2522d5fce269a2026be8139f5c7e5585ef402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88c207f7cd7a5720a1ddc55ac93c0a3755a7f052385b6f40eda1fc327109077b60b507d585e52612f327a40caaf789c13e787de0548643aad5d40119892cc808efdfd00bdfc6ab817f8ea51bb11ba2773149a93b4b3af0a2a99153d8b5d130997713c4b8a0fe9ffe371f035fa6f1532304fe4fbc446aedbef79247c8cbb73507;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed738f969eee34d41e23191b94e87abed69edd189c68ebde3850db15d9133964ce43c873c5f7bc76ff44563b0c02f797bf19f8d8c0c32b627dcaa8a15255ad6735eb27e39a9e35b6361116552bce3dec28cab0c117c923172cf198354ec0a29e655c53b5a54a5b2a8180b6d3bae4d8bc1cabc3221f0182ec08da33a1c3daa709;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2d7af3828d5c3b5ec8627a586ef57db12d27d1c65aee07cdd1ed59a8c3e157ead3a5b54cddbdd21aa6678d1ecb593fb2f9edf145d0dbac75cdccbc30af39bc15fe2b0f2738c392f23b4e3670c227ad9e55274ac3b3079b394c4f36142df1bbb1d9a50c3e6d2e1146117cd96a6a019f84d135e1610aa7a57e694f7f59400ae6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2f67eebc5ff5080e24eb09600fcc1077a07e2d8792d6545a8849deb520c8ea7b76e377603515e43af458336fb5f77babe6aae543c88da6f2a8ae147606e9529178a16c02a829c4877eb7d1f01f8408287ae37ce135c46181a9cb9b258a89b4e9f36da6008a654816702a7b486451418d620c0b7c4a89287d79c9799f2d21e76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd8bed595ca87fabd839ecb8cf69af2373cc3f91262758016c2805c3d355a4cd0fea5e762d9307738b0985c8e429ce30d09681c6a4fe2891184a0e68adfd99a0592eb448eea59922bc7fd73fdba4a7554ae112377e64b1b63c1aeef10bf64a38705fa674d4722694f2d59d56b174cd7b2bc927e2d47c63b219d7a4f895962105;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb84c57f182c581490d6d38512793c13ded6ab9bf768f1e7026d7b3e1c8aa399755f54148191ee1725296cf47ff23d7b74a374d52f74d0d8b3efe0bc936efc3f4faf4a8fed280727cebfa68268f641a19fa3ba44d1fe961970107110ef8735e1d311d3c26da8951ae8eb11260c7b8dfee8cd9ab1c9c7a4641ee545294c88493;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ef95443d94b9b65b93e68a0c9e16658fd33d70579a08811b0e301fabfc904b90518fc3a0be0d868e0bf791c04208a6abbd005df7db7185a668f136d2db7a9e03f86e61405f0e3fed7ae040630a5c08b4b8979251afabb38790f7310cbceff404b2561c1e1ca98765d9b81e8a8b84201e12431c37d0a65e9d72a16701a12c402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5153872b48da97958cfa5fd6da99388b9698910bef8c397b0996fd04e9b096b59b2f5b5e85a0eb5a67afc43d3d9a6755b369e2540d1706167e86e74131d679cf252a2745a10b4a7de73c07ff4a442eec750ed539882f19a21095cef6cfb0069f02ee4f8fdbeab201cb2dc87c946bc54744d826fa2e9e685070ef8b08e6a2dae2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa3bd745cf733e8b6dd9a45eee5c33fdb368f0e3b84d28700b966245503bb32b6927d1b86e76e13e5bce3d89eb504b6a8bbf289355fc819dd2df13a498019709a84b82fc0338be76b3460e37967907ec7d9cf295cd3fdcaab5a2955ad0b848cc6e5ce1ed28c51438ffec26a6dda0e354f0cab96a8f9d67de0e61c499dd1da4ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc51820ce10e559010c653a92dbb54a55e2141582d24a76ab62c039859302407adaa4e5f6eef166e312a42b35a56105c7e04d6b8c747a1a3e0e797a36680b3155500c74275ad1ba6389939f49559dbed15a0028dcbe59153704e84f9ab09822a79352d3f609d253fb02c097259731974787d69d5038f9229d48d4ad607db1424;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a8c32a022e687ed4ccbcdcedbdc976b038286f65ddab6f78378d94ecdc88ae15b4799752cc8e042495a261b50c5135941f97f84fb2a34488c521982bb842129aa226efd5daf834bbef34a69c9efc9442df55ae4408ca873414cb437d390f33939edb89f3434a60ddfd9525faaa3a78f5c2b0a9d5fd451ebacc68cbf17614b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d54a9e6bd9c829b2f3e82b8795911eefeb90c303bf132a6b03e54d553cb3d40d575e210651cac2fd83e7c32e424f97324e35080337216ab901e8693ba5bc9b4a0179785d3da13466c1932af23d9c6f439861a2f00c5b053c40113978c616042a538a11e9baf16770d8f31e879e57217d14965b2fce9933ba973b10c8a2f218b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f15573d9d09294e384360911e212193db7606e19da7a976c4948ce2687f8f2316c837b50553edde6c34867153e5a3165a051a2a0546dcdecd8499f9bb6b2acbebcb0d9d15e9636898c40886ab704a50cfade87132a4b3caf264ae7ab1308a9196b5db7fee851f52e26747cbdf05b47c336dcd74d177067eed6638d26a66fc80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f7ac4367f97cf7b6ebe84a4430f9c6201f5d194f3eab8fdf4715a4e4c989319d16ae9855bd5e8f418f70422c33a2603d839e3057319f16faea6f3cae7cfb991eee2ef16522ae2bd7a6328cfda7c093c7527f3b05faecfafd98c06335fb6694250590191e20ef2a626d0eeff39795812ebadaf6d561ea54a5539238637e61138;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d30197b86bee921c73b31153cef3008deac522f7b31cbdfbc45499d61c6654009253bd54102b6faeaab47e3f1e513ada31d6ae2dd29de75022880b177dd3bb782a051352b7dc06e36cb41a4cef6704f8451887118486dddaedb1199c1edf62dcfc368dd7b032b3e4ae7561c2ddb8a413c91e6d9115eefe76cf98308896e818;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h762f8aea8b5a31703646c3d23df7b51ee5eaa5055a2b8da7933ec50210928898c3e57fdcb9bd4c34126e0c341ef2cdbfb22756fe746a2710d5304192c7e9d80587875045550a3c3800d7d227abf25060c54d04a840d5c84638bec1dc80cedb6cf97f4ee19e3c390b842250fb15a0881fadd0e6d1923ded8ba9a71ae0bba8f308;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd4bd48a3229b9822b60978d35d27e6a3bb140be1867fdfee78866dbdf6d6dbfda18d4579c60c0044e55c508f3adb4566b5aa4991d3ecde7a834084b14976cf1d90d87e911988c7f1c2e667ce0ab6e914e22ab2972d5445744521e94a4c0db4a9e657fd4238a43967b9ef732979ff23cabb5722a5af2ff3293651782e1704a55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80e3d55ccc356916c2c37221e5cfd4d8addbb98528d634b24b4f2ecd376f9425041b8696b534554e88c6382074baead1255dd9f4bc0ff3142166124640281905015fcfbaf02bca3f518c741c7a56ade40da62ae3240561df3cb8a13de15b027c8bc4e0b9e261c60d38f12fd1d801371c72af541b2672403a03bdff198e661be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba909fefed0c6267d3e8028cce53ef0e8ddcf9308bec8760c7320869dd8b767ce325b50a51b9c9e8bd762b383c003de60a5911e4ab68b2039014f7ffc8f602a07f30e6bfd27f02c2624fd6ebc099bc9ad802df680bb472b8fc8e3e7d73c8f37fbe554eca251a54fbe60265f678eb10460699e9e99040c50b1b598159e445e0c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd12b678da452d6e0dfdabc85840b332daf04296643e9961ec9241b0724223a128edd00a9aefba58a255dc220c1d691ee5e95328f38a3ee73d716623ee48827d721cef5d577f7c130f480823ac8f8fa9670a4fd614353aabfd8da59a419ba5e4cec37f0918cab92e303492bbec96692100ce56f50b66bffef8917734094999002;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19ef5c6d2fa68b2e7b82f50dd2f58470d51525c32b433df0f5409daa5e13d65ff3e4e415a83d0a4726c83df5355f21520e3f7f74cc4b75c7c1a915f74d7144a68ef3f0780e39fcbad69f0272c5627399996dc38394b06c820d568428268abc0a387c9ad22336d3c5d844030948c9648417a4c8e98158a513a19c68bd8408b0e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68ea9ade1cd117c7f62a6aa6b3d675eed4e2e4fb7826e55fdbf88a9b1a99186d515fdd71f2b91935754459dd532e5cafd39552eef03d808d3eb47475baccc694d52abdee504623637ac2b7ab1f90aec5b62e45c181ad99a1d599a447c89e479552eeabf7bdd24bed107e73a2a784a8bc14747d078c29cdb927db94b2e9cd0c69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3213b51587ac367995e4fcc0cf4068752c8fa7c35eb175fd580fce4fd62a3f68c5e395c44c56d6ec7bea7b977b5fe078d32ccd36b14fae72b3e78ee6264bd3f3b967078c726946ae4aebb0f434b5bdd8c722bdfccddfb4cdb3cc2e46fe0f7f9b563fe1cc4f9c5b90c700e4908b2230095bafc32cb17abf4b0d83fdbb6a5dc9be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1694a7f300907dfb576bf012cf83d8e3e1bcfd4efae67a38e4998f0eda5794c5458c96668022508047a58b3e6a185ae2c7c38cbafe572a9b0c40824d85cb17b728beebd1ad1396581c61f44ce25387bd07e5c4693cd533b282ff97d987ca966750642483fe41ad6e49c31625ddbc429997b58eadca2509508f46e7225df4c4de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h993db0072c73a9310d539c545c64bd3f1856d25468e5904ea43a90813a7dfec268f3ad1f44c64e549c3ad8b77f34b534b847821f6923dc1478e461f2c36864e94c5cceb23b20ff1eebe7418292280d473963e3e05cb44013bd8f1e4a2e3905323222e59b9e3adffc2895298d671ddc81ec40cc73a91fe32d33b98fb042972ed5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f3ac346d5cfd4eee4dd5c0d9dcb2d9256f04fc95ba1bc84fdef368370c882afe15ff5e5530baa319bdf00b1618ae73f8030a64fc4f08bae01f3d7995ea8968a82c947edcf7d3775cd37c52d143ff4b97c0d3ce7cd7b716434d0302428b22c180f8fe6d7f31930fd6de32a1ea65a6fdb45f8a12a0d94193f7864d6fa29b71fff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h978adf6ad584779bbada01f547ca61fbb381507a08418fdbd41fd4d4fd929123ce19bf43d8e6c1c488583184a5d99b64b127b9790addc1a032c5f06ebfc963c28cc8af8d3672fcd3203f6252025716e67862fe983f26b51b6d968ed97952a0e64d0c71f9b8857d497a3624280771372f79f9b57fc73702bb0052b7e4846a5323;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2570ee0c9d9d61037eb3604287283710971d1b04a669da142c966ddacd88852b1f3aaf057f5b93789bc6f3833aa84adab69d1abb56d8caf71b0fd2994197d897c039ebf46d2cbe746515b1005ab495e3f1a4792e7f9489e0b70d981292b6e909c1d15b20f08f264a43991f313c73e63d988a415e0284001e022ca8e65f144458;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f1f224488dccd4e832a75621483e43c981eff423b39f949dd3d7ed8367f9d1b7dd276d32d3697d71e3b63dca62dac20afec4bb6fdcc22bc9d5bfe8d886fb5d73554ac529ecf5e980a8690292e9ab5605832ec38057b9f16a67713c58c7fe6fff05144b8dece1cbd4a27a93d5be766e340d26510d46e60ccfce4dca4a339be9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a60d5845be46e563532937b38f0b310a17c2921a3ee0de99fc9fef9c2e9c4d27b434148994d7c290c34efd5fad291b281ac6de30cbb6d8d6305bc9288532a6129dcf664b46387fb01ede3e999544a724efc2259a763da5ab78bc9b87011ce0c59113d0f5a0a67b548d6c6654a452ed7fc296d700144a113c01175391d740905;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he93725f1b8daa7225764e6343e590e72e97faba2287e3d578e92613846eda85abd67f107946a7556d53014305ec2c62351d50210fcbfd81c140e8ef8d4ef5ea382c2ded732f6983cb9d74129d677f63b6580721cd250453df0b89f994a977a45866ddfa17c135aa5abf606d86d2e2cfcbfae667f14563797cff63886fb082698;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ddef3161a02f89763fdf230a3ddcf5a4d92a42d1fb9ff14873e2e10555901cdf15caebd4f8ace081f3cce738b75b16b61756bc67cce033bd0246c6d87ad656e03396109c3c21ab7b5c325605dd95b7fb2d461a04e5942c3283475becf00e089e4cb47e17b150b4ac9ca7e9d12c91e0c496c6f49810c6ad061821c6d184029c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeaf11c56e91211f3c98bc63346bd850e36ac417c90bc599b5e6216f2470280a462b48a772984fa90e7765f7c69f2ff07300a8f38d3f2ce1064de386ea5d4957ddb582c189d1e6e2b43e220a4411e0cf7ce5cb3fe0e48305f8a3e6c303a7eeeee7be21ac0498991ec32968a19cb410cf589fe5738e7498a11b221609bf3f5f4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67ede043af26fe00eb0647fc139fda04fd3be32eca07f8ccff87ba8c0d3ce101855213e22a707ebef468a0329fd3c25ac32ba14b8e054389564bef1bde43f6aa49cd5b956e3f7b9b4f59891efe2090241a8b3594f4b3552cff3b2edc49afcb491fa7698e7a02aed31cece455f5407072cb0b4bda8e6d0cdb2e121de7bb31c354;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4d1841a1ccc6f87d05396942737e3664edea584d62d551a700f03bd7b6bbd8ab2e82eb735ef6d4a64bf3aa2477fd8b64cb5ee3c47fdb93bb0e98b9de777e8b5dbf57edc98a9e1b870c8a441e45dab00fb58b0f0695dab02943a15c5a1edc50a7575b436905e2270a26614468b300151df4b2095fd9909296edee3662492d817;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bc5b11fb47a185a25a66bd130dc15429ae461da0534290e391e567aa1b6d9bb6d2f4be4d3f2b9876623e026246f732f6a36fe51602d4b04d0877b999e3740a892b2b3f89d72c6f7e624c99fddae54038417d560de167302abc21100119a14e2a62f09357bf95c2ae89aa1e072c2aeaa250571328b699644b6e93f8c6ff8754;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca117dd386d164e43567acf1cb0e30f48e0c78fe61bdcedd5cf6cf85a0e8410ae23d760f40287c6c439130b2661bb8d7f37ab6811a8db5c7b4c8d8af9e0b352494763b6764a7b6608cdd1b179efb3b0cb3dbce6952726226e8111413317107c197ea1913f4f6f240c8dfc84443a6298828c889521219d1836ae148ad359db2c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3da52ea6ec6fb03f2ee7e68cfb59d51de5c6d41bb4292579b6fea46b1eff852d9436560d4341693e5fd925fd4108f91c0a165f9837337b0dc40e4564c515f2c23a4a552bd64431d5b61eeddb6c03c2f87fd491bbbb67439e43eb4bb93d18dd438ef0902172abd52b735476963d31fc27490704b0eb8c96591ec92f17939c151c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hece06c4a29d3acaf4d4eb0e4741f912d239539b6aa9e541b1265742b412c01102e9cb568ccfe32b9913ac4806fb96b9fb90ade26f5d6d30dbe6d01f5b37eae8a5da825ac1cca8dee51f8b0c16f10e34580310fdb6ec8d6815ebae66bd3222efb340b3022141e995514aa7ab315fb3541f74dcc418e247dfe372a99043997e2de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd40ce9e3f366203ee66d383b512183d44fb178463764f3df672c19f7d68c2893800d8bb0c31ffad684263ba552934b4b042f7712946c171503a5addd451d277cd9ce7b2760148fbc13dbf1bc519c92c890860a831070b3c7bfacd9163257506dcf8143842ac1d0a1475dc35c8f135a4b8171c9a77ed6c62b1ae6c8cfc6f46ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h869c1c85b86da65bb1a57a86a86e82f94e198c894626f3d3a0cc9f443d3ec5ad88fabc4edf2fdecef0d96ee4976bc6804d34493cbf0d0fa7065368365eb65d1a00adb3aa18c41f6f9a5f1f93a6ccbcac9847768ef1efc77069b71bd1f424406f29f355a3b7d8de5e39fffbbf380f529838dfca743d8aada09c44a659c4b8ba09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4c308aa4ff304b2c6d9c395bd5cf14f7dc284f18f6a5b4e33f881de9b6f20ec4162b0a99c6c1970cc53fa13878ca43d33b2080979562c70e874abbb0f90478836d0b9b3975d49a9598e1726b188049b31442c01f883a4c31c753257ece9e6ee45a18e27e232bc2684ed40f294c17d00cd34a4cde80e78317a28b63ab3413ab3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc56f1a26a7b97c18cec0a05e80a99f14de1034e8383fbff8264c817b74b1347f4d9e08f1d6519321684467319453060de231f4e52b4e832475f620a9b43df922a4f7ca466dd0b32e4d65e2ebb050d921c80d8ec23bf0587606e4899430de4d8f586bd99e76af49ac1ae2e394071986522fd1f1aebb1d0a24461c2f699615d8d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff7644bd3900c1e34ca2c6dd60a474e58cacb648420f9a05dbf49c5c8e4a9075132933139ff91cd7699eeb5e71e45ba6f8459758f6e293f5df90e4c884bd40c801dbb6d73f8b29e5864cdb5caeef9ea5ef3ff7c93ff3be75cbed65ed846279de29d725b0ffd55a808dbbaa0897b501689466c0e4d34519297e4e04d7ef68305;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc98ab73bbe69997213213e300cad49fd6bc4af5d4419b657a87a7c56430a651a813051e870befc7e2c16aab08058b5fdbdd06b1471cdf19a5eafbadb8a93ab95ccf1712a4af2b6d4f53bdf549e30a15ce3bd99937cae0abeea847cb0f3ea4c28b879bc3e444f79fddca3daf6f4cbab717e4bd12f4ca765ebe15dadd59e814184;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h197b239cf7daab7529e26821f3f0f7d2a0fbf3d2fd03cf1c8cb3e8fe672633abb15d6d2ececac26369576c02e3f8d980af6a5f38536cb9904d3714077c698544613e2a102abc58e1aaca80350be504eee790e683ca4abf8085a0d4ad7609ebfccf2e7553826d49e7f096afd051aa024f96bb6f5894fe4f5e86bdc853b757cd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66aa95322190da9b91528c6cac9290ad10c0bcbd2525d21426680af91f8af126c751dd8c6d40d7ccfe0850fd6ce94dec0b0782764d1fb174c0ad29aa7706d1a2adc6b55ce22c3a8562dec64bea041b1063bff5f181d21e0a8a03967550d3d006dd8359a33b1839cfc3880d0de0aeba4ef6f6dbce33c4b2a890394e68aa742623;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd48ad2087a3cc0d65d693312ea7fc76dfca510194caa97db543762cd23eb168e366213b371ceddca42844f4a4527b24f4603185593b01c16a1c07b29151891b6386c638212764ed8a36518e4b1c6b2551a235b34dadcabed1466a8413dec8bab101d2ad6cf0f827342bbe8d30f940195bde0c123a65bc342c8f242777594889;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1388ae471fbf0e9ce78b2f004758d7727463e18d29c96f71fb2fc2f7ed9ca716c5d28b37335856eb1b2098e56f39d0568a9b152b318ef9666549fcb2cef485731c303cbf2db12cabc01188ff4f9abd0ab1f485720dd25da01dd921bb1f487b75a15c32faa8042d588186e21b3e2adf003d1c2845a0c7ccb9215e48462ff1727;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcafdaa92dd1e5d92dbe9f3a58855e2f54d60d976be8b2d7edd9da0568dd33d48069ba70f62fb0287045905619f410173e55d687d7c291beff43ab81bcec54894f07ffa718e967a77fc29b9ee8e07a08a752c12657e3d836004e67185f4317d3c165115525a99f8eb832c836eb2818596d4c9ad26009d8e922a6879986dcf14a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd4577425f85eb8ba777d02aab2b593fdfd857c11c9ebdaee6b5b35c03faf1de500ef14364dd3ca2cfa1aa409918047888295d5d6734742a5118ea88c711c672152b07a2eb5150b29f35bd7e10a5f41613eee463554a779206c03b0860aa2bdbd0de20078a719190770da05469f7719445a5c334516d017b611f79c8445bd484;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h368630c486f0ffdf4ddc053ab23ded6b40a1f03693f3d38a302a6e2b94f4823c393a56557048d37d3e77f1c8c2bf1e04d76b64d955ccf8d0c2166f2a2c8357b512d9f4bcca0830f57cf3d3108e86c45e37c9d3fb743d1524bde39dd58d3a3dfd2159b9955d4c8e1e68c0941f179986bd797aedbdf0e8363020dc7f8249f8e3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65515ad9c33bc97caa7ecdaf364d26816bfb16fc2e11f485922b679cafddc7f4d1cb6ba1c822ac19231dc7622263245bdffcb5f3369a8cfe51ebed2ab9152d44fe5c5238666e6528e469aa98515bcd7363bc3b9cdd4afed11718fc130d11d3efdc4201a9a3382e0b5e8260d73d99e2f27e11e2b09686495aea5727d723d1f10c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40be368f16a7b2b8fdd944a3cb1b3591d661c2cdf0289358b425538a22751d18e1747eccb6c55aab8869f6b5f8e542e5f40e241f7c7b20a2651900a0f975522ddc1772226a6847e326680949ff6a10acd296ca43fbb0f13098d59052f14a7819365533155bfc18cba1f66ac40e7e273ba5fc47ebe7dd006ea5313d113e7d20b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe94db6b22e3680425fd63a5cb58dd3032f59926aac0383859d93ac376bb82bc2d6134d94fbaf89a8bd4a247e32df06099392abe30ff66752eb21043892f12874e06ada3b46ef7939d4a63fb7e193979d434c5ce44590a8eaa06a6e8bc9d9c2d124d7012ec5fc76d093b3608ef3fc0879ab637d60d8a616a68551f1af8073a2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73a76e863e00ed1d33b36da038372e2ab2e3d58b9750d0925de76f8d9ed656db5901d3b67df000efe9a30dffca032357ab7de5d083ef4f470a6ca2d06a5746ff314ecfef664e3e88cd92fb81e71285073ca89bd248d0466bad8a0201d89c6454c3d533eb6a11bb9a30a1ea14eacdc54df1a26037b481b82b2e92c56bcf1844e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4daa21393fa1b8ebb6806e4afd0675c19d2e59462feaaaadf76b223e3ec4cfd50b8b7476211e127e3d246e37b07132af7a6a6395b2d1390014a0aae873290cb9bca26bf3f78708781306126273ca9584aa78a19bfce0791be85a24b2479bb9274039fe9650e91bd3ca0050e37c11c7affb5f1d108e86911e898eb23c1b5b2382;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90051d7eb067e76cd9d23d7e16300ff1d6b79585db172c0335d04b38fc7484e4f200035456be980f7519b03d976b527cc3edebb39b4e29e34c93c11b7790f65bb1934111fb661135228dae02dde29ca1a0ee34566a28f944030066cfbac055b4344fa3de50b892278bc109246608c5c028c928d22e6b55e1921cd09f5f0c01b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbc1e2dd4b856e14d2d5ce0ee2dc3331576cf72c3ae775d61f3eac5e7df974bece5c49471cbb4f16328b7c739ec5ac71ad83f3e25ab7df970830326288e7bfc36cd3259081a6821084884b89087b184bf0b1a73be0140ce08ae3b6bd9cafb937d87be92213f0749f7fb23809c3db6a222ad571a97fe43ddd70d53580e3676784;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f25979d68c1d7345ff1bfb5a2662e7d5d5781d7fd7e2b5cf1fa0eb8d90c1168b496e5b8057d8b39f2b56969c36830e348ffcf92d1824913429fda6a8b34748d497fd334271b4b1c805122326846742c73c111cdc739ebc10f35c053f43f4f78268b9f27d6772cbaf98a75316a9f927d87e9279362544a62640bbf3a68464c62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had268708b5e95c706f0e0c1f83448a0d5cdf1e5764c827241d439b350912d0493674c122e778423f00bd34f2681223e36cc5fff1c9cacbc7296018d86c3c22716d8cf577bd73bb5e2ca42b958666cbbdbfc26d7bd4cb42b7be1fa61d008edff645a4965a74e2fc081fde74a6d4cce22f311e1b69abd76a9af3560f93acb0bb3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h156e936228b38813bc916630abb7669cbfa52bcec9fe2055bb13f1d51e59d0a417d8ee1e173bafd8a762e334afe867d1a3be08dd03a6d31883b5fec45c7be5c4747996aa31b269781670ffc26014877b51b6fb07304f5a305ac6d6ecfbd8503453f16eeac8e87608daadcd54af1e695b482d56b005d027dbc9db5ef61f85b47d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf889cbb039c5e1682759f1d5eb0c70284b14043be7f25027ca4a38c8b1bf9356586231a840e515d87366eebcf6a516475dc705ea97a17ce550021bf81b2dac21983784b83af8f359d000f9001d9bc2168d25170bf7705931c5d1939cdbf45f1439dec065619780aa34e22f9db17e1cf63a056cee6fe22f8ce3359d39ed8eef29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d85d611e04f393d982bf7f41818687e46ea674bb94a1e3e9c8e44863f6d12e08552b0be0682621abe0e6bca0ad03fd9e400aab3f73391add62ed6dc278534477186ee9e035336e84566e91b2a1d13c23f42e92f87daa9f05d479c35a07e640365672305c8d3722bd8de9fe57489adf6b893734d839b6a425476ff59575749b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h472f5a6c999c86795014e4d417f2f28e6cd0cecb40b7f57cab623f14d45418dda3bf803b75f71f0872a2d5fbf31ee8f37762321962e34a0cf8213d659276192bba02cdc194ce1e91381e565ea9fd542e281c5290e9de18e47a52c2a6f23efc828bfd9c5ad6cf6187a34a1f6cd25c325f65094b12adfd643ba9c77f45c472ac53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbffc91cc97331b13e8f484a2892d9f41621fceefc4f70bdf84d8a8faf9412715bef403f8edccec7ea44153446424f8a017229b67fd8be10abc0c5997e383ff72683dcf3c75f1b4ba8b89b975d011868fffc2eec94ebc2460a1ae636b6a8d168a09d9be980fc0c75c5e15cea71c770f95bd183e67e5454e4769ae3b058fa6b01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7953b28caaba5c05f013ba448927ead07ed35a40e7d017067e724b97da237f2ed664994aa65980f3e942e5c1d708da2a596085dae1ca0c6bbe16137da96c631ac5ee3e7a1be76471e08056a660069bdcf3a7b31d6a7048fc9ebbb51d3acf6f65f33da83314b3ef97ba1d866769b857d07c365bca51ed07fa1713fa40ccd8d8c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h347316c75962ebca03cd8f5f6dd9974c645d0d3e0a19829a75ca75cbacd4d1482c66d166e8da4b5a2b0b80cb76d36019b20f4faf7ff64acf67dc0bb83941f8ad92025ab5bfbc16be4a2ca85b3a81dbcf593a69bf6bce66dd1793e21be87d5c631a2b83d09550ae3bb2c33877d19204159f66493a46e0a4b6fce807b969f6c246;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9057483fa9b7d41a4f80b3459564b0fe5db1a46b16abcbbc1aa37a45eddbc944bbcce54ae3b7f8d745fb27097a909f175240f747e4e61a109c65837528485dbfd80393cfddbe82014763355599217a4eafa7fe0513a9e1c4e47d62d76fff7c95f48c943f51ee3d39735333fd78e6cf5d63ef751212998f26aa9dc1a1529923b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcee6c0657ce7cd4a3100b68efdeebd01cd9fe6fcf6c763e36e863315832b658876f971d6fabdcebd6197a03994de819ed2d5f0ab4d8b46b5378c2e1e11d02937b12252709cc7d749c6c93e198b8a0600d19109e0e1e907091f8e058ca0d7c5073153c951dd30dd4f0ced97197741cfe5f04987738cbb74677ec68e77ba2667f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebd0894633671c1ea1bbd7a980d496b0451d95f92dda4d29e9e0383bf613c5ca9762d49c46dd88acc88ab94c484187782e865d21e98d60efa9818ed106c0d684f4638c6c98570d858fcc2c75415e256d192f9ab0779ce8cebf9c14f9f029ca83d7a2566737dc7eca355e4c84323a966452dd99291da47ae8352fae066d1c2a5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7dfa3d354904f1717f727e65025390193e8b027f048db472abe84f4812e0fe35422be821c2e90537c10a277f053f525589dd2b1d09ef87b8e0cb2c22c30a64f6f0f0c1e0a401a7c2e4159c8f430f6a9bed4cdb891114cb4dd103d543e5b722e645fd7a0fab820613404a21cbf141485597dbd6675c2b6ad832cc07dd93dcfd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h575890ec00deeb42901917dc7fbaa402e106c945b3fa7b60cd4035ebcd2fea7f78622f3b65422b0a304577a541d94832440ce7014ec6fc3011addfc66e7ad1efb11316994fcd3a6bc13c788087c5f464cca2127e7981fe3b0558508cfbd6aecc8ad9ecbb77e4edfc31a903bb23bff745e043476c81e51fb5ffdf0c0d07f833e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c6a438ddd94a37cdfa2f1dbba4642f7a271904071b4889b5159a710fb8d5465c8f70410b7c0138f13653dc0f242ca0e327c1f2fcf70cc37dd8dcf4dd8f77ee3c245ac4b34589507673341cd891ce2f1a0b48a0f76e0caf3e16cc439bbf3b4a6544ba237b7f7ecf17a7ef5847e1f9e012942acdc0ca7e1c4a6a270d15fc10098;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33c2060ec1a2a1b6c5afb87fc24a79d8ff76882926a52333adecc193e66235ee2a8bca5838713f7533f565e35b170cd977267c5efd18dbbae0edac16970f7d14b5e5932448ab0a5ca8f39868bc68442da122a3472f1d11b46412bebb8e1354b76edcd7e3af665715d3068504a78ea43e35dcc59fac40f06e929231a047a138f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4756d2816c898211d130160654e4b3c2858f7ae17a1a0f23c567e2e91e84188ee1ce84e8b48decc36226e6cb2b664f09f997438c711eb03ee2026c83cd154b1ee7a1924b140be569a47259d6c3a83affc737f5bae1d347b80eaa78cf4fff7f1c7ce5306f3951f673cd01919b80d88baa65bfcd2c9c821f589971c2f8173e3ad5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he56fba445da902b693490bc45ad828d979625c9c2ad279c14bdb906f7c876a664e73869705e6c82554b1f9f90ca4a04e4dc3ef00ece020c84b89b35b52b0bb872dba68c6bf917dcffaed7182abd7b2fb21395825fb58f093937f9a1d9ac39c24730d1797c4e5ac0760af1d6edbfdd8821e860635dc1b423e1b5a73ca5d7fd7af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbde4869c0ab90460271010ed56e2ab9d377dddb8a98632eb769e901d220db2781ce5064fbd6bf49d5f3ae962ad7e50c817c8b7831ce02b3096397dfd1566a6324872b7e273533f5af030fffc027fb54655cd29ff92e847ee68767cb39ab0ad0d8a7f0e608ed4d91ac110d8be7b0d45e2f7de0c14403e411d2bffc2a96fd4d679;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d1cf77a9ae8f5fb1f08e3709fad50197d2ee7a31e246977b9d10730581e1e9133641bd53988dc6dcca2fb4992f2ced0eb4adfc19e6bc2f61dbc9f96b3ac414d2cded0d2089e12ef50c4ce74b8f85bd3aee5203b89a7e10c01bf7c4787b1f2bed20e6e15202eb7936ee3b29d8223459a0398dbd3a554f01de908e213ef54475c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f2498ed2c1be5f1ea9efa851cb7bb40053319b65f66941c7717378508d47c582e3f1d0f6a4686e20347ec2a17a1b8bc48af2f785d3db9c59505cd0c1a4320df6585a24d8e4601a83eff54f8147c170db5b8be0c9641c7b8ead0e6e91478b8cb7dc0a0cedcb9f6836b958402608ee2e5d917d1b1a19468c3b89516e09a8cc995;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c5856aa9bb366282c0c5ec247636fb3722c16972144ca63433ff0f4af08d441fe7fb162d8b673e790c6c5d60043a7eed6d713a0ec1f5b5be8a86bc3817b4b05aa0f1decacb37a9e0d1912bb89d9c7a064cfd93529f1b3d5196b3f02ec71574087eb1b743fe4d325b26255c5e838d0f7a6cf9404a85bdfac885d2c65a46c15a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6103b336c4155d974ec91a3bf5ae1d11ca971519f5ee0142b0a483841a834617c10824e0472a00d51101c460b55eb293958f73d4e2c259bc0945a20c32584e3d6a64241e7b6d92af93afcc983663a5e6ba5d7aaef0fa7e875719ecf75a9e1d06438e4a2d42211092c3a2a59c37bd1a068077caf8504afd7ca0cc6f2817783b69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85eff8be8f3374478a97a9eb5858a3ad35b4c25b4420a6bf4e383c1acf99b60313a5503d323a8c207549c3906e430748ea8a7f3d4df088562d1fa02f2d218d7443899fad0499f06b147716431ebcff8f133efc3794de10ba726033634fff9420d5581d7a18e29d1a33fca9e3f23b9ee118fe3d215dcdec098049f5c16212e300;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h326a3151580ad1e44151dd34f98a0e21d71fe55a93e50c0d2efb706f9afcc6dd03982a457a59f8b959a382f4f45fdd9d85322a7be291f22298a16603d75ccf1f417f2eec0a1bffe5c6935fbbc6aebf03254f54d1eef1892042ab4c1d0fb62aed26ed376aa6cb77627b8f6c0e7c50b0f69b50a403b62205a8cf4035e65628357e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9107ea1bef5329b6020b798b96d9920c8b7f20d7cf0f13ce094046df9470eadbe34ce0842d2ec26d3e8c171c9a5635e40535abf345b794d47eaf933820b8de0a13d7025b2548f7289d308ababbb3934ea6f974418150bf7df9bc1a0e6beb27a1c888d8fcf8a54bed309a107b12831f26955eb70432ac03c291869d412c67ff89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc789b4857dc4a9c16f06f7f929d0fd1a8644f1628628e1e0f990f32ca9ec021584a5cd982fc8c8437eb7bc2acfe9c2372b28c44e4fd862c8805bf89f6433a8c1b584ae2dfe763e8209417a088dc6b9ab09c4ea75ebec378e1fbb5fafe7828f473532f8d133a5691dea6c4bb928ddf2621edf599a90c92ba7768854a488ef3d4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb928b782ece0e987a930d2a8d99dc727a7bce727c0161d9566bc08371d3957825318a633b7aac80c8cd637d32f8e171b9b748083386c608daaf1d8be8a366f1f07b4413ab47b5f62a50660b47c406bd376a15ad93affcd99d01390d81c5e6275d245785fbfd79c81fe6c95dd02d8364766a0146037e0d1aa638c074426075ee4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47ba0d8391deccadd52323dca6d8a5103c80cf994223e213d030a294303ca9dd40c21584296172e23874cac129a5c84ff0150a8a91ec60e6bb9271196e1d44355fd66f3b6d42cf40db3f9ef23ad7ab5c78cdaa41b05c3c18f6e0905ebd6f32ea82cdfc7dd716ac24a180b88d97ad306200ab9c390fcfe820a94dc7d6e4487d32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d51445789f5c918fa97f76927f3bb745881b94d42f29fd8b9c6c0961cb14ce666d7d14a623220b2f0dfbe1870c8ecee30c88234da09640759c95969663a93d3b8f4d17da1c0dfb9ed2ad61639772e5893a28ed7f08cb7dc3594c6e59f754e06ac3e535fe2513c76b471481d7e6c4a81a5ba11bdc110ff889826d011633955e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13c815793e44e18b47b93d65746fbd80b29a2d5c28e85f660b8b0d089ca118d23e776ef2b5ced8e1d0e32a64d906ac0129d7b902af678a89a7810b57bc36044135d5d5c99dd327e16de883b104568bdccf8b0bfd6e3c7b65aadc39b94811fe60e59261586984ede76b0740682ffade7f1fab600e30690d0cbe10c240a056ddad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha39a1809351b79b505954024cd6edd990ad12d293612399b10238f00824cc78c912f1ef3a1401382955d6a3e87fad4611179a6ab479eef99391dca2dfa7f956dd35a0d1558c0c35ab5590a71b2838e3507c91e917e0b0f08b3acbf00cf2207d5ca9c19a323e8c5c652f114a5269a8778f8d9dfa7c4cc9cfc8af0c373978557e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59a7fc5c7bd21e0894e4cabf8e5408f2ea5cd457ce3f9fb5868a7d0cad0262b1d3eb3661392a7c815e12e14f6e261c55b8d961125a9dab1e1552b670546f8937ee4a61a8349c5d478d96ee853193018a7572769f049130bec7bb728c8534c58e3256ba2e361dba3c5097e2e29f90da5fc032cf007ef7327d82826d0f5531b6ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b3effaa97a67d03a4dc6cc9c99d6bd5bae106038f5d4fd6d67bfc0cc7a771bc03cf2f3c32ab322452c06444cc3fbe769b8352f82a6bac8ef8774b9a39a034b44de37c3f1367b05419f02415a7c6b0f902a034676b0487f8061a32a9238932359138c0367500d7f8a23d70cf82aca954fe421025afe16cc8da5f6fa333113802;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h405f5af9e9a2bc8d3eca57506ab0cca416d9c10c408c50552c76377d2586f49c40ddf56859e8dcffff72e59bd085c9765f7352b1cd756ebd966ed96d672dee98104e04d61e03cdd93c6e1877fcf58e73fce5616d53e2bdbebe37ae81b79690996b83dbcd6fa9209906b135a8fb24c3723e695fb3598b219bb51090b82726ec8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e92ec184e838d29364b67b7c48954de7ddebeb835b70eb2c314673f9d2768bbe8b205c75e7ef31f4e13f7d6aff9159e7aaa513d1f32c3e8210dc6376cadb628e0ad69ab83766155b6202a883da89ec69461ebb160b090935756b48e552411f930d4f83bac0db5c3abbecc344cc24de73062cdc06e858751bacc7c99d5de1d40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab35098dc74bb6b1a8e7b4bb776fa25cf84efa53dd9821310ba0eb4363781fd915e29b12b9ce3b665d3490cf311ca5c1389940ef54a5c79b1a32b249e9fab0b5541c9f34e94037aba3546ad2dfad9ff1a9ebf438c836fbbe56f6395bfe529abc8717108f0aad300f85628f2bd70ff9e41081605bc410032511d7619dd2da3d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82aaa51028d7e34b4be0f58602afef82b445e1c0ea247e8da963191aa864b62303f4ba70d9befe5a29c4a011de69484856bd9b96a5d9a3e7eaa418b4589164002314bf3e08ca31170454a5f1160afbbca558d9bbe64e0a4eb259ca0d95989ed9da79ae624a94d1a2c4e28d63fc88e4c5d65dc3c393f98deec24dfd3a652208b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3a2d0ec5229c1062ba284b6763f91b1c2e7c8276df20c19c4e5b759623b0d07182b18e76fd576484d34cf81cde799d8658b1a310d5cc1908c213018d258a558575956e164e9315e466462a02650f0024705aab1e8d5972d0d7e41a8745ff592a3c885d040679f3794c13a916005a10cff829223451459444d3854f8af7a50a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c16a7eb70a4ace1cc232a6de61668b5cafc8cdc27d4ac02b514654fd420fa38cf2d185850eee147fa87c04de4afc84cc9e9e3144de9b8d02d289195cc44d50cbade13d284e10ebf5556d319d6bc1897b7a610944e901a3c874ceacbfe4f3c6dda51f8475f035f79f32cc8bd0edbf397da189e92ca4257f79ce310f9d35fdd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40516136e8797084e6d15331bc71f8ade22481d7376555719a7384901f59405fa891b191f0910ae89296ae62d14ee4463a7df0285c3d0100a656b006541858a837fd10201b1f4bd4cf3b3d1bff6c0fb66fb399bcadf5692fc4f7392a44c510e71c9bfd7ae0577692f352e86800f804f9d0a7ee7b184d94e7a9bfd29703570943;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f24cbff33b7c9ac5d55cde932736f9ea37684de9af5dfc6eb3e4812b596971076c9db1c550d53590e785c3e526a7ae320953e58e82bad70451c3040ea60acaa597c05ee50feeba96d68247b241bb48585946b3bf1397575d31cbe6cc5d5721883d477ba0d9549d2c0b7db5e5d3a878969c2727256e88359b7280b8e78f579f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7273e4517bbc5c7b6371712fc8d2ad6f5b14824427db69eac83e6b27a53936e5ec1461aa80c978179da6763da15c071a1d9ffec0efe704bb9ca6890d159169e0295a78dd3dca7d1c784be6a575715f424235e2896325dab7cda30aae9f196ceae17293ae13c48ebd2ceeb0af9fbec803d095637a57369781a6769657df759b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49fa0f81e0ebad18332abac9f4f8128f665353fa63dc1871865093eed40b7d387f5047e77be8d16ddbe8c9fe62c30c281c1864763f44dadaab4f912c666a91e6d26ac21a10517eb55dd34b286ba5fb994d816b7613629fc36074e9b31d74fb4ee41b331f402ffab5f12620fe104334c41531dec4c297595a3e29bf8ae5ff4dba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52c5403c528ea4cdbf2e9c11ee05e3cd5de3275bd4e6555d93c7f73e6bf32aa3c39f09e7a9fd1bd19e706b908955cdf159034272da447cfee82ad2df3b02f163bb4868e865bbbfc8d82832ad73317a1a46efee523b14c65bbb4c3ffb34c948653c7106f31c7249216b69413106c386415e2caabbc16c79ba5b5e39c6f146284;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ab026a7b82524acf9d870244ba7c4d88702195c0229102258c1bd0dda198a33fe0c4800c876570ed8c2920c509aa558ac9a37fc0f765113985b257b8d6b78243e4d2ad238321bba07390eefee7d2c118ee4fa0d0eb89fd1d11abd6cc9e05e7b5dde2f0d31e74b083b4d87428636f6ac6464bfda36d5a24b3a03413ea8abc9b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c4d19912495b3518509e48b08426a4c4f121ba2176adcec48c908326f1220c3b549c2b5923cf67c234b04b516197f11eb645be6fa22bef70610b78315b0dfb0bee17e6bf85004261e0755e359950555fe96b835fe8b4b7e66a31d282477cf4dd3a13108484f33c6d3bf705f3c75188b0419c3d9d8e2315deef92c6c17ebc865;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66c2b9ebefedcb8611bc42c07098d06cca42e8aaad04cdacaa0cbe3f26156d6bf5897c1ea75d50a7c882d8d4d6db9f02cfed2232ae63174928370c6a5e2794ab361c44a60b89251816a9ece6dd2aefe99227603094fd9882cb7e15db483d28ae837c66eb420da3ac63fb74ae3345d0232b8d34226bf6f66a1b61bcfc57ae4a0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa6a29bf509798e51b0e5e6e5c6649fde3c06d32d8d6aa86b61fc67077e24b3123ab5971b6ad81e3009fe9b719f1ff88f8d17b923a218d0bca46120e84f01304c3c417f7f50ed9f988ff8429735fd9f29046df9239caf032d6e41efe99e453046218d26eba09ea1a58ba5b7f86704806f296f6261b84ccd6d345ae123f2c2b3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a1ab3db74f34fd50577e5f8ed18b18a3e650fda4a1f948d761a18cb19ed4a42e8466cbb423c6dab68eec796cd57f762b23a08309c9e92e84d92f78b527bd7ec875bc7de878ec9a9fbe9c07958e59d6f9069087870de00fbd71cda8c5a5a8876f4ebc24e8556956a980f7d0e28d04eaa0b8ef9e4f8cc6426c327ccd3be152457;
        #1
        $finish();
    end
endmodule
